module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    reg [127:0] src32;
    reg [127:0] src33;
    reg [127:0] src34;
    reg [127:0] src35;
    reg [127:0] src36;
    reg [127:0] src37;
    reg [127:0] src38;
    reg [127:0] src39;
    reg [127:0] src40;
    reg [127:0] src41;
    reg [127:0] src42;
    reg [127:0] src43;
    reg [127:0] src44;
    reg [127:0] src45;
    reg [127:0] src46;
    reg [127:0] src47;
    reg [127:0] src48;
    reg [127:0] src49;
    reg [127:0] src50;
    reg [127:0] src51;
    reg [127:0] src52;
    reg [127:0] src53;
    reg [127:0] src54;
    reg [127:0] src55;
    reg [127:0] src56;
    reg [127:0] src57;
    reg [127:0] src58;
    reg [127:0] src59;
    reg [127:0] src60;
    reg [127:0] src61;
    reg [127:0] src62;
    reg [127:0] src63;
    compressor_CLA128_64 compressor_CLA128_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
        src16 <= 128'h0;
        src17 <= 128'h0;
        src18 <= 128'h0;
        src19 <= 128'h0;
        src20 <= 128'h0;
        src21 <= 128'h0;
        src22 <= 128'h0;
        src23 <= 128'h0;
        src24 <= 128'h0;
        src25 <= 128'h0;
        src26 <= 128'h0;
        src27 <= 128'h0;
        src28 <= 128'h0;
        src29 <= 128'h0;
        src30 <= 128'h0;
        src31 <= 128'h0;
        src32 <= 128'h0;
        src33 <= 128'h0;
        src34 <= 128'h0;
        src35 <= 128'h0;
        src36 <= 128'h0;
        src37 <= 128'h0;
        src38 <= 128'h0;
        src39 <= 128'h0;
        src40 <= 128'h0;
        src41 <= 128'h0;
        src42 <= 128'h0;
        src43 <= 128'h0;
        src44 <= 128'h0;
        src45 <= 128'h0;
        src46 <= 128'h0;
        src47 <= 128'h0;
        src48 <= 128'h0;
        src49 <= 128'h0;
        src50 <= 128'h0;
        src51 <= 128'h0;
        src52 <= 128'h0;
        src53 <= 128'h0;
        src54 <= 128'h0;
        src55 <= 128'h0;
        src56 <= 128'h0;
        src57 <= 128'h0;
        src58 <= 128'h0;
        src59 <= 128'h0;
        src60 <= 128'h0;
        src61 <= 128'h0;
        src62 <= 128'h0;
        src63 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA128_64(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    input [127:0]src16,
    input [127:0]src17,
    input [127:0]src18,
    input [127:0]src19,
    input [127:0]src20,
    input [127:0]src21,
    input [127:0]src22,
    input [127:0]src23,
    input [127:0]src24,
    input [127:0]src25,
    input [127:0]src26,
    input [127:0]src27,
    input [127:0]src28,
    input [127:0]src29,
    input [127:0]src30,
    input [127:0]src31,
    input [127:0]src32,
    input [127:0]src33,
    input [127:0]src34,
    input [127:0]src35,
    input [127:0]src36,
    input [127:0]src37,
    input [127:0]src38,
    input [127:0]src39,
    input [127:0]src40,
    input [127:0]src41,
    input [127:0]src42,
    input [127:0]src43,
    input [127:0]src44,
    input [127:0]src45,
    input [127:0]src46,
    input [127:0]src47,
    input [127:0]src48,
    input [127:0]src49,
    input [127:0]src50,
    input [127:0]src51,
    input [127:0]src52,
    input [127:0]src53,
    input [127:0]src54,
    input [127:0]src55,
    input [127:0]src56,
    input [127:0]src57,
    input [127:0]src58,
    input [127:0]src59,
    input [127:0]src60,
    input [127:0]src61,
    input [127:0]src62,
    input [127:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [0:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [0:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [0:0] comp_out69;
    wire [1:0] comp_out70;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[1], 1'h0, comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], 1'h0, comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], 1'h0, comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      input wire [127:0] src16,
      input wire [127:0] src17,
      input wire [127:0] src18,
      input wire [127:0] src19,
      input wire [127:0] src20,
      input wire [127:0] src21,
      input wire [127:0] src22,
      input wire [127:0] src23,
      input wire [127:0] src24,
      input wire [127:0] src25,
      input wire [127:0] src26,
      input wire [127:0] src27,
      input wire [127:0] src28,
      input wire [127:0] src29,
      input wire [127:0] src30,
      input wire [127:0] src31,
      input wire [127:0] src32,
      input wire [127:0] src33,
      input wire [127:0] src34,
      input wire [127:0] src35,
      input wire [127:0] src36,
      input wire [127:0] src37,
      input wire [127:0] src38,
      input wire [127:0] src39,
      input wire [127:0] src40,
      input wire [127:0] src41,
      input wire [127:0] src42,
      input wire [127:0] src43,
      input wire [127:0] src44,
      input wire [127:0] src45,
      input wire [127:0] src46,
      input wire [127:0] src47,
      input wire [127:0] src48,
      input wire [127:0] src49,
      input wire [127:0] src50,
      input wire [127:0] src51,
      input wire [127:0] src52,
      input wire [127:0] src53,
      input wire [127:0] src54,
      input wire [127:0] src55,
      input wire [127:0] src56,
      input wire [127:0] src57,
      input wire [127:0] src58,
      input wire [127:0] src59,
      input wire [127:0] src60,
      input wire [127:0] src61,
      input wire [127:0] src62,
      input wire [127:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [0:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [0:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [0:0] dst69,
      output wire [1:0] dst70);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [127:0] stage0_16;
   wire [127:0] stage0_17;
   wire [127:0] stage0_18;
   wire [127:0] stage0_19;
   wire [127:0] stage0_20;
   wire [127:0] stage0_21;
   wire [127:0] stage0_22;
   wire [127:0] stage0_23;
   wire [127:0] stage0_24;
   wire [127:0] stage0_25;
   wire [127:0] stage0_26;
   wire [127:0] stage0_27;
   wire [127:0] stage0_28;
   wire [127:0] stage0_29;
   wire [127:0] stage0_30;
   wire [127:0] stage0_31;
   wire [127:0] stage0_32;
   wire [127:0] stage0_33;
   wire [127:0] stage0_34;
   wire [127:0] stage0_35;
   wire [127:0] stage0_36;
   wire [127:0] stage0_37;
   wire [127:0] stage0_38;
   wire [127:0] stage0_39;
   wire [127:0] stage0_40;
   wire [127:0] stage0_41;
   wire [127:0] stage0_42;
   wire [127:0] stage0_43;
   wire [127:0] stage0_44;
   wire [127:0] stage0_45;
   wire [127:0] stage0_46;
   wire [127:0] stage0_47;
   wire [127:0] stage0_48;
   wire [127:0] stage0_49;
   wire [127:0] stage0_50;
   wire [127:0] stage0_51;
   wire [127:0] stage0_52;
   wire [127:0] stage0_53;
   wire [127:0] stage0_54;
   wire [127:0] stage0_55;
   wire [127:0] stage0_56;
   wire [127:0] stage0_57;
   wire [127:0] stage0_58;
   wire [127:0] stage0_59;
   wire [127:0] stage0_60;
   wire [127:0] stage0_61;
   wire [127:0] stage0_62;
   wire [127:0] stage0_63;
   wire [29:0] stage1_0;
   wire [32:0] stage1_1;
   wire [46:0] stage1_2;
   wire [66:0] stage1_3;
   wire [65:0] stage1_4;
   wire [51:0] stage1_5;
   wire [88:0] stage1_6;
   wire [70:0] stage1_7;
   wire [65:0] stage1_8;
   wire [60:0] stage1_9;
   wire [40:0] stage1_10;
   wire [63:0] stage1_11;
   wire [55:0] stage1_12;
   wire [53:0] stage1_13;
   wire [65:0] stage1_14;
   wire [67:0] stage1_15;
   wire [88:0] stage1_16;
   wire [66:0] stage1_17;
   wire [41:0] stage1_18;
   wire [54:0] stage1_19;
   wire [71:0] stage1_20;
   wire [54:0] stage1_21;
   wire [70:0] stage1_22;
   wire [53:0] stage1_23;
   wire [61:0] stage1_24;
   wire [60:0] stage1_25;
   wire [83:0] stage1_26;
   wire [55:0] stage1_27;
   wire [47:0] stage1_28;
   wire [79:0] stage1_29;
   wire [71:0] stage1_30;
   wire [59:0] stage1_31;
   wire [82:0] stage1_32;
   wire [62:0] stage1_33;
   wire [67:0] stage1_34;
   wire [47:0] stage1_35;
   wire [60:0] stage1_36;
   wire [96:0] stage1_37;
   wire [43:0] stage1_38;
   wire [92:0] stage1_39;
   wire [62:0] stage1_40;
   wire [39:0] stage1_41;
   wire [50:0] stage1_42;
   wire [78:0] stage1_43;
   wire [49:0] stage1_44;
   wire [57:0] stage1_45;
   wire [79:0] stage1_46;
   wire [69:0] stage1_47;
   wire [45:0] stage1_48;
   wire [50:0] stage1_49;
   wire [70:0] stage1_50;
   wire [47:0] stage1_51;
   wire [60:0] stage1_52;
   wire [61:0] stage1_53;
   wire [51:0] stage1_54;
   wire [67:0] stage1_55;
   wire [56:0] stage1_56;
   wire [57:0] stage1_57;
   wire [59:0] stage1_58;
   wire [55:0] stage1_59;
   wire [52:0] stage1_60;
   wire [58:0] stage1_61;
   wire [97:0] stage1_62;
   wire [52:0] stage1_63;
   wire [29:0] stage1_64;
   wire [17:0] stage1_65;
   wire [19:0] stage2_0;
   wire [12:0] stage2_1;
   wire [24:0] stage2_2;
   wire [27:0] stage2_3;
   wire [25:0] stage2_4;
   wire [28:0] stage2_5;
   wire [25:0] stage2_6;
   wire [38:0] stage2_7;
   wire [31:0] stage2_8;
   wire [41:0] stage2_9;
   wire [30:0] stage2_10;
   wire [21:0] stage2_11;
   wire [27:0] stage2_12;
   wire [16:0] stage2_13;
   wire [38:0] stage2_14;
   wire [30:0] stage2_15;
   wire [23:0] stage2_16;
   wire [33:0] stage2_17;
   wire [30:0] stage2_18;
   wire [26:0] stage2_19;
   wire [33:0] stage2_20;
   wire [21:0] stage2_21;
   wire [34:0] stage2_22;
   wire [27:0] stage2_23;
   wire [27:0] stage2_24;
   wire [31:0] stage2_25;
   wire [26:0] stage2_26;
   wire [32:0] stage2_27;
   wire [26:0] stage2_28;
   wire [20:0] stage2_29;
   wire [51:0] stage2_30;
   wire [27:0] stage2_31;
   wire [24:0] stage2_32;
   wire [28:0] stage2_33;
   wire [31:0] stage2_34;
   wire [29:0] stage2_35;
   wire [32:0] stage2_36;
   wire [36:0] stage2_37;
   wire [35:0] stage2_38;
   wire [21:0] stage2_39;
   wire [34:0] stage2_40;
   wire [31:0] stage2_41;
   wire [17:0] stage2_42;
   wire [20:0] stage2_43;
   wire [29:0] stage2_44;
   wire [34:0] stage2_45;
   wire [22:0] stage2_46;
   wire [35:0] stage2_47;
   wire [30:0] stage2_48;
   wire [15:0] stage2_49;
   wire [32:0] stage2_50;
   wire [30:0] stage2_51;
   wire [17:0] stage2_52;
   wire [38:0] stage2_53;
   wire [28:0] stage2_54;
   wire [19:0] stage2_55;
   wire [26:0] stage2_56;
   wire [32:0] stage2_57;
   wire [23:0] stage2_58;
   wire [34:0] stage2_59;
   wire [21:0] stage2_60;
   wire [28:0] stage2_61;
   wire [37:0] stage2_62;
   wire [37:0] stage2_63;
   wire [25:0] stage2_64;
   wire [17:0] stage2_65;
   wire [5:0] stage2_66;
   wire [1:0] stage2_67;
   wire [4:0] stage3_0;
   wire [7:0] stage3_1;
   wire [5:0] stage3_2;
   wire [21:0] stage3_3;
   wire [11:0] stage3_4;
   wire [23:0] stage3_5;
   wire [9:0] stage3_6;
   wire [11:0] stage3_7;
   wire [15:0] stage3_8;
   wire [19:0] stage3_9;
   wire [11:0] stage3_10;
   wire [12:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [9:0] stage3_14;
   wire [25:0] stage3_15;
   wire [11:0] stage3_16;
   wire [11:0] stage3_17;
   wire [12:0] stage3_18;
   wire [15:0] stage3_19;
   wire [13:0] stage3_20;
   wire [17:0] stage3_21;
   wire [8:0] stage3_22;
   wire [12:0] stage3_23;
   wire [15:0] stage3_24;
   wire [19:0] stage3_25;
   wire [12:0] stage3_26;
   wire [13:0] stage3_27;
   wire [16:0] stage3_28;
   wire [7:0] stage3_29;
   wire [14:0] stage3_30;
   wire [19:0] stage3_31;
   wire [11:0] stage3_32;
   wire [11:0] stage3_33;
   wire [17:0] stage3_34;
   wire [9:0] stage3_35;
   wire [14:0] stage3_36;
   wire [14:0] stage3_37;
   wire [12:0] stage3_38;
   wire [13:0] stage3_39;
   wire [17:0] stage3_40;
   wire [11:0] stage3_41;
   wire [19:0] stage3_42;
   wire [9:0] stage3_43;
   wire [7:0] stage3_44;
   wire [14:0] stage3_45;
   wire [11:0] stage3_46;
   wire [10:0] stage3_47;
   wire [18:0] stage3_48;
   wire [11:0] stage3_49;
   wire [6:0] stage3_50;
   wire [12:0] stage3_51;
   wire [19:0] stage3_52;
   wire [8:0] stage3_53;
   wire [23:0] stage3_54;
   wire [11:0] stage3_55;
   wire [7:0] stage3_56;
   wire [11:0] stage3_57;
   wire [11:0] stage3_58;
   wire [13:0] stage3_59;
   wire [13:0] stage3_60;
   wire [20:0] stage3_61;
   wire [15:0] stage3_62;
   wire [17:0] stage3_63;
   wire [12:0] stage3_64;
   wire [11:0] stage3_65;
   wire [6:0] stage3_66;
   wire [6:0] stage3_67;
   wire [0:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [9:0] stage4_3;
   wire [13:0] stage4_4;
   wire [8:0] stage4_5;
   wire [8:0] stage4_6;
   wire [6:0] stage4_7;
   wire [5:0] stage4_8;
   wire [6:0] stage4_9;
   wire [10:0] stage4_10;
   wire [5:0] stage4_11;
   wire [5:0] stage4_12;
   wire [4:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [7:0] stage4_17;
   wire [5:0] stage4_18;
   wire [6:0] stage4_19;
   wire [10:0] stage4_20;
   wire [3:0] stage4_21;
   wire [4:0] stage4_22;
   wire [5:0] stage4_23;
   wire [10:0] stage4_24;
   wire [7:0] stage4_25;
   wire [10:0] stage4_26;
   wire [5:0] stage4_27;
   wire [5:0] stage4_28;
   wire [9:0] stage4_29;
   wire [3:0] stage4_30;
   wire [6:0] stage4_31;
   wire [6:0] stage4_32;
   wire [5:0] stage4_33;
   wire [5:0] stage4_34;
   wire [5:0] stage4_35;
   wire [6:0] stage4_36;
   wire [6:0] stage4_37;
   wire [5:0] stage4_38;
   wire [7:0] stage4_39;
   wire [11:0] stage4_40;
   wire [10:0] stage4_41;
   wire [5:0] stage4_42;
   wire [4:0] stage4_43;
   wire [5:0] stage4_44;
   wire [5:0] stage4_45;
   wire [5:0] stage4_46;
   wire [6:0] stage4_47;
   wire [4:0] stage4_48;
   wire [5:0] stage4_49;
   wire [6:0] stage4_50;
   wire [2:0] stage4_51;
   wire [16:0] stage4_52;
   wire [5:0] stage4_53;
   wire [11:0] stage4_54;
   wire [3:0] stage4_55;
   wire [7:0] stage4_56;
   wire [5:0] stage4_57;
   wire [3:0] stage4_58;
   wire [5:0] stage4_59;
   wire [5:0] stage4_60;
   wire [9:0] stage4_61;
   wire [5:0] stage4_62;
   wire [8:0] stage4_63;
   wire [8:0] stage4_64;
   wire [4:0] stage4_65;
   wire [4:0] stage4_66;
   wire [3:0] stage4_67;
   wire [1:0] stage4_68;
   wire [0:0] stage4_69;
   wire [0:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [3:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [3:0] stage5_6;
   wire [2:0] stage5_7;
   wire [3:0] stage5_8;
   wire [3:0] stage5_9;
   wire [6:0] stage5_10;
   wire [1:0] stage5_11;
   wire [5:0] stage5_12;
   wire [4:0] stage5_13;
   wire [0:0] stage5_14;
   wire [8:0] stage5_15;
   wire [3:0] stage5_16;
   wire [2:0] stage5_17;
   wire [1:0] stage5_18;
   wire [2:0] stage5_19;
   wire [8:0] stage5_20;
   wire [4:0] stage5_21;
   wire [3:0] stage5_22;
   wire [0:0] stage5_23;
   wire [5:0] stage5_24;
   wire [2:0] stage5_25;
   wire [3:0] stage5_26;
   wire [7:0] stage5_27;
   wire [1:0] stage5_28;
   wire [5:0] stage5_29;
   wire [3:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [2:0] stage5_33;
   wire [7:0] stage5_34;
   wire [0:0] stage5_35;
   wire [1:0] stage5_36;
   wire [2:0] stage5_37;
   wire [3:0] stage5_38;
   wire [4:0] stage5_39;
   wire [2:0] stage5_40;
   wire [3:0] stage5_41;
   wire [3:0] stage5_42;
   wire [3:0] stage5_43;
   wire [3:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [4:0] stage5_47;
   wire [5:0] stage5_48;
   wire [0:0] stage5_49;
   wire [1:0] stage5_50;
   wire [2:0] stage5_51;
   wire [6:0] stage5_52;
   wire [3:0] stage5_53;
   wire [2:0] stage5_54;
   wire [3:0] stage5_55;
   wire [5:0] stage5_56;
   wire [1:0] stage5_57;
   wire [3:0] stage5_58;
   wire [2:0] stage5_59;
   wire [1:0] stage5_60;
   wire [2:0] stage5_61;
   wire [2:0] stage5_62;
   wire [3:0] stage5_63;
   wire [5:0] stage5_64;
   wire [2:0] stage5_65;
   wire [1:0] stage5_66;
   wire [2:0] stage5_67;
   wire [1:0] stage5_68;
   wire [0:0] stage5_69;
   wire [0:0] stage5_70;
   wire [0:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [1:0] stage6_36;
   wire [1:0] stage6_37;
   wire [0:0] stage6_38;
   wire [1:0] stage6_39;
   wire [1:0] stage6_40;
   wire [1:0] stage6_41;
   wire [1:0] stage6_42;
   wire [1:0] stage6_43;
   wire [1:0] stage6_44;
   wire [1:0] stage6_45;
   wire [1:0] stage6_46;
   wire [1:0] stage6_47;
   wire [1:0] stage6_48;
   wire [1:0] stage6_49;
   wire [1:0] stage6_50;
   wire [1:0] stage6_51;
   wire [1:0] stage6_52;
   wire [1:0] stage6_53;
   wire [1:0] stage6_54;
   wire [1:0] stage6_55;
   wire [1:0] stage6_56;
   wire [1:0] stage6_57;
   wire [1:0] stage6_58;
   wire [1:0] stage6_59;
   wire [1:0] stage6_60;
   wire [1:0] stage6_61;
   wire [1:0] stage6_62;
   wire [0:0] stage6_63;
   wire [1:0] stage6_64;
   wire [1:0] stage6_65;
   wire [1:0] stage6_66;
   wire [1:0] stage6_67;
   wire [1:0] stage6_68;
   wire [0:0] stage6_69;
   wire [1:0] stage6_70;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;
   assign dst39 = stage6_39;
   assign dst40 = stage6_40;
   assign dst41 = stage6_41;
   assign dst42 = stage6_42;
   assign dst43 = stage6_43;
   assign dst44 = stage6_44;
   assign dst45 = stage6_45;
   assign dst46 = stage6_46;
   assign dst47 = stage6_47;
   assign dst48 = stage6_48;
   assign dst49 = stage6_49;
   assign dst50 = stage6_50;
   assign dst51 = stage6_51;
   assign dst52 = stage6_52;
   assign dst53 = stage6_53;
   assign dst54 = stage6_54;
   assign dst55 = stage6_55;
   assign dst56 = stage6_56;
   assign dst57 = stage6_57;
   assign dst58 = stage6_58;
   assign dst59 = stage6_59;
   assign dst60 = stage6_60;
   assign dst61 = stage6_61;
   assign dst62 = stage6_62;
   assign dst63 = stage6_63;
   assign dst64 = stage6_64;
   assign dst65 = stage6_65;
   assign dst66 = stage6_66;
   assign dst67 = stage6_67;
   assign dst68 = stage6_68;
   assign dst69 = stage6_69;
   assign dst70 = stage6_70;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_2[2]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_2[3]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[4]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[5]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[6]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[7]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[8]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[9]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[10]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[11]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[12]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[13]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[14]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[15]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[16]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[17]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[18]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[19]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[18],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[19],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[20],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[21],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[22],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[23],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[24],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[25],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[26],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[27],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[0],stage1_4[28],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[1],stage1_4[29],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[2],stage1_4[30],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[3],stage1_4[31],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[4],stage1_4[32],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[5],stage1_4[33],stage1_3[35],stage1_2[35]}
   );
   gpc606_5 gpc36 (
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[6],stage1_4[34],stage1_3[36],stage1_2[36]}
   );
   gpc606_5 gpc37 (
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[7],stage1_4[35],stage1_3[37],stage1_2[37]}
   );
   gpc606_5 gpc38 (
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[8],stage1_4[36],stage1_3[38],stage1_2[38]}
   );
   gpc615_5 gpc39 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_3[36]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[9],stage1_4[37],stage1_3[39],stage1_2[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage0_4[42]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[7],stage1_5[10],stage1_4[38],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage0_4[43]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[8],stage1_5[11],stage1_4[39],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage0_4[44]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[9],stage1_5[12],stage1_4[40],stage1_3[42]}
   );
   gpc615_5 gpc43 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[45]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[10],stage1_5[13],stage1_4[41],stage1_3[43]}
   );
   gpc615_5 gpc44 (
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage0_4[46]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[11],stage1_5[14],stage1_4[42],stage1_3[44]}
   );
   gpc615_5 gpc45 (
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage0_4[47]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[12],stage1_5[15],stage1_4[43],stage1_3[45]}
   );
   gpc615_5 gpc46 (
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage0_4[48]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[13],stage1_5[16],stage1_4[44],stage1_3[46]}
   );
   gpc615_5 gpc47 (
      {stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage0_4[49]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[14],stage1_5[17],stage1_4[45],stage1_3[47]}
   );
   gpc615_5 gpc48 (
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage0_4[50]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[15],stage1_5[18],stage1_4[46],stage1_3[48]}
   );
   gpc615_5 gpc49 (
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage0_4[51]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[16],stage1_5[19],stage1_4[47],stage1_3[49]}
   );
   gpc615_5 gpc50 (
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage0_4[52]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[17],stage1_5[20],stage1_4[48],stage1_3[50]}
   );
   gpc615_5 gpc51 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[53]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[18],stage1_5[21],stage1_4[49],stage1_3[51]}
   );
   gpc615_5 gpc52 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[54]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[19],stage1_5[22],stage1_4[50],stage1_3[52]}
   );
   gpc615_5 gpc53 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[55]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[20],stage1_5[23],stage1_4[51],stage1_3[53]}
   );
   gpc615_5 gpc54 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[56]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[21],stage1_5[24],stage1_4[52],stage1_3[54]}
   );
   gpc615_5 gpc55 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[57]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[22],stage1_5[25],stage1_4[53],stage1_3[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[16],stage1_6[23],stage1_5[26],stage1_4[54]}
   );
   gpc606_5 gpc57 (
      {stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[17],stage1_6[24],stage1_5[27],stage1_4[55]}
   );
   gpc606_5 gpc58 (
      {stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[18],stage1_6[25],stage1_5[28],stage1_4[56]}
   );
   gpc606_5 gpc59 (
      {stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[19],stage1_6[26],stage1_5[29],stage1_4[57]}
   );
   gpc606_5 gpc60 (
      {stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[20],stage1_6[27],stage1_5[30],stage1_4[58]}
   );
   gpc606_5 gpc61 (
      {stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[21],stage1_6[28],stage1_5[31],stage1_4[59]}
   );
   gpc606_5 gpc62 (
      {stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[22],stage1_6[29],stage1_5[32],stage1_4[60]}
   );
   gpc606_5 gpc63 (
      {stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[23],stage1_6[30],stage1_5[33],stage1_4[61]}
   );
   gpc606_5 gpc64 (
      {stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[24],stage1_6[31],stage1_5[34],stage1_4[62]}
   );
   gpc606_5 gpc65 (
      {stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[25],stage1_6[32],stage1_5[35],stage1_4[63]}
   );
   gpc615_5 gpc66 (
      {stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122]},
      {stage0_5[96]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[26],stage1_6[33],stage1_5[36],stage1_4[64]}
   );
   gpc615_5 gpc67 (
      {stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_5[97]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[27],stage1_6[34],stage1_5[37],stage1_4[65]}
   );
   gpc615_5 gpc68 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102]},
      {stage0_6[72]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[12],stage1_7[28],stage1_6[35],stage1_5[38]}
   );
   gpc615_5 gpc69 (
      {stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_6[73]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[13],stage1_7[29],stage1_6[36],stage1_5[39]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[74]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[14],stage1_7[30],stage1_6[37],stage1_5[40]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[75]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[15],stage1_7[31],stage1_6[38],stage1_5[41]}
   );
   gpc623_5 gpc72 (
      {stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage0_7[24], stage0_7[25]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[16],stage1_7[32],stage1_6[39]}
   );
   gpc606_5 gpc73 (
      {stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[17],stage1_7[33]}
   );
   gpc606_5 gpc74 (
      {stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[18],stage1_7[34]}
   );
   gpc606_5 gpc75 (
      {stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[19],stage1_7[35]}
   );
   gpc606_5 gpc76 (
      {stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[20],stage1_7[36]}
   );
   gpc606_5 gpc77 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], stage0_7[54], stage0_7[55]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[21],stage1_7[37]}
   );
   gpc606_5 gpc78 (
      {stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[6],stage1_9[10],stage1_8[22],stage1_7[38]}
   );
   gpc606_5 gpc79 (
      {stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65], stage0_7[66], stage0_7[67]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[7],stage1_9[11],stage1_8[23],stage1_7[39]}
   );
   gpc606_5 gpc80 (
      {stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71], stage0_7[72], stage0_7[73]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[8],stage1_9[12],stage1_8[24],stage1_7[40]}
   );
   gpc606_5 gpc81 (
      {stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77], stage0_7[78], stage0_7[79]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[9],stage1_9[13],stage1_8[25],stage1_7[41]}
   );
   gpc606_5 gpc82 (
      {stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83], stage0_7[84], stage0_7[85]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[10],stage1_9[14],stage1_8[26],stage1_7[42]}
   );
   gpc606_5 gpc83 (
      {stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89], stage0_7[90], stage0_7[91]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[11],stage1_9[15],stage1_8[27],stage1_7[43]}
   );
   gpc606_5 gpc84 (
      {stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95], stage0_7[96], stage0_7[97]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[12],stage1_9[16],stage1_8[28],stage1_7[44]}
   );
   gpc615_5 gpc85 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[6]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[13],stage1_9[17],stage1_8[29],stage1_7[45]}
   );
   gpc606_5 gpc86 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[13],stage1_10[14],stage1_9[18],stage1_8[30]}
   );
   gpc606_5 gpc87 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[14],stage1_10[15],stage1_9[19],stage1_8[31]}
   );
   gpc606_5 gpc88 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[15],stage1_10[16],stage1_9[20],stage1_8[32]}
   );
   gpc606_5 gpc89 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[16],stage1_10[17],stage1_9[21],stage1_8[33]}
   );
   gpc606_5 gpc90 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[17],stage1_10[18],stage1_9[22],stage1_8[34]}
   );
   gpc606_5 gpc91 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[18],stage1_10[19],stage1_9[23],stage1_8[35]}
   );
   gpc606_5 gpc92 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[19],stage1_10[20],stage1_9[24],stage1_8[36]}
   );
   gpc606_5 gpc93 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[20],stage1_10[21],stage1_9[25],stage1_8[37]}
   );
   gpc606_5 gpc94 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[21],stage1_10[22],stage1_9[26],stage1_8[38]}
   );
   gpc606_5 gpc95 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[22],stage1_10[23],stage1_9[27],stage1_8[39]}
   );
   gpc606_5 gpc96 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[23],stage1_10[24],stage1_9[28],stage1_8[40]}
   );
   gpc606_5 gpc97 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[24],stage1_10[25],stage1_9[29],stage1_8[41]}
   );
   gpc606_5 gpc98 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[25],stage1_10[26],stage1_9[30],stage1_8[42]}
   );
   gpc606_5 gpc99 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[26],stage1_10[27],stage1_9[31],stage1_8[43]}
   );
   gpc606_5 gpc100 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[27],stage1_10[28],stage1_9[32],stage1_8[44]}
   );
   gpc606_5 gpc101 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[28],stage1_10[29],stage1_9[33],stage1_8[45]}
   );
   gpc606_5 gpc102 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[29],stage1_10[30],stage1_9[34],stage1_8[46]}
   );
   gpc615_5 gpc103 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82]},
      {stage0_10[102]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[17],stage1_11[30],stage1_10[31],stage1_9[35]}
   );
   gpc615_5 gpc104 (
      {stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_10[103]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[18],stage1_11[31],stage1_10[32],stage1_9[36]}
   );
   gpc615_5 gpc105 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_10[104]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[19],stage1_11[32],stage1_10[33],stage1_9[37]}
   );
   gpc615_5 gpc106 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_10[105]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[20],stage1_11[33],stage1_10[34],stage1_9[38]}
   );
   gpc615_5 gpc107 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102]},
      {stage0_10[106]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[21],stage1_11[34],stage1_10[35],stage1_9[39]}
   );
   gpc615_5 gpc108 (
      {stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_10[107]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[22],stage1_11[35],stage1_10[36],stage1_9[40]}
   );
   gpc615_5 gpc109 (
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112]},
      {stage0_11[36]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[6],stage1_12[23],stage1_11[36],stage1_10[37]}
   );
   gpc615_5 gpc110 (
      {stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117]},
      {stage0_11[37]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[7],stage1_12[24],stage1_11[37],stage1_10[38]}
   );
   gpc615_5 gpc111 (
      {stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121], stage0_10[122]},
      {stage0_11[38]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[8],stage1_12[25],stage1_11[38],stage1_10[39]}
   );
   gpc615_5 gpc112 (
      {stage0_10[123], stage0_10[124], stage0_10[125], stage0_10[126], stage0_10[127]},
      {stage0_11[39]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[9],stage1_12[26],stage1_11[39],stage1_10[40]}
   );
   gpc117_4 gpc113 (
      {stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage0_12[24]},
      {stage0_13[0]},
      {stage1_14[4],stage1_13[10],stage1_12[27],stage1_11[40]}
   );
   gpc117_4 gpc114 (
      {stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_12[25]},
      {stage0_13[1]},
      {stage1_14[5],stage1_13[11],stage1_12[28],stage1_11[41]}
   );
   gpc117_4 gpc115 (
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_12[26]},
      {stage0_13[2]},
      {stage1_14[6],stage1_13[12],stage1_12[29],stage1_11[42]}
   );
   gpc117_4 gpc116 (
      {stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67]},
      {stage0_12[27]},
      {stage0_13[3]},
      {stage1_14[7],stage1_13[13],stage1_12[30],stage1_11[43]}
   );
   gpc615_5 gpc117 (
      {stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71], stage0_11[72]},
      {stage0_12[28]},
      {stage0_13[4], stage0_13[5], stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9]},
      {stage1_15[0],stage1_14[8],stage1_13[14],stage1_12[31],stage1_11[44]}
   );
   gpc615_5 gpc118 (
      {stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage0_12[29]},
      {stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15]},
      {stage1_15[1],stage1_14[9],stage1_13[15],stage1_12[32],stage1_11[45]}
   );
   gpc615_5 gpc119 (
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82]},
      {stage0_12[30]},
      {stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21]},
      {stage1_15[2],stage1_14[10],stage1_13[16],stage1_12[33],stage1_11[46]}
   );
   gpc615_5 gpc120 (
      {stage0_11[83], stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87]},
      {stage0_12[31]},
      {stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27]},
      {stage1_15[3],stage1_14[11],stage1_13[17],stage1_12[34],stage1_11[47]}
   );
   gpc615_5 gpc121 (
      {stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91], stage0_11[92]},
      {stage0_12[32]},
      {stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33]},
      {stage1_15[4],stage1_14[12],stage1_13[18],stage1_12[35],stage1_11[48]}
   );
   gpc615_5 gpc122 (
      {stage0_11[93], stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97]},
      {stage0_12[33]},
      {stage0_13[34], stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39]},
      {stage1_15[5],stage1_14[13],stage1_13[19],stage1_12[36],stage1_11[49]}
   );
   gpc615_5 gpc123 (
      {stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102]},
      {stage0_12[34]},
      {stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45]},
      {stage1_15[6],stage1_14[14],stage1_13[20],stage1_12[37],stage1_11[50]}
   );
   gpc615_5 gpc124 (
      {stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage0_12[35]},
      {stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage1_15[7],stage1_14[15],stage1_13[21],stage1_12[38],stage1_11[51]}
   );
   gpc615_5 gpc125 (
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112]},
      {stage0_12[36]},
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57]},
      {stage1_15[8],stage1_14[16],stage1_13[22],stage1_12[39],stage1_11[52]}
   );
   gpc615_5 gpc126 (
      {stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117]},
      {stage0_12[37]},
      {stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63]},
      {stage1_15[9],stage1_14[17],stage1_13[23],stage1_12[40],stage1_11[53]}
   );
   gpc1406_5 gpc127 (
      {stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[10],stage1_14[18],stage1_13[24],stage1_12[41]}
   );
   gpc606_5 gpc128 (
      {stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49]},
      {stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9]},
      {stage1_16[1],stage1_15[11],stage1_14[19],stage1_13[25],stage1_12[42]}
   );
   gpc606_5 gpc129 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage1_16[2],stage1_15[12],stage1_14[20],stage1_13[26],stage1_12[43]}
   );
   gpc606_5 gpc130 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21]},
      {stage1_16[3],stage1_15[13],stage1_14[21],stage1_13[27],stage1_12[44]}
   );
   gpc606_5 gpc131 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage1_16[4],stage1_15[14],stage1_14[22],stage1_13[28],stage1_12[45]}
   );
   gpc606_5 gpc132 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33]},
      {stage1_16[5],stage1_15[15],stage1_14[23],stage1_13[29],stage1_12[46]}
   );
   gpc606_5 gpc133 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[34], stage0_14[35], stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39]},
      {stage1_16[6],stage1_15[16],stage1_14[24],stage1_13[30],stage1_12[47]}
   );
   gpc606_5 gpc134 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[40], stage0_14[41], stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45]},
      {stage1_16[7],stage1_15[17],stage1_14[25],stage1_13[31],stage1_12[48]}
   );
   gpc606_5 gpc135 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51]},
      {stage1_16[8],stage1_15[18],stage1_14[26],stage1_13[32],stage1_12[49]}
   );
   gpc606_5 gpc136 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57]},
      {stage1_16[9],stage1_15[19],stage1_14[27],stage1_13[33],stage1_12[50]}
   );
   gpc606_5 gpc137 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[58], stage0_14[59], stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63]},
      {stage1_16[10],stage1_15[20],stage1_14[28],stage1_13[34],stage1_12[51]}
   );
   gpc606_5 gpc138 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69]},
      {stage1_16[11],stage1_15[21],stage1_14[29],stage1_13[35],stage1_12[52]}
   );
   gpc606_5 gpc139 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75]},
      {stage1_16[12],stage1_15[22],stage1_14[30],stage1_13[36],stage1_12[53]}
   );
   gpc606_5 gpc140 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81]},
      {stage1_16[13],stage1_15[23],stage1_14[31],stage1_13[37],stage1_12[54]}
   );
   gpc606_5 gpc141 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[82], stage0_14[83], stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87]},
      {stage1_16[14],stage1_15[24],stage1_14[32],stage1_13[38],stage1_12[55]}
   );
   gpc606_5 gpc142 (
      {stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[15],stage1_15[25],stage1_14[33],stage1_13[39]}
   );
   gpc606_5 gpc143 (
      {stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[1],stage1_16[16],stage1_15[26],stage1_14[34],stage1_13[40]}
   );
   gpc606_5 gpc144 (
      {stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[2],stage1_16[17],stage1_15[27],stage1_14[35],stage1_13[41]}
   );
   gpc606_5 gpc145 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage1_17[3],stage1_16[18],stage1_15[28],stage1_14[36],stage1_13[42]}
   );
   gpc606_5 gpc146 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30]},
      {stage1_17[4],stage1_16[19],stage1_15[29],stage1_14[37],stage1_13[43]}
   );
   gpc615_5 gpc147 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98]},
      {stage0_14[88]},
      {stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36]},
      {stage1_17[5],stage1_16[20],stage1_15[30],stage1_14[38],stage1_13[44]}
   );
   gpc615_5 gpc148 (
      {stage0_13[99], stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103]},
      {stage0_14[89]},
      {stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41], stage0_15[42]},
      {stage1_17[6],stage1_16[21],stage1_15[31],stage1_14[39],stage1_13[45]}
   );
   gpc615_5 gpc149 (
      {stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108]},
      {stage0_14[90]},
      {stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47], stage0_15[48]},
      {stage1_17[7],stage1_16[22],stage1_15[32],stage1_14[40],stage1_13[46]}
   );
   gpc615_5 gpc150 (
      {stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_14[91]},
      {stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53], stage0_15[54]},
      {stage1_17[8],stage1_16[23],stage1_15[33],stage1_14[41],stage1_13[47]}
   );
   gpc615_5 gpc151 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118]},
      {stage0_14[92]},
      {stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59], stage0_15[60]},
      {stage1_17[9],stage1_16[24],stage1_15[34],stage1_14[42],stage1_13[48]}
   );
   gpc615_5 gpc152 (
      {stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_14[93]},
      {stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65], stage0_15[66]},
      {stage1_17[10],stage1_16[25],stage1_15[35],stage1_14[43],stage1_13[49]}
   );
   gpc615_5 gpc153 (
      {stage0_14[94], stage0_14[95], stage0_14[96], stage0_14[97], stage0_14[98]},
      {stage0_15[67]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[11],stage1_16[26],stage1_15[36],stage1_14[44]}
   );
   gpc615_5 gpc154 (
      {stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102], stage0_14[103]},
      {stage0_15[68]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[12],stage1_16[27],stage1_15[37],stage1_14[45]}
   );
   gpc615_5 gpc155 (
      {stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108]},
      {stage0_15[69]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[13],stage1_16[28],stage1_15[38],stage1_14[46]}
   );
   gpc1343_5 gpc156 (
      {stage0_15[70], stage0_15[71], stage0_15[72]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21]},
      {stage0_17[0], stage0_17[1], stage0_17[2]},
      {stage0_18[0]},
      {stage1_19[0],stage1_18[3],stage1_17[14],stage1_16[29],stage1_15[39]}
   );
   gpc606_5 gpc157 (
      {stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77], stage0_15[78]},
      {stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7], stage0_17[8]},
      {stage1_19[1],stage1_18[4],stage1_17[15],stage1_16[30],stage1_15[40]}
   );
   gpc606_5 gpc158 (
      {stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83], stage0_15[84]},
      {stage0_17[9], stage0_17[10], stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14]},
      {stage1_19[2],stage1_18[5],stage1_17[16],stage1_16[31],stage1_15[41]}
   );
   gpc606_5 gpc159 (
      {stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89], stage0_15[90]},
      {stage0_17[15], stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage1_19[3],stage1_18[6],stage1_17[17],stage1_16[32],stage1_15[42]}
   );
   gpc615_5 gpc160 (
      {stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage0_16[22]},
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26]},
      {stage1_19[4],stage1_18[7],stage1_17[18],stage1_16[33],stage1_15[43]}
   );
   gpc615_5 gpc161 (
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100]},
      {stage0_16[23]},
      {stage0_17[27], stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32]},
      {stage1_19[5],stage1_18[8],stage1_17[19],stage1_16[34],stage1_15[44]}
   );
   gpc615_5 gpc162 (
      {stage0_15[101], stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105]},
      {stage0_16[24]},
      {stage0_17[33], stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38]},
      {stage1_19[6],stage1_18[9],stage1_17[20],stage1_16[35],stage1_15[45]}
   );
   gpc606_5 gpc163 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5], stage0_18[6]},
      {stage1_20[0],stage1_19[7],stage1_18[10],stage1_17[21],stage1_16[36]}
   );
   gpc606_5 gpc164 (
      {stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36]},
      {stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11], stage0_18[12]},
      {stage1_20[1],stage1_19[8],stage1_18[11],stage1_17[22],stage1_16[37]}
   );
   gpc606_5 gpc165 (
      {stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17], stage0_18[18]},
      {stage1_20[2],stage1_19[9],stage1_18[12],stage1_17[23],stage1_16[38]}
   );
   gpc606_5 gpc166 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48]},
      {stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23], stage0_18[24]},
      {stage1_20[3],stage1_19[10],stage1_18[13],stage1_17[24],stage1_16[39]}
   );
   gpc606_5 gpc167 (
      {stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54]},
      {stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29], stage0_18[30]},
      {stage1_20[4],stage1_19[11],stage1_18[14],stage1_17[25],stage1_16[40]}
   );
   gpc606_5 gpc168 (
      {stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60]},
      {stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35], stage0_18[36]},
      {stage1_20[5],stage1_19[12],stage1_18[15],stage1_17[26],stage1_16[41]}
   );
   gpc606_5 gpc169 (
      {stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66]},
      {stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41], stage0_18[42]},
      {stage1_20[6],stage1_19[13],stage1_18[16],stage1_17[27],stage1_16[42]}
   );
   gpc606_5 gpc170 (
      {stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72]},
      {stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47], stage0_18[48]},
      {stage1_20[7],stage1_19[14],stage1_18[17],stage1_17[28],stage1_16[43]}
   );
   gpc606_5 gpc171 (
      {stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78]},
      {stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53], stage0_18[54]},
      {stage1_20[8],stage1_19[15],stage1_18[18],stage1_17[29],stage1_16[44]}
   );
   gpc606_5 gpc172 (
      {stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84]},
      {stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59], stage0_18[60]},
      {stage1_20[9],stage1_19[16],stage1_18[19],stage1_17[30],stage1_16[45]}
   );
   gpc606_5 gpc173 (
      {stage0_17[39], stage0_17[40], stage0_17[41], stage0_17[42], stage0_17[43], stage0_17[44]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[10],stage1_19[17],stage1_18[20],stage1_17[31]}
   );
   gpc606_5 gpc174 (
      {stage0_17[45], stage0_17[46], stage0_17[47], stage0_17[48], stage0_17[49], stage0_17[50]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[11],stage1_19[18],stage1_18[21],stage1_17[32]}
   );
   gpc606_5 gpc175 (
      {stage0_17[51], stage0_17[52], stage0_17[53], stage0_17[54], stage0_17[55], stage0_17[56]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[12],stage1_19[19],stage1_18[22],stage1_17[33]}
   );
   gpc606_5 gpc176 (
      {stage0_17[57], stage0_17[58], stage0_17[59], stage0_17[60], stage0_17[61], stage0_17[62]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[13],stage1_19[20],stage1_18[23],stage1_17[34]}
   );
   gpc606_5 gpc177 (
      {stage0_17[63], stage0_17[64], stage0_17[65], stage0_17[66], stage0_17[67], stage0_17[68]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[14],stage1_19[21],stage1_18[24],stage1_17[35]}
   );
   gpc606_5 gpc178 (
      {stage0_17[69], stage0_17[70], stage0_17[71], stage0_17[72], stage0_17[73], stage0_17[74]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[15],stage1_19[22],stage1_18[25],stage1_17[36]}
   );
   gpc606_5 gpc179 (
      {stage0_17[75], stage0_17[76], stage0_17[77], stage0_17[78], stage0_17[79], stage0_17[80]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[16],stage1_19[23],stage1_18[26],stage1_17[37]}
   );
   gpc606_5 gpc180 (
      {stage0_17[81], stage0_17[82], stage0_17[83], stage0_17[84], stage0_17[85], stage0_17[86]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[17],stage1_19[24],stage1_18[27],stage1_17[38]}
   );
   gpc606_5 gpc181 (
      {stage0_17[87], stage0_17[88], stage0_17[89], stage0_17[90], stage0_17[91], stage0_17[92]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[18],stage1_19[25],stage1_18[28],stage1_17[39]}
   );
   gpc615_5 gpc182 (
      {stage0_17[93], stage0_17[94], stage0_17[95], stage0_17[96], stage0_17[97]},
      {stage0_18[61]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[19],stage1_19[26],stage1_18[29],stage1_17[40]}
   );
   gpc615_5 gpc183 (
      {stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101], stage0_17[102]},
      {stage0_18[62]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[20],stage1_19[27],stage1_18[30],stage1_17[41]}
   );
   gpc606_5 gpc184 (
      {stage0_18[63], stage0_18[64], stage0_18[65], stage0_18[66], stage0_18[67], stage0_18[68]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[11],stage1_20[21],stage1_19[28],stage1_18[31]}
   );
   gpc606_5 gpc185 (
      {stage0_18[69], stage0_18[70], stage0_18[71], stage0_18[72], stage0_18[73], stage0_18[74]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[12],stage1_20[22],stage1_19[29],stage1_18[32]}
   );
   gpc606_5 gpc186 (
      {stage0_18[75], stage0_18[76], stage0_18[77], stage0_18[78], stage0_18[79], stage0_18[80]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[13],stage1_20[23],stage1_19[30],stage1_18[33]}
   );
   gpc606_5 gpc187 (
      {stage0_18[81], stage0_18[82], stage0_18[83], stage0_18[84], stage0_18[85], stage0_18[86]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[14],stage1_20[24],stage1_19[31],stage1_18[34]}
   );
   gpc606_5 gpc188 (
      {stage0_18[87], stage0_18[88], stage0_18[89], stage0_18[90], stage0_18[91], stage0_18[92]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[15],stage1_20[25],stage1_19[32],stage1_18[35]}
   );
   gpc606_5 gpc189 (
      {stage0_18[93], stage0_18[94], stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[16],stage1_20[26],stage1_19[33],stage1_18[36]}
   );
   gpc606_5 gpc190 (
      {stage0_18[99], stage0_18[100], stage0_18[101], stage0_18[102], stage0_18[103], stage0_18[104]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[17],stage1_20[27],stage1_19[34],stage1_18[37]}
   );
   gpc606_5 gpc191 (
      {stage0_18[105], stage0_18[106], stage0_18[107], stage0_18[108], stage0_18[109], stage0_18[110]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[18],stage1_20[28],stage1_19[35],stage1_18[38]}
   );
   gpc606_5 gpc192 (
      {stage0_18[111], stage0_18[112], stage0_18[113], stage0_18[114], stage0_18[115], stage0_18[116]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[19],stage1_20[29],stage1_19[36],stage1_18[39]}
   );
   gpc606_5 gpc193 (
      {stage0_18[117], stage0_18[118], stage0_18[119], stage0_18[120], stage0_18[121], stage0_18[122]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[20],stage1_20[30],stage1_19[37],stage1_18[40]}
   );
   gpc615_5 gpc194 (
      {stage0_18[123], stage0_18[124], stage0_18[125], stage0_18[126], stage0_18[127]},
      {stage0_19[66]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[21],stage1_20[31],stage1_19[38],stage1_18[41]}
   );
   gpc606_5 gpc195 (
      {stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71], stage0_19[72]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[11],stage1_21[22],stage1_20[32],stage1_19[39]}
   );
   gpc615_5 gpc196 (
      {stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage0_20[66]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[12],stage1_21[23],stage1_20[33],stage1_19[40]}
   );
   gpc615_5 gpc197 (
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82]},
      {stage0_20[67]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[13],stage1_21[24],stage1_20[34],stage1_19[41]}
   );
   gpc615_5 gpc198 (
      {stage0_19[83], stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87]},
      {stage0_20[68]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[14],stage1_21[25],stage1_20[35],stage1_19[42]}
   );
   gpc615_5 gpc199 (
      {stage0_19[88], stage0_19[89], stage0_19[90], stage0_19[91], stage0_19[92]},
      {stage0_20[69]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[15],stage1_21[26],stage1_20[36],stage1_19[43]}
   );
   gpc615_5 gpc200 (
      {stage0_19[93], stage0_19[94], stage0_19[95], stage0_19[96], stage0_19[97]},
      {stage0_20[70]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[16],stage1_21[27],stage1_20[37],stage1_19[44]}
   );
   gpc615_5 gpc201 (
      {stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101], stage0_19[102]},
      {stage0_20[71]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[17],stage1_21[28],stage1_20[38],stage1_19[45]}
   );
   gpc615_5 gpc202 (
      {stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage0_20[72]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[18],stage1_21[29],stage1_20[39],stage1_19[46]}
   );
   gpc615_5 gpc203 (
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112]},
      {stage0_20[73]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[19],stage1_21[30],stage1_20[40],stage1_19[47]}
   );
   gpc615_5 gpc204 (
      {stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117]},
      {stage0_20[74]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[20],stage1_21[31],stage1_20[41],stage1_19[48]}
   );
   gpc615_5 gpc205 (
      {stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122]},
      {stage0_20[75]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[21],stage1_21[32],stage1_20[42],stage1_19[49]}
   );
   gpc606_5 gpc206 (
      {stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[11],stage1_22[22],stage1_21[33],stage1_20[43]}
   );
   gpc606_5 gpc207 (
      {stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[12],stage1_22[23],stage1_21[34],stage1_20[44]}
   );
   gpc606_5 gpc208 (
      {stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[13],stage1_22[24],stage1_21[35],stage1_20[45]}
   );
   gpc615_5 gpc209 (
      {stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_21[66]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[14],stage1_22[25],stage1_21[36],stage1_20[46]}
   );
   gpc615_5 gpc210 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103]},
      {stage0_21[67]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[15],stage1_22[26],stage1_21[37],stage1_20[47]}
   );
   gpc606_5 gpc211 (
      {stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72], stage0_21[73]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[5],stage1_23[16],stage1_22[27],stage1_21[38]}
   );
   gpc606_5 gpc212 (
      {stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78], stage0_21[79]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[6],stage1_23[17],stage1_22[28],stage1_21[39]}
   );
   gpc606_5 gpc213 (
      {stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84], stage0_21[85]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[7],stage1_23[18],stage1_22[29],stage1_21[40]}
   );
   gpc615_5 gpc214 (
      {stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_22[30]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[8],stage1_23[19],stage1_22[30],stage1_21[41]}
   );
   gpc615_5 gpc215 (
      {stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_22[31]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[9],stage1_23[20],stage1_22[31],stage1_21[42]}
   );
   gpc615_5 gpc216 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100]},
      {stage0_22[32]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[10],stage1_23[21],stage1_22[32],stage1_21[43]}
   );
   gpc615_5 gpc217 (
      {stage0_21[101], stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105]},
      {stage0_22[33]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[11],stage1_23[22],stage1_22[33],stage1_21[44]}
   );
   gpc615_5 gpc218 (
      {stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109], stage0_21[110]},
      {stage0_22[34]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[12],stage1_23[23],stage1_22[34],stage1_21[45]}
   );
   gpc615_5 gpc219 (
      {stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage0_22[35]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[13],stage1_23[24],stage1_22[35],stage1_21[46]}
   );
   gpc615_5 gpc220 (
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120]},
      {stage0_22[36]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[14],stage1_23[25],stage1_22[36],stage1_21[47]}
   );
   gpc606_5 gpc221 (
      {stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[10],stage1_24[15],stage1_23[26],stage1_22[37]}
   );
   gpc606_5 gpc222 (
      {stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[11],stage1_24[16],stage1_23[27],stage1_22[38]}
   );
   gpc606_5 gpc223 (
      {stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[12],stage1_24[17],stage1_23[28],stage1_22[39]}
   );
   gpc606_5 gpc224 (
      {stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[13],stage1_24[18],stage1_23[29],stage1_22[40]}
   );
   gpc606_5 gpc225 (
      {stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[14],stage1_24[19],stage1_23[30],stage1_22[41]}
   );
   gpc606_5 gpc226 (
      {stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[15],stage1_24[20],stage1_23[31],stage1_22[42]}
   );
   gpc606_5 gpc227 (
      {stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[16],stage1_24[21],stage1_23[32],stage1_22[43]}
   );
   gpc606_5 gpc228 (
      {stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[17],stage1_24[22],stage1_23[33],stage1_22[44]}
   );
   gpc606_5 gpc229 (
      {stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[18],stage1_24[23],stage1_23[34],stage1_22[45]}
   );
   gpc615_5 gpc230 (
      {stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage0_23[60]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[19],stage1_24[24],stage1_23[35],stage1_22[46]}
   );
   gpc615_5 gpc231 (
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100]},
      {stage0_23[61]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[20],stage1_24[25],stage1_23[36],stage1_22[47]}
   );
   gpc615_5 gpc232 (
      {stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105]},
      {stage0_23[62]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[21],stage1_24[26],stage1_23[37],stage1_22[48]}
   );
   gpc606_5 gpc233 (
      {stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[12],stage1_25[22],stage1_24[27],stage1_23[38]}
   );
   gpc606_5 gpc234 (
      {stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[13],stage1_25[23],stage1_24[28],stage1_23[39]}
   );
   gpc606_5 gpc235 (
      {stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[14],stage1_25[24],stage1_24[29],stage1_23[40]}
   );
   gpc606_5 gpc236 (
      {stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[15],stage1_25[25],stage1_24[30],stage1_23[41]}
   );
   gpc606_5 gpc237 (
      {stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[16],stage1_25[26],stage1_24[31],stage1_23[42]}
   );
   gpc606_5 gpc238 (
      {stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[17],stage1_25[27],stage1_24[32],stage1_23[43]}
   );
   gpc606_5 gpc239 (
      {stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[18],stage1_25[28],stage1_24[33],stage1_23[44]}
   );
   gpc606_5 gpc240 (
      {stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[19],stage1_25[29],stage1_24[34],stage1_23[45]}
   );
   gpc606_5 gpc241 (
      {stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[20],stage1_25[30],stage1_24[35],stage1_23[46]}
   );
   gpc615_5 gpc242 (
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121]},
      {stage0_24[72]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[21],stage1_25[31],stage1_24[36],stage1_23[47]}
   );
   gpc606_5 gpc243 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[22],stage1_25[32],stage1_24[37]}
   );
   gpc606_5 gpc244 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[23],stage1_25[33],stage1_24[38]}
   );
   gpc606_5 gpc245 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[24],stage1_25[34],stage1_24[39]}
   );
   gpc606_5 gpc246 (
      {stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[25],stage1_25[35],stage1_24[40]}
   );
   gpc606_5 gpc247 (
      {stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[26],stage1_25[36],stage1_24[41]}
   );
   gpc606_5 gpc248 (
      {stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[27],stage1_25[37],stage1_24[42]}
   );
   gpc606_5 gpc249 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[6],stage1_27[16],stage1_26[28],stage1_25[38]}
   );
   gpc606_5 gpc250 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[7],stage1_27[17],stage1_26[29],stage1_25[39]}
   );
   gpc606_5 gpc251 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[8],stage1_27[18],stage1_26[30],stage1_25[40]}
   );
   gpc606_5 gpc252 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[9],stage1_27[19],stage1_26[31],stage1_25[41]}
   );
   gpc606_5 gpc253 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[10],stage1_27[20],stage1_26[32],stage1_25[42]}
   );
   gpc606_5 gpc254 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[11],stage1_27[21],stage1_26[33],stage1_25[43]}
   );
   gpc606_5 gpc255 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[12],stage1_27[22],stage1_26[34],stage1_25[44]}
   );
   gpc606_5 gpc256 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[13],stage1_27[23],stage1_26[35],stage1_25[45]}
   );
   gpc606_5 gpc257 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[14],stage1_27[24],stage1_26[36],stage1_25[46]}
   );
   gpc1163_5 gpc258 (
      {stage0_26[36], stage0_26[37], stage0_26[38]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage0_28[0]},
      {stage0_29[0]},
      {stage1_30[0],stage1_29[9],stage1_28[15],stage1_27[25],stage1_26[37]}
   );
   gpc1163_5 gpc259 (
      {stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage0_28[1]},
      {stage0_29[1]},
      {stage1_30[1],stage1_29[10],stage1_28[16],stage1_27[26],stage1_26[38]}
   );
   gpc1163_5 gpc260 (
      {stage0_26[42], stage0_26[43], stage0_26[44]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage0_28[2]},
      {stage0_29[2]},
      {stage1_30[2],stage1_29[11],stage1_28[17],stage1_27[27],stage1_26[39]}
   );
   gpc1163_5 gpc261 (
      {stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage0_28[3]},
      {stage0_29[3]},
      {stage1_30[3],stage1_29[12],stage1_28[18],stage1_27[28],stage1_26[40]}
   );
   gpc1163_5 gpc262 (
      {stage0_26[48], stage0_26[49], stage0_26[50]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage0_28[4]},
      {stage0_29[4]},
      {stage1_30[4],stage1_29[13],stage1_28[19],stage1_27[29],stage1_26[41]}
   );
   gpc207_4 gpc263 (
      {stage0_26[51], stage0_26[52], stage0_26[53], stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57]},
      {stage0_28[5], stage0_28[6]},
      {stage1_29[14],stage1_28[20],stage1_27[30],stage1_26[42]}
   );
   gpc606_5 gpc264 (
      {stage0_26[58], stage0_26[59], stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63]},
      {stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12]},
      {stage1_30[5],stage1_29[15],stage1_28[21],stage1_27[31],stage1_26[43]}
   );
   gpc606_5 gpc265 (
      {stage0_26[64], stage0_26[65], stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69]},
      {stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18]},
      {stage1_30[6],stage1_29[16],stage1_28[22],stage1_27[32],stage1_26[44]}
   );
   gpc606_5 gpc266 (
      {stage0_26[70], stage0_26[71], stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75]},
      {stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24]},
      {stage1_30[7],stage1_29[17],stage1_28[23],stage1_27[33],stage1_26[45]}
   );
   gpc606_5 gpc267 (
      {stage0_26[76], stage0_26[77], stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81]},
      {stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29], stage0_28[30]},
      {stage1_30[8],stage1_29[18],stage1_28[24],stage1_27[34],stage1_26[46]}
   );
   gpc606_5 gpc268 (
      {stage0_26[82], stage0_26[83], stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87]},
      {stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36]},
      {stage1_30[9],stage1_29[19],stage1_28[25],stage1_27[35],stage1_26[47]}
   );
   gpc615_5 gpc269 (
      {stage0_26[88], stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92]},
      {stage0_27[84]},
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage1_30[10],stage1_29[20],stage1_28[26],stage1_27[36],stage1_26[48]}
   );
   gpc2135_5 gpc270 (
      {stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage0_28[43], stage0_28[44], stage0_28[45]},
      {stage0_29[5]},
      {stage0_30[0], stage0_30[1]},
      {stage1_31[0],stage1_30[11],stage1_29[21],stage1_28[27],stage1_27[37]}
   );
   gpc606_5 gpc271 (
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[12],stage1_29[22],stage1_28[28],stage1_27[38]}
   );
   gpc606_5 gpc272 (
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[13],stage1_29[23],stage1_28[29],stage1_27[39]}
   );
   gpc606_5 gpc273 (
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[14],stage1_29[24],stage1_28[30],stage1_27[40]}
   );
   gpc606_5 gpc274 (
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[15],stage1_29[25],stage1_28[31],stage1_27[41]}
   );
   gpc606_5 gpc275 (
      {stage0_28[46], stage0_28[47], stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51]},
      {stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6], stage0_30[7]},
      {stage1_32[0],stage1_31[5],stage1_30[16],stage1_29[26],stage1_28[32]}
   );
   gpc606_5 gpc276 (
      {stage0_28[52], stage0_28[53], stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57]},
      {stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12], stage0_30[13]},
      {stage1_32[1],stage1_31[6],stage1_30[17],stage1_29[27],stage1_28[33]}
   );
   gpc606_5 gpc277 (
      {stage0_28[58], stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63]},
      {stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18], stage0_30[19]},
      {stage1_32[2],stage1_31[7],stage1_30[18],stage1_29[28],stage1_28[34]}
   );
   gpc606_5 gpc278 (
      {stage0_28[64], stage0_28[65], stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69]},
      {stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24], stage0_30[25]},
      {stage1_32[3],stage1_31[8],stage1_30[19],stage1_29[29],stage1_28[35]}
   );
   gpc606_5 gpc279 (
      {stage0_28[70], stage0_28[71], stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75]},
      {stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30], stage0_30[31]},
      {stage1_32[4],stage1_31[9],stage1_30[20],stage1_29[30],stage1_28[36]}
   );
   gpc606_5 gpc280 (
      {stage0_28[76], stage0_28[77], stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81]},
      {stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36], stage0_30[37]},
      {stage1_32[5],stage1_31[10],stage1_30[21],stage1_29[31],stage1_28[37]}
   );
   gpc606_5 gpc281 (
      {stage0_28[82], stage0_28[83], stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87]},
      {stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42], stage0_30[43]},
      {stage1_32[6],stage1_31[11],stage1_30[22],stage1_29[32],stage1_28[38]}
   );
   gpc606_5 gpc282 (
      {stage0_28[88], stage0_28[89], stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93]},
      {stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48], stage0_30[49]},
      {stage1_32[7],stage1_31[12],stage1_30[23],stage1_29[33],stage1_28[39]}
   );
   gpc606_5 gpc283 (
      {stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99]},
      {stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54], stage0_30[55]},
      {stage1_32[8],stage1_31[13],stage1_30[24],stage1_29[34],stage1_28[40]}
   );
   gpc606_5 gpc284 (
      {stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105]},
      {stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60], stage0_30[61]},
      {stage1_32[9],stage1_31[14],stage1_30[25],stage1_29[35],stage1_28[41]}
   );
   gpc615_5 gpc285 (
      {stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109], stage0_28[110]},
      {stage0_29[30]},
      {stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66], stage0_30[67]},
      {stage1_32[10],stage1_31[15],stage1_30[26],stage1_29[36],stage1_28[42]}
   );
   gpc615_5 gpc286 (
      {stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_29[31]},
      {stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72], stage0_30[73]},
      {stage1_32[11],stage1_31[16],stage1_30[27],stage1_29[37],stage1_28[43]}
   );
   gpc615_5 gpc287 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_29[32]},
      {stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78], stage0_30[79]},
      {stage1_32[12],stage1_31[17],stage1_30[28],stage1_29[38],stage1_28[44]}
   );
   gpc615_5 gpc288 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_29[33]},
      {stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84], stage0_30[85]},
      {stage1_32[13],stage1_31[18],stage1_30[29],stage1_29[39],stage1_28[45]}
   );
   gpc135_4 gpc289 (
      {stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37], stage0_29[38]},
      {stage0_30[86], stage0_30[87], stage0_30[88]},
      {stage0_31[0]},
      {stage1_32[14],stage1_31[19],stage1_30[30],stage1_29[40]}
   );
   gpc606_5 gpc290 (
      {stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43], stage0_29[44]},
      {stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6]},
      {stage1_33[0],stage1_32[15],stage1_31[20],stage1_30[31],stage1_29[41]}
   );
   gpc606_5 gpc291 (
      {stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49], stage0_29[50]},
      {stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12]},
      {stage1_33[1],stage1_32[16],stage1_31[21],stage1_30[32],stage1_29[42]}
   );
   gpc606_5 gpc292 (
      {stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55], stage0_29[56]},
      {stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18]},
      {stage1_33[2],stage1_32[17],stage1_31[22],stage1_30[33],stage1_29[43]}
   );
   gpc606_5 gpc293 (
      {stage0_29[57], stage0_29[58], stage0_29[59], stage0_29[60], stage0_29[61], stage0_29[62]},
      {stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24]},
      {stage1_33[3],stage1_32[18],stage1_31[23],stage1_30[34],stage1_29[44]}
   );
   gpc606_5 gpc294 (
      {stage0_29[63], stage0_29[64], stage0_29[65], stage0_29[66], stage0_29[67], stage0_29[68]},
      {stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30]},
      {stage1_33[4],stage1_32[19],stage1_31[24],stage1_30[35],stage1_29[45]}
   );
   gpc606_5 gpc295 (
      {stage0_29[69], stage0_29[70], stage0_29[71], stage0_29[72], stage0_29[73], stage0_29[74]},
      {stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36]},
      {stage1_33[5],stage1_32[20],stage1_31[25],stage1_30[36],stage1_29[46]}
   );
   gpc606_5 gpc296 (
      {stage0_29[75], stage0_29[76], stage0_29[77], stage0_29[78], stage0_29[79], stage0_29[80]},
      {stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42]},
      {stage1_33[6],stage1_32[21],stage1_31[26],stage1_30[37],stage1_29[47]}
   );
   gpc606_5 gpc297 (
      {stage0_29[81], stage0_29[82], stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86]},
      {stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48]},
      {stage1_33[7],stage1_32[22],stage1_31[27],stage1_30[38],stage1_29[48]}
   );
   gpc606_5 gpc298 (
      {stage0_29[87], stage0_29[88], stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92]},
      {stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54]},
      {stage1_33[8],stage1_32[23],stage1_31[28],stage1_30[39],stage1_29[49]}
   );
   gpc606_5 gpc299 (
      {stage0_29[93], stage0_29[94], stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98]},
      {stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60]},
      {stage1_33[9],stage1_32[24],stage1_31[29],stage1_30[40],stage1_29[50]}
   );
   gpc615_5 gpc300 (
      {stage0_30[89], stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93]},
      {stage0_31[61]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[10],stage1_32[25],stage1_31[30],stage1_30[41]}
   );
   gpc615_5 gpc301 (
      {stage0_30[94], stage0_30[95], stage0_30[96], stage0_30[97], stage0_30[98]},
      {stage0_31[62]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[11],stage1_32[26],stage1_31[31],stage1_30[42]}
   );
   gpc2116_5 gpc302 (
      {stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67], stage0_31[68]},
      {stage0_32[12]},
      {stage0_33[0]},
      {stage0_34[0], stage0_34[1]},
      {stage1_35[0],stage1_34[2],stage1_33[12],stage1_32[27],stage1_31[32]}
   );
   gpc615_5 gpc303 (
      {stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage0_32[13]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[1],stage1_34[3],stage1_33[13],stage1_32[28],stage1_31[33]}
   );
   gpc615_5 gpc304 (
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78]},
      {stage0_32[14]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[2],stage1_34[4],stage1_33[14],stage1_32[29],stage1_31[34]}
   );
   gpc615_5 gpc305 (
      {stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage0_32[15]},
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage1_35[3],stage1_34[5],stage1_33[15],stage1_32[30],stage1_31[35]}
   );
   gpc615_5 gpc306 (
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88]},
      {stage0_32[16]},
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage1_35[4],stage1_34[6],stage1_33[16],stage1_32[31],stage1_31[36]}
   );
   gpc615_5 gpc307 (
      {stage0_31[89], stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93]},
      {stage0_32[17]},
      {stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29], stage0_33[30]},
      {stage1_35[5],stage1_34[7],stage1_33[17],stage1_32[32],stage1_31[37]}
   );
   gpc615_5 gpc308 (
      {stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97], stage0_31[98]},
      {stage0_32[18]},
      {stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35], stage0_33[36]},
      {stage1_35[6],stage1_34[8],stage1_33[18],stage1_32[33],stage1_31[38]}
   );
   gpc615_5 gpc309 (
      {stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage0_32[19]},
      {stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41], stage0_33[42]},
      {stage1_35[7],stage1_34[9],stage1_33[19],stage1_32[34],stage1_31[39]}
   );
   gpc615_5 gpc310 (
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108]},
      {stage0_32[20]},
      {stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47], stage0_33[48]},
      {stage1_35[8],stage1_34[10],stage1_33[20],stage1_32[35],stage1_31[40]}
   );
   gpc606_5 gpc311 (
      {stage0_32[21], stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26]},
      {stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5], stage0_34[6], stage0_34[7]},
      {stage1_36[0],stage1_35[9],stage1_34[11],stage1_33[21],stage1_32[36]}
   );
   gpc606_5 gpc312 (
      {stage0_32[27], stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32]},
      {stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11], stage0_34[12], stage0_34[13]},
      {stage1_36[1],stage1_35[10],stage1_34[12],stage1_33[22],stage1_32[37]}
   );
   gpc606_5 gpc313 (
      {stage0_32[33], stage0_32[34], stage0_32[35], stage0_32[36], stage0_32[37], stage0_32[38]},
      {stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17], stage0_34[18], stage0_34[19]},
      {stage1_36[2],stage1_35[11],stage1_34[13],stage1_33[23],stage1_32[38]}
   );
   gpc606_5 gpc314 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23], stage0_34[24], stage0_34[25]},
      {stage1_36[3],stage1_35[12],stage1_34[14],stage1_33[24],stage1_32[39]}
   );
   gpc606_5 gpc315 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29], stage0_34[30], stage0_34[31]},
      {stage1_36[4],stage1_35[13],stage1_34[15],stage1_33[25],stage1_32[40]}
   );
   gpc606_5 gpc316 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35], stage0_34[36], stage0_34[37]},
      {stage1_36[5],stage1_35[14],stage1_34[16],stage1_33[26],stage1_32[41]}
   );
   gpc606_5 gpc317 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41], stage0_34[42], stage0_34[43]},
      {stage1_36[6],stage1_35[15],stage1_34[17],stage1_33[27],stage1_32[42]}
   );
   gpc606_5 gpc318 (
      {stage0_32[63], stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47], stage0_34[48], stage0_34[49]},
      {stage1_36[7],stage1_35[16],stage1_34[18],stage1_33[28],stage1_32[43]}
   );
   gpc606_5 gpc319 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73], stage0_32[74]},
      {stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53], stage0_34[54], stage0_34[55]},
      {stage1_36[8],stage1_35[17],stage1_34[19],stage1_33[29],stage1_32[44]}
   );
   gpc606_5 gpc320 (
      {stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78], stage0_32[79], stage0_32[80]},
      {stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59], stage0_34[60], stage0_34[61]},
      {stage1_36[9],stage1_35[18],stage1_34[20],stage1_33[30],stage1_32[45]}
   );
   gpc606_5 gpc321 (
      {stage0_32[81], stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86]},
      {stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65], stage0_34[66], stage0_34[67]},
      {stage1_36[10],stage1_35[19],stage1_34[21],stage1_33[31],stage1_32[46]}
   );
   gpc606_5 gpc322 (
      {stage0_32[87], stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92]},
      {stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71], stage0_34[72], stage0_34[73]},
      {stage1_36[11],stage1_35[20],stage1_34[22],stage1_33[32],stage1_32[47]}
   );
   gpc606_5 gpc323 (
      {stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53], stage0_33[54]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[12],stage1_35[21],stage1_34[23],stage1_33[33]}
   );
   gpc606_5 gpc324 (
      {stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59], stage0_33[60]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[13],stage1_35[22],stage1_34[24],stage1_33[34]}
   );
   gpc606_5 gpc325 (
      {stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65], stage0_33[66]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[14],stage1_35[23],stage1_34[25],stage1_33[35]}
   );
   gpc606_5 gpc326 (
      {stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71], stage0_33[72]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[15],stage1_35[24],stage1_34[26],stage1_33[36]}
   );
   gpc606_5 gpc327 (
      {stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77], stage0_33[78]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[16],stage1_35[25],stage1_34[27],stage1_33[37]}
   );
   gpc615_5 gpc328 (
      {stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage0_34[74]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[17],stage1_35[26],stage1_34[28],stage1_33[38]}
   );
   gpc615_5 gpc329 (
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88]},
      {stage0_34[75]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[18],stage1_35[27],stage1_34[29],stage1_33[39]}
   );
   gpc615_5 gpc330 (
      {stage0_33[89], stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93]},
      {stage0_34[76]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[19],stage1_35[28],stage1_34[30],stage1_33[40]}
   );
   gpc615_5 gpc331 (
      {stage0_33[94], stage0_33[95], stage0_33[96], stage0_33[97], stage0_33[98]},
      {stage0_34[77]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[20],stage1_35[29],stage1_34[31],stage1_33[41]}
   );
   gpc615_5 gpc332 (
      {stage0_33[99], stage0_33[100], stage0_33[101], stage0_33[102], stage0_33[103]},
      {stage0_34[78]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[21],stage1_35[30],stage1_34[32],stage1_33[42]}
   );
   gpc615_5 gpc333 (
      {stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107], stage0_33[108]},
      {stage0_34[79]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[22],stage1_35[31],stage1_34[33],stage1_33[43]}
   );
   gpc606_5 gpc334 (
      {stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83], stage0_34[84], stage0_34[85]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[11],stage1_36[23],stage1_35[32],stage1_34[34]}
   );
   gpc606_5 gpc335 (
      {stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89], stage0_34[90], stage0_34[91]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[12],stage1_36[24],stage1_35[33],stage1_34[35]}
   );
   gpc615_5 gpc336 (
      {stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95], stage0_34[96]},
      {stage0_35[66]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[13],stage1_36[25],stage1_35[34],stage1_34[36]}
   );
   gpc615_5 gpc337 (
      {stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage0_36[18]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[3],stage1_37[14],stage1_36[26],stage1_35[35]}
   );
   gpc615_5 gpc338 (
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76]},
      {stage0_36[19]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[4],stage1_37[15],stage1_36[27],stage1_35[36]}
   );
   gpc615_5 gpc339 (
      {stage0_35[77], stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81]},
      {stage0_36[20]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[5],stage1_37[16],stage1_36[28],stage1_35[37]}
   );
   gpc615_5 gpc340 (
      {stage0_35[82], stage0_35[83], stage0_35[84], stage0_35[85], stage0_35[86]},
      {stage0_36[21]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[6],stage1_37[17],stage1_36[29],stage1_35[38]}
   );
   gpc615_5 gpc341 (
      {stage0_35[87], stage0_35[88], stage0_35[89], stage0_35[90], stage0_35[91]},
      {stage0_36[22]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[7],stage1_37[18],stage1_36[30],stage1_35[39]}
   );
   gpc615_5 gpc342 (
      {stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95], stage0_35[96]},
      {stage0_36[23]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[8],stage1_37[19],stage1_36[31],stage1_35[40]}
   );
   gpc615_5 gpc343 (
      {stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage0_36[24]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[9],stage1_37[20],stage1_36[32],stage1_35[41]}
   );
   gpc615_5 gpc344 (
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106]},
      {stage0_36[25]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[10],stage1_37[21],stage1_36[33],stage1_35[42]}
   );
   gpc615_5 gpc345 (
      {stage0_35[107], stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111]},
      {stage0_36[26]},
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage1_39[8],stage1_38[11],stage1_37[22],stage1_36[34],stage1_35[43]}
   );
   gpc615_5 gpc346 (
      {stage0_35[112], stage0_35[113], stage0_35[114], stage0_35[115], stage0_35[116]},
      {stage0_36[27]},
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage1_39[9],stage1_38[12],stage1_37[23],stage1_36[35],stage1_35[44]}
   );
   gpc615_5 gpc347 (
      {stage0_35[117], stage0_35[118], stage0_35[119], stage0_35[120], stage0_35[121]},
      {stage0_36[28]},
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage1_39[10],stage1_38[13],stage1_37[24],stage1_36[36],stage1_35[45]}
   );
   gpc615_5 gpc348 (
      {stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125], stage0_35[126]},
      {stage0_36[29]},
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage1_39[11],stage1_38[14],stage1_37[25],stage1_36[37],stage1_35[46]}
   );
   gpc606_5 gpc349 (
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[12],stage1_38[15],stage1_37[26],stage1_36[38]}
   );
   gpc606_5 gpc350 (
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[13],stage1_38[16],stage1_37[27],stage1_36[39]}
   );
   gpc606_5 gpc351 (
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[14],stage1_38[17],stage1_37[28],stage1_36[40]}
   );
   gpc606_5 gpc352 (
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[15],stage1_38[18],stage1_37[29],stage1_36[41]}
   );
   gpc606_5 gpc353 (
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[16],stage1_38[19],stage1_37[30],stage1_36[42]}
   );
   gpc606_5 gpc354 (
      {stage0_36[60], stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[17],stage1_38[20],stage1_37[31],stage1_36[43]}
   );
   gpc606_5 gpc355 (
      {stage0_36[66], stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[18],stage1_38[21],stage1_37[32],stage1_36[44]}
   );
   gpc606_5 gpc356 (
      {stage0_36[72], stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[19],stage1_38[22],stage1_37[33],stage1_36[45]}
   );
   gpc606_5 gpc357 (
      {stage0_36[78], stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[20],stage1_38[23],stage1_37[34],stage1_36[46]}
   );
   gpc606_5 gpc358 (
      {stage0_36[84], stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[21],stage1_38[24],stage1_37[35],stage1_36[47]}
   );
   gpc606_5 gpc359 (
      {stage0_36[90], stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[22],stage1_38[25],stage1_37[36],stage1_36[48]}
   );
   gpc606_5 gpc360 (
      {stage0_36[96], stage0_36[97], stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[23],stage1_38[26],stage1_37[37],stage1_36[49]}
   );
   gpc606_5 gpc361 (
      {stage0_36[102], stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[24],stage1_38[27],stage1_37[38],stage1_36[50]}
   );
   gpc606_5 gpc362 (
      {stage0_36[108], stage0_36[109], stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[25],stage1_38[28],stage1_37[39],stage1_36[51]}
   );
   gpc606_5 gpc363 (
      {stage0_36[114], stage0_36[115], stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[26],stage1_38[29],stage1_37[40],stage1_36[52]}
   );
   gpc615_5 gpc364 (
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94]},
      {stage0_39[0]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[0],stage1_40[15],stage1_39[27],stage1_38[30]}
   );
   gpc615_5 gpc365 (
      {stage0_38[95], stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99]},
      {stage0_39[1]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[1],stage1_40[16],stage1_39[28],stage1_38[31]}
   );
   gpc615_5 gpc366 (
      {stage0_38[100], stage0_38[101], stage0_38[102], stage0_38[103], stage0_38[104]},
      {stage0_39[2]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[2],stage1_40[17],stage1_39[29],stage1_38[32]}
   );
   gpc615_5 gpc367 (
      {stage0_38[105], stage0_38[106], stage0_38[107], stage0_38[108], stage0_38[109]},
      {stage0_39[3]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[3],stage1_40[18],stage1_39[30],stage1_38[33]}
   );
   gpc615_5 gpc368 (
      {stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113], stage0_38[114]},
      {stage0_39[4]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[4],stage1_40[19],stage1_39[31],stage1_38[34]}
   );
   gpc615_5 gpc369 (
      {stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage0_39[5]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[5],stage1_40[20],stage1_39[32],stage1_38[35]}
   );
   gpc606_5 gpc370 (
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[6],stage1_41[6],stage1_40[21],stage1_39[33]}
   );
   gpc606_5 gpc371 (
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[7],stage1_41[7],stage1_40[22],stage1_39[34]}
   );
   gpc615_5 gpc372 (
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22]},
      {stage0_40[36]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[8],stage1_41[8],stage1_40[23],stage1_39[35]}
   );
   gpc615_5 gpc373 (
      {stage0_39[23], stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27]},
      {stage0_40[37]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[9],stage1_41[9],stage1_40[24],stage1_39[36]}
   );
   gpc615_5 gpc374 (
      {stage0_39[28], stage0_39[29], stage0_39[30], stage0_39[31], stage0_39[32]},
      {stage0_40[38]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[10],stage1_41[10],stage1_40[25],stage1_39[37]}
   );
   gpc615_5 gpc375 (
      {stage0_39[33], stage0_39[34], stage0_39[35], stage0_39[36], stage0_39[37]},
      {stage0_40[39]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[11],stage1_41[11],stage1_40[26],stage1_39[38]}
   );
   gpc615_5 gpc376 (
      {stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41], stage0_39[42]},
      {stage0_40[40]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[12],stage1_41[12],stage1_40[27],stage1_39[39]}
   );
   gpc615_5 gpc377 (
      {stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage0_40[41]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[13],stage1_41[13],stage1_40[28],stage1_39[40]}
   );
   gpc615_5 gpc378 (
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52]},
      {stage0_40[42]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[14],stage1_41[14],stage1_40[29],stage1_39[41]}
   );
   gpc615_5 gpc379 (
      {stage0_39[53], stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57]},
      {stage0_40[43]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[15],stage1_41[15],stage1_40[30],stage1_39[42]}
   );
   gpc615_5 gpc380 (
      {stage0_39[58], stage0_39[59], stage0_39[60], stage0_39[61], stage0_39[62]},
      {stage0_40[44]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[16],stage1_41[16],stage1_40[31],stage1_39[43]}
   );
   gpc615_5 gpc381 (
      {stage0_39[63], stage0_39[64], stage0_39[65], stage0_39[66], stage0_39[67]},
      {stage0_40[45]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[17],stage1_41[17],stage1_40[32],stage1_39[44]}
   );
   gpc615_5 gpc382 (
      {stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71], stage0_39[72]},
      {stage0_40[46]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[18],stage1_41[18],stage1_40[33],stage1_39[45]}
   );
   gpc615_5 gpc383 (
      {stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage0_40[47]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[19],stage1_41[19],stage1_40[34],stage1_39[46]}
   );
   gpc615_5 gpc384 (
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82]},
      {stage0_40[48]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[20],stage1_41[20],stage1_40[35],stage1_39[47]}
   );
   gpc1163_5 gpc385 (
      {stage0_40[49], stage0_40[50], stage0_40[51]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage0_42[0]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[15],stage1_42[21],stage1_41[21],stage1_40[36]}
   );
   gpc606_5 gpc386 (
      {stage0_40[52], stage0_40[53], stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57]},
      {stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5], stage0_42[6]},
      {stage1_44[1],stage1_43[16],stage1_42[22],stage1_41[22],stage1_40[37]}
   );
   gpc606_5 gpc387 (
      {stage0_40[58], stage0_40[59], stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63]},
      {stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11], stage0_42[12]},
      {stage1_44[2],stage1_43[17],stage1_42[23],stage1_41[23],stage1_40[38]}
   );
   gpc606_5 gpc388 (
      {stage0_40[64], stage0_40[65], stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69]},
      {stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17], stage0_42[18]},
      {stage1_44[3],stage1_43[18],stage1_42[24],stage1_41[24],stage1_40[39]}
   );
   gpc606_5 gpc389 (
      {stage0_40[70], stage0_40[71], stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75]},
      {stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23], stage0_42[24]},
      {stage1_44[4],stage1_43[19],stage1_42[25],stage1_41[25],stage1_40[40]}
   );
   gpc606_5 gpc390 (
      {stage0_40[76], stage0_40[77], stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81]},
      {stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29], stage0_42[30]},
      {stage1_44[5],stage1_43[20],stage1_42[26],stage1_41[26],stage1_40[41]}
   );
   gpc606_5 gpc391 (
      {stage0_40[82], stage0_40[83], stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87]},
      {stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35], stage0_42[36]},
      {stage1_44[6],stage1_43[21],stage1_42[27],stage1_41[27],stage1_40[42]}
   );
   gpc606_5 gpc392 (
      {stage0_40[88], stage0_40[89], stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93]},
      {stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41], stage0_42[42]},
      {stage1_44[7],stage1_43[22],stage1_42[28],stage1_41[28],stage1_40[43]}
   );
   gpc606_5 gpc393 (
      {stage0_40[94], stage0_40[95], stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99]},
      {stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47], stage0_42[48]},
      {stage1_44[8],stage1_43[23],stage1_42[29],stage1_41[29],stage1_40[44]}
   );
   gpc606_5 gpc394 (
      {stage0_40[100], stage0_40[101], stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105]},
      {stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53], stage0_42[54]},
      {stage1_44[9],stage1_43[24],stage1_42[30],stage1_41[30],stage1_40[45]}
   );
   gpc606_5 gpc395 (
      {stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111]},
      {stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59], stage0_42[60]},
      {stage1_44[10],stage1_43[25],stage1_42[31],stage1_41[31],stage1_40[46]}
   );
   gpc615_5 gpc396 (
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100]},
      {stage0_42[61]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[11],stage1_43[26],stage1_42[32],stage1_41[32]}
   );
   gpc615_5 gpc397 (
      {stage0_41[101], stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105]},
      {stage0_42[62]},
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage1_45[1],stage1_44[12],stage1_43[27],stage1_42[33],stage1_41[33]}
   );
   gpc615_5 gpc398 (
      {stage0_41[106], stage0_41[107], stage0_41[108], stage0_41[109], stage0_41[110]},
      {stage0_42[63]},
      {stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17], stage0_43[18]},
      {stage1_45[2],stage1_44[13],stage1_43[28],stage1_42[34],stage1_41[34]}
   );
   gpc615_5 gpc399 (
      {stage0_41[111], stage0_41[112], stage0_41[113], stage0_41[114], stage0_41[115]},
      {stage0_42[64]},
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23], stage0_43[24]},
      {stage1_45[3],stage1_44[14],stage1_43[29],stage1_42[35],stage1_41[35]}
   );
   gpc615_5 gpc400 (
      {stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119], stage0_41[120]},
      {stage0_42[65]},
      {stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29], stage0_43[30]},
      {stage1_45[4],stage1_44[15],stage1_43[30],stage1_42[36],stage1_41[36]}
   );
   gpc615_5 gpc401 (
      {stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_42[66]},
      {stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35], stage0_43[36]},
      {stage1_45[5],stage1_44[16],stage1_43[31],stage1_42[37],stage1_41[37]}
   );
   gpc615_5 gpc402 (
      {stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage0_43[37]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[6],stage1_44[17],stage1_43[32],stage1_42[38]}
   );
   gpc615_5 gpc403 (
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76]},
      {stage0_43[38]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[7],stage1_44[18],stage1_43[33],stage1_42[39]}
   );
   gpc615_5 gpc404 (
      {stage0_42[77], stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81]},
      {stage0_43[39]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[8],stage1_44[19],stage1_43[34],stage1_42[40]}
   );
   gpc615_5 gpc405 (
      {stage0_42[82], stage0_42[83], stage0_42[84], stage0_42[85], stage0_42[86]},
      {stage0_43[40]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[9],stage1_44[20],stage1_43[35],stage1_42[41]}
   );
   gpc615_5 gpc406 (
      {stage0_42[87], stage0_42[88], stage0_42[89], stage0_42[90], stage0_42[91]},
      {stage0_43[41]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[10],stage1_44[21],stage1_43[36],stage1_42[42]}
   );
   gpc615_5 gpc407 (
      {stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95], stage0_42[96]},
      {stage0_43[42]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[11],stage1_44[22],stage1_43[37],stage1_42[43]}
   );
   gpc615_5 gpc408 (
      {stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage0_43[43]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[12],stage1_44[23],stage1_43[38],stage1_42[44]}
   );
   gpc615_5 gpc409 (
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106]},
      {stage0_43[44]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[13],stage1_44[24],stage1_43[39],stage1_42[45]}
   );
   gpc615_5 gpc410 (
      {stage0_42[107], stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111]},
      {stage0_43[45]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[14],stage1_44[25],stage1_43[40],stage1_42[46]}
   );
   gpc615_5 gpc411 (
      {stage0_42[112], stage0_42[113], stage0_42[114], stage0_42[115], stage0_42[116]},
      {stage0_43[46]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[15],stage1_44[26],stage1_43[41],stage1_42[47]}
   );
   gpc615_5 gpc412 (
      {stage0_42[117], stage0_42[118], stage0_42[119], stage0_42[120], stage0_42[121]},
      {stage0_43[47]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[16],stage1_44[27],stage1_43[42],stage1_42[48]}
   );
   gpc615_5 gpc413 (
      {stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125], stage0_42[126]},
      {stage0_43[48]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[17],stage1_44[28],stage1_43[43],stage1_42[49]}
   );
   gpc615_5 gpc414 (
      {stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage0_44[72]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[12],stage1_45[18],stage1_44[29],stage1_43[44]}
   );
   gpc615_5 gpc415 (
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58]},
      {stage0_44[73]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[13],stage1_45[19],stage1_44[30],stage1_43[45]}
   );
   gpc615_5 gpc416 (
      {stage0_43[59], stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63]},
      {stage0_44[74]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[14],stage1_45[20],stage1_44[31],stage1_43[46]}
   );
   gpc615_5 gpc417 (
      {stage0_43[64], stage0_43[65], stage0_43[66], stage0_43[67], stage0_43[68]},
      {stage0_44[75]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[15],stage1_45[21],stage1_44[32],stage1_43[47]}
   );
   gpc615_5 gpc418 (
      {stage0_43[69], stage0_43[70], stage0_43[71], stage0_43[72], stage0_43[73]},
      {stage0_44[76]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[16],stage1_45[22],stage1_44[33],stage1_43[48]}
   );
   gpc615_5 gpc419 (
      {stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77], stage0_43[78]},
      {stage0_44[77]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[17],stage1_45[23],stage1_44[34],stage1_43[49]}
   );
   gpc615_5 gpc420 (
      {stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage0_44[78]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[18],stage1_45[24],stage1_44[35],stage1_43[50]}
   );
   gpc615_5 gpc421 (
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88]},
      {stage0_44[79]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[19],stage1_45[25],stage1_44[36],stage1_43[51]}
   );
   gpc615_5 gpc422 (
      {stage0_43[89], stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93]},
      {stage0_44[80]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[20],stage1_45[26],stage1_44[37],stage1_43[52]}
   );
   gpc615_5 gpc423 (
      {stage0_43[94], stage0_43[95], stage0_43[96], stage0_43[97], stage0_43[98]},
      {stage0_44[81]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[21],stage1_45[27],stage1_44[38],stage1_43[53]}
   );
   gpc615_5 gpc424 (
      {stage0_43[99], stage0_43[100], stage0_43[101], stage0_43[102], stage0_43[103]},
      {stage0_44[82]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[22],stage1_45[28],stage1_44[39],stage1_43[54]}
   );
   gpc606_5 gpc425 (
      {stage0_44[83], stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[11],stage1_46[23],stage1_45[29],stage1_44[40]}
   );
   gpc606_5 gpc426 (
      {stage0_44[89], stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[12],stage1_46[24],stage1_45[30],stage1_44[41]}
   );
   gpc606_5 gpc427 (
      {stage0_44[95], stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[13],stage1_46[25],stage1_45[31],stage1_44[42]}
   );
   gpc606_5 gpc428 (
      {stage0_44[101], stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[14],stage1_46[26],stage1_45[32],stage1_44[43]}
   );
   gpc606_5 gpc429 (
      {stage0_44[107], stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[15],stage1_46[27],stage1_45[33],stage1_44[44]}
   );
   gpc606_5 gpc430 (
      {stage0_44[113], stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[16],stage1_46[28],stage1_45[34],stage1_44[45]}
   );
   gpc606_5 gpc431 (
      {stage0_44[119], stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[17],stage1_46[29],stage1_45[35],stage1_44[46]}
   );
   gpc606_5 gpc432 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[7],stage1_47[18],stage1_46[30],stage1_45[36]}
   );
   gpc606_5 gpc433 (
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[8],stage1_47[19],stage1_46[31],stage1_45[37]}
   );
   gpc606_5 gpc434 (
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[9],stage1_47[20],stage1_46[32],stage1_45[38]}
   );
   gpc606_5 gpc435 (
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[10],stage1_47[21],stage1_46[33],stage1_45[39]}
   );
   gpc606_5 gpc436 (
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[11],stage1_47[22],stage1_46[34],stage1_45[40]}
   );
   gpc606_5 gpc437 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[12],stage1_47[23],stage1_46[35],stage1_45[41]}
   );
   gpc606_5 gpc438 (
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[13],stage1_47[24],stage1_46[36],stage1_45[42]}
   );
   gpc606_5 gpc439 (
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[14],stage1_47[25],stage1_46[37],stage1_45[43]}
   );
   gpc606_5 gpc440 (
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[8],stage1_48[15],stage1_47[26],stage1_46[38]}
   );
   gpc606_5 gpc441 (
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[9],stage1_48[16],stage1_47[27],stage1_46[39]}
   );
   gpc606_5 gpc442 (
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[10],stage1_48[17],stage1_47[28],stage1_46[40]}
   );
   gpc606_5 gpc443 (
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[11],stage1_48[18],stage1_47[29],stage1_46[41]}
   );
   gpc615_5 gpc444 (
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70]},
      {stage0_47[48]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[12],stage1_48[19],stage1_47[30],stage1_46[42]}
   );
   gpc615_5 gpc445 (
      {stage0_46[71], stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75]},
      {stage0_47[49]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[13],stage1_48[20],stage1_47[31],stage1_46[43]}
   );
   gpc615_5 gpc446 (
      {stage0_46[76], stage0_46[77], stage0_46[78], stage0_46[79], stage0_46[80]},
      {stage0_47[50]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[14],stage1_48[21],stage1_47[32],stage1_46[44]}
   );
   gpc615_5 gpc447 (
      {stage0_46[81], stage0_46[82], stage0_46[83], stage0_46[84], stage0_46[85]},
      {stage0_47[51]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[15],stage1_48[22],stage1_47[33],stage1_46[45]}
   );
   gpc1325_5 gpc448 (
      {stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89], stage0_46[90]},
      {stage0_47[52], stage0_47[53]},
      {stage0_48[48], stage0_48[49], stage0_48[50]},
      {stage0_49[0]},
      {stage1_50[8],stage1_49[16],stage1_48[23],stage1_47[34],stage1_46[46]}
   );
   gpc1325_5 gpc449 (
      {stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage0_47[54], stage0_47[55]},
      {stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage0_49[1]},
      {stage1_50[9],stage1_49[17],stage1_48[24],stage1_47[35],stage1_46[47]}
   );
   gpc2135_5 gpc450 (
      {stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59], stage0_47[60]},
      {stage0_48[54], stage0_48[55], stage0_48[56]},
      {stage0_49[2]},
      {stage0_50[0], stage0_50[1]},
      {stage1_51[0],stage1_50[10],stage1_49[18],stage1_48[25],stage1_47[36]}
   );
   gpc606_5 gpc451 (
      {stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65], stage0_47[66]},
      {stage0_49[3], stage0_49[4], stage0_49[5], stage0_49[6], stage0_49[7], stage0_49[8]},
      {stage1_51[1],stage1_50[11],stage1_49[19],stage1_48[26],stage1_47[37]}
   );
   gpc606_5 gpc452 (
      {stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71], stage0_47[72]},
      {stage0_49[9], stage0_49[10], stage0_49[11], stage0_49[12], stage0_49[13], stage0_49[14]},
      {stage1_51[2],stage1_50[12],stage1_49[20],stage1_48[27],stage1_47[38]}
   );
   gpc615_5 gpc453 (
      {stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage0_48[57]},
      {stage0_49[15], stage0_49[16], stage0_49[17], stage0_49[18], stage0_49[19], stage0_49[20]},
      {stage1_51[3],stage1_50[13],stage1_49[21],stage1_48[28],stage1_47[39]}
   );
   gpc615_5 gpc454 (
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82]},
      {stage0_48[58]},
      {stage0_49[21], stage0_49[22], stage0_49[23], stage0_49[24], stage0_49[25], stage0_49[26]},
      {stage1_51[4],stage1_50[14],stage1_49[22],stage1_48[29],stage1_47[40]}
   );
   gpc615_5 gpc455 (
      {stage0_47[83], stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87]},
      {stage0_48[59]},
      {stage0_49[27], stage0_49[28], stage0_49[29], stage0_49[30], stage0_49[31], stage0_49[32]},
      {stage1_51[5],stage1_50[15],stage1_49[23],stage1_48[30],stage1_47[41]}
   );
   gpc615_5 gpc456 (
      {stage0_47[88], stage0_47[89], stage0_47[90], stage0_47[91], stage0_47[92]},
      {stage0_48[60]},
      {stage0_49[33], stage0_49[34], stage0_49[35], stage0_49[36], stage0_49[37], stage0_49[38]},
      {stage1_51[6],stage1_50[16],stage1_49[24],stage1_48[31],stage1_47[42]}
   );
   gpc615_5 gpc457 (
      {stage0_47[93], stage0_47[94], stage0_47[95], stage0_47[96], stage0_47[97]},
      {stage0_48[61]},
      {stage0_49[39], stage0_49[40], stage0_49[41], stage0_49[42], stage0_49[43], stage0_49[44]},
      {stage1_51[7],stage1_50[17],stage1_49[25],stage1_48[32],stage1_47[43]}
   );
   gpc615_5 gpc458 (
      {stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101], stage0_47[102]},
      {stage0_48[62]},
      {stage0_49[45], stage0_49[46], stage0_49[47], stage0_49[48], stage0_49[49], stage0_49[50]},
      {stage1_51[8],stage1_50[18],stage1_49[26],stage1_48[33],stage1_47[44]}
   );
   gpc606_5 gpc459 (
      {stage0_48[63], stage0_48[64], stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68]},
      {stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5], stage0_50[6], stage0_50[7]},
      {stage1_52[0],stage1_51[9],stage1_50[19],stage1_49[27],stage1_48[34]}
   );
   gpc606_5 gpc460 (
      {stage0_48[69], stage0_48[70], stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74]},
      {stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11], stage0_50[12], stage0_50[13]},
      {stage1_52[1],stage1_51[10],stage1_50[20],stage1_49[28],stage1_48[35]}
   );
   gpc606_5 gpc461 (
      {stage0_48[75], stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80]},
      {stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17], stage0_50[18], stage0_50[19]},
      {stage1_52[2],stage1_51[11],stage1_50[21],stage1_49[29],stage1_48[36]}
   );
   gpc606_5 gpc462 (
      {stage0_48[81], stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85], stage0_48[86]},
      {stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23], stage0_50[24], stage0_50[25]},
      {stage1_52[3],stage1_51[12],stage1_50[22],stage1_49[30],stage1_48[37]}
   );
   gpc606_5 gpc463 (
      {stage0_48[87], stage0_48[88], stage0_48[89], stage0_48[90], stage0_48[91], stage0_48[92]},
      {stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29], stage0_50[30], stage0_50[31]},
      {stage1_52[4],stage1_51[13],stage1_50[23],stage1_49[31],stage1_48[38]}
   );
   gpc606_5 gpc464 (
      {stage0_48[93], stage0_48[94], stage0_48[95], stage0_48[96], stage0_48[97], stage0_48[98]},
      {stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35], stage0_50[36], stage0_50[37]},
      {stage1_52[5],stage1_51[14],stage1_50[24],stage1_49[32],stage1_48[39]}
   );
   gpc606_5 gpc465 (
      {stage0_48[99], stage0_48[100], stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104]},
      {stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41], stage0_50[42], stage0_50[43]},
      {stage1_52[6],stage1_51[15],stage1_50[25],stage1_49[33],stage1_48[40]}
   );
   gpc606_5 gpc466 (
      {stage0_48[105], stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110]},
      {stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47], stage0_50[48], stage0_50[49]},
      {stage1_52[7],stage1_51[16],stage1_50[26],stage1_49[34],stage1_48[41]}
   );
   gpc606_5 gpc467 (
      {stage0_48[111], stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116]},
      {stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53], stage0_50[54], stage0_50[55]},
      {stage1_52[8],stage1_51[17],stage1_50[27],stage1_49[35],stage1_48[42]}
   );
   gpc615_5 gpc468 (
      {stage0_48[117], stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121]},
      {stage0_49[51]},
      {stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59], stage0_50[60], stage0_50[61]},
      {stage1_52[9],stage1_51[18],stage1_50[28],stage1_49[36],stage1_48[43]}
   );
   gpc615_5 gpc469 (
      {stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125], stage0_48[126]},
      {stage0_49[52]},
      {stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65], stage0_50[66], stage0_50[67]},
      {stage1_52[10],stage1_51[19],stage1_50[29],stage1_49[37],stage1_48[44]}
   );
   gpc606_5 gpc470 (
      {stage0_49[53], stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[11],stage1_51[20],stage1_50[30],stage1_49[38]}
   );
   gpc606_5 gpc471 (
      {stage0_49[59], stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[12],stage1_51[21],stage1_50[31],stage1_49[39]}
   );
   gpc606_5 gpc472 (
      {stage0_49[65], stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[13],stage1_51[22],stage1_50[32],stage1_49[40]}
   );
   gpc606_5 gpc473 (
      {stage0_49[71], stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[14],stage1_51[23],stage1_50[33],stage1_49[41]}
   );
   gpc606_5 gpc474 (
      {stage0_49[77], stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[15],stage1_51[24],stage1_50[34],stage1_49[42]}
   );
   gpc606_5 gpc475 (
      {stage0_49[83], stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[16],stage1_51[25],stage1_50[35],stage1_49[43]}
   );
   gpc606_5 gpc476 (
      {stage0_49[89], stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[17],stage1_51[26],stage1_50[36],stage1_49[44]}
   );
   gpc606_5 gpc477 (
      {stage0_49[95], stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[18],stage1_51[27],stage1_50[37],stage1_49[45]}
   );
   gpc606_5 gpc478 (
      {stage0_49[101], stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[19],stage1_51[28],stage1_50[38],stage1_49[46]}
   );
   gpc606_5 gpc479 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[20],stage1_51[29],stage1_50[39],stage1_49[47]}
   );
   gpc606_5 gpc480 (
      {stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[21],stage1_51[30],stage1_50[40],stage1_49[48]}
   );
   gpc606_5 gpc481 (
      {stage0_49[119], stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[22],stage1_51[31],stage1_50[41],stage1_49[49]}
   );
   gpc623_5 gpc482 (
      {stage0_49[125], stage0_49[126], stage0_49[127]},
      {stage0_50[68], stage0_50[69]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[23],stage1_51[32],stage1_50[42],stage1_49[50]}
   );
   gpc606_5 gpc483 (
      {stage0_50[70], stage0_50[71], stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[13],stage1_52[24],stage1_51[33],stage1_50[43]}
   );
   gpc606_5 gpc484 (
      {stage0_50[76], stage0_50[77], stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[14],stage1_52[25],stage1_51[34],stage1_50[44]}
   );
   gpc606_5 gpc485 (
      {stage0_50[82], stage0_50[83], stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[15],stage1_52[26],stage1_51[35],stage1_50[45]}
   );
   gpc606_5 gpc486 (
      {stage0_50[88], stage0_50[89], stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[16],stage1_52[27],stage1_51[36],stage1_50[46]}
   );
   gpc606_5 gpc487 (
      {stage0_50[94], stage0_50[95], stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[17],stage1_52[28],stage1_51[37],stage1_50[47]}
   );
   gpc606_5 gpc488 (
      {stage0_50[100], stage0_50[101], stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[18],stage1_52[29],stage1_51[38],stage1_50[48]}
   );
   gpc606_5 gpc489 (
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[6],stage1_53[19],stage1_52[30],stage1_51[39]}
   );
   gpc606_5 gpc490 (
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[7],stage1_53[20],stage1_52[31],stage1_51[40]}
   );
   gpc606_5 gpc491 (
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[8],stage1_53[21],stage1_52[32],stage1_51[41]}
   );
   gpc606_5 gpc492 (
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[9],stage1_53[22],stage1_52[33],stage1_51[42]}
   );
   gpc606_5 gpc493 (
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[10],stage1_53[23],stage1_52[34],stage1_51[43]}
   );
   gpc606_5 gpc494 (
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[11],stage1_53[24],stage1_52[35],stage1_51[44]}
   );
   gpc606_5 gpc495 (
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[12],stage1_53[25],stage1_52[36],stage1_51[45]}
   );
   gpc606_5 gpc496 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[13],stage1_53[26],stage1_52[37],stage1_51[46]}
   );
   gpc606_5 gpc497 (
      {stage0_51[126], stage0_51[127], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[14],stage1_53[27],stage1_52[38],stage1_51[47]}
   );
   gpc606_5 gpc498 (
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[9],stage1_54[15],stage1_53[28],stage1_52[39]}
   );
   gpc606_5 gpc499 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[10],stage1_54[16],stage1_53[29],stage1_52[40]}
   );
   gpc606_5 gpc500 (
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[11],stage1_54[17],stage1_53[30],stage1_52[41]}
   );
   gpc606_5 gpc501 (
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[12],stage1_54[18],stage1_53[31],stage1_52[42]}
   );
   gpc606_5 gpc502 (
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[13],stage1_54[19],stage1_53[32],stage1_52[43]}
   );
   gpc606_5 gpc503 (
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[14],stage1_54[20],stage1_53[33],stage1_52[44]}
   );
   gpc606_5 gpc504 (
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[15],stage1_54[21],stage1_53[34],stage1_52[45]}
   );
   gpc606_5 gpc505 (
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[16],stage1_54[22],stage1_53[35],stage1_52[46]}
   );
   gpc606_5 gpc506 (
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[17],stage1_54[23],stage1_53[36],stage1_52[47]}
   );
   gpc606_5 gpc507 (
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[18],stage1_54[24],stage1_53[37],stage1_52[48]}
   );
   gpc606_5 gpc508 (
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[19],stage1_54[25],stage1_53[38],stage1_52[49]}
   );
   gpc606_5 gpc509 (
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[20],stage1_54[26],stage1_53[39],stage1_52[50]}
   );
   gpc606_5 gpc510 (
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[21],stage1_54[27],stage1_53[40],stage1_52[51]}
   );
   gpc606_5 gpc511 (
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[22],stage1_54[28],stage1_53[41],stage1_52[52]}
   );
   gpc1343_5 gpc512 (
      {stage0_53[54], stage0_53[55], stage0_53[56]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87]},
      {stage0_55[0], stage0_55[1], stage0_55[2]},
      {stage0_56[0]},
      {stage1_57[0],stage1_56[14],stage1_55[23],stage1_54[29],stage1_53[42]}
   );
   gpc606_5 gpc513 (
      {stage0_53[57], stage0_53[58], stage0_53[59], stage0_53[60], stage0_53[61], stage0_53[62]},
      {stage0_55[3], stage0_55[4], stage0_55[5], stage0_55[6], stage0_55[7], stage0_55[8]},
      {stage1_57[1],stage1_56[15],stage1_55[24],stage1_54[30],stage1_53[43]}
   );
   gpc606_5 gpc514 (
      {stage0_53[63], stage0_53[64], stage0_53[65], stage0_53[66], stage0_53[67], stage0_53[68]},
      {stage0_55[9], stage0_55[10], stage0_55[11], stage0_55[12], stage0_55[13], stage0_55[14]},
      {stage1_57[2],stage1_56[16],stage1_55[25],stage1_54[31],stage1_53[44]}
   );
   gpc606_5 gpc515 (
      {stage0_53[69], stage0_53[70], stage0_53[71], stage0_53[72], stage0_53[73], stage0_53[74]},
      {stage0_55[15], stage0_55[16], stage0_55[17], stage0_55[18], stage0_55[19], stage0_55[20]},
      {stage1_57[3],stage1_56[17],stage1_55[26],stage1_54[32],stage1_53[45]}
   );
   gpc606_5 gpc516 (
      {stage0_53[75], stage0_53[76], stage0_53[77], stage0_53[78], stage0_53[79], stage0_53[80]},
      {stage0_55[21], stage0_55[22], stage0_55[23], stage0_55[24], stage0_55[25], stage0_55[26]},
      {stage1_57[4],stage1_56[18],stage1_55[27],stage1_54[33],stage1_53[46]}
   );
   gpc606_5 gpc517 (
      {stage0_53[81], stage0_53[82], stage0_53[83], stage0_53[84], stage0_53[85], stage0_53[86]},
      {stage0_55[27], stage0_55[28], stage0_55[29], stage0_55[30], stage0_55[31], stage0_55[32]},
      {stage1_57[5],stage1_56[19],stage1_55[28],stage1_54[34],stage1_53[47]}
   );
   gpc606_5 gpc518 (
      {stage0_53[87], stage0_53[88], stage0_53[89], stage0_53[90], stage0_53[91], stage0_53[92]},
      {stage0_55[33], stage0_55[34], stage0_55[35], stage0_55[36], stage0_55[37], stage0_55[38]},
      {stage1_57[6],stage1_56[20],stage1_55[29],stage1_54[35],stage1_53[48]}
   );
   gpc606_5 gpc519 (
      {stage0_53[93], stage0_53[94], stage0_53[95], stage0_53[96], stage0_53[97], stage0_53[98]},
      {stage0_55[39], stage0_55[40], stage0_55[41], stage0_55[42], stage0_55[43], stage0_55[44]},
      {stage1_57[7],stage1_56[21],stage1_55[30],stage1_54[36],stage1_53[49]}
   );
   gpc606_5 gpc520 (
      {stage0_53[99], stage0_53[100], stage0_53[101], stage0_53[102], stage0_53[103], stage0_53[104]},
      {stage0_55[45], stage0_55[46], stage0_55[47], stage0_55[48], stage0_55[49], stage0_55[50]},
      {stage1_57[8],stage1_56[22],stage1_55[31],stage1_54[37],stage1_53[50]}
   );
   gpc615_5 gpc521 (
      {stage0_53[105], stage0_53[106], stage0_53[107], stage0_53[108], stage0_53[109]},
      {stage0_54[88]},
      {stage0_55[51], stage0_55[52], stage0_55[53], stage0_55[54], stage0_55[55], stage0_55[56]},
      {stage1_57[9],stage1_56[23],stage1_55[32],stage1_54[38],stage1_53[51]}
   );
   gpc615_5 gpc522 (
      {stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113], stage0_53[114]},
      {stage0_54[89]},
      {stage0_55[57], stage0_55[58], stage0_55[59], stage0_55[60], stage0_55[61], stage0_55[62]},
      {stage1_57[10],stage1_56[24],stage1_55[33],stage1_54[39],stage1_53[52]}
   );
   gpc615_5 gpc523 (
      {stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage0_54[90]},
      {stage0_55[63], stage0_55[64], stage0_55[65], stage0_55[66], stage0_55[67], stage0_55[68]},
      {stage1_57[11],stage1_56[25],stage1_55[34],stage1_54[40],stage1_53[53]}
   );
   gpc606_5 gpc524 (
      {stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95], stage0_54[96]},
      {stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6]},
      {stage1_58[0],stage1_57[12],stage1_56[26],stage1_55[35],stage1_54[41]}
   );
   gpc606_5 gpc525 (
      {stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101], stage0_54[102]},
      {stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12]},
      {stage1_58[1],stage1_57[13],stage1_56[27],stage1_55[36],stage1_54[42]}
   );
   gpc615_5 gpc526 (
      {stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage0_55[69]},
      {stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18]},
      {stage1_58[2],stage1_57[14],stage1_56[28],stage1_55[37],stage1_54[43]}
   );
   gpc615_5 gpc527 (
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112]},
      {stage0_55[70]},
      {stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24]},
      {stage1_58[3],stage1_57[15],stage1_56[29],stage1_55[38],stage1_54[44]}
   );
   gpc615_5 gpc528 (
      {stage0_54[113], stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117]},
      {stage0_55[71]},
      {stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30]},
      {stage1_58[4],stage1_57[16],stage1_56[30],stage1_55[39],stage1_54[45]}
   );
   gpc615_5 gpc529 (
      {stage0_54[118], stage0_54[119], stage0_54[120], stage0_54[121], stage0_54[122]},
      {stage0_55[72]},
      {stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36]},
      {stage1_58[5],stage1_57[17],stage1_56[31],stage1_55[40],stage1_54[46]}
   );
   gpc1163_5 gpc530 (
      {stage0_55[73], stage0_55[74], stage0_55[75]},
      {stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42]},
      {stage0_57[0]},
      {stage0_58[0]},
      {stage1_59[0],stage1_58[6],stage1_57[18],stage1_56[32],stage1_55[41]}
   );
   gpc1163_5 gpc531 (
      {stage0_55[76], stage0_55[77], stage0_55[78]},
      {stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48]},
      {stage0_57[1]},
      {stage0_58[1]},
      {stage1_59[1],stage1_58[7],stage1_57[19],stage1_56[33],stage1_55[42]}
   );
   gpc606_5 gpc532 (
      {stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83], stage0_55[84]},
      {stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6], stage0_57[7]},
      {stage1_59[2],stage1_58[8],stage1_57[20],stage1_56[34],stage1_55[43]}
   );
   gpc606_5 gpc533 (
      {stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89], stage0_55[90]},
      {stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11], stage0_57[12], stage0_57[13]},
      {stage1_59[3],stage1_58[9],stage1_57[21],stage1_56[35],stage1_55[44]}
   );
   gpc606_5 gpc534 (
      {stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95], stage0_55[96]},
      {stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17], stage0_57[18], stage0_57[19]},
      {stage1_59[4],stage1_58[10],stage1_57[22],stage1_56[36],stage1_55[45]}
   );
   gpc606_5 gpc535 (
      {stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101], stage0_55[102]},
      {stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23], stage0_57[24], stage0_57[25]},
      {stage1_59[5],stage1_58[11],stage1_57[23],stage1_56[37],stage1_55[46]}
   );
   gpc615_5 gpc536 (
      {stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage0_56[49]},
      {stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29], stage0_57[30], stage0_57[31]},
      {stage1_59[6],stage1_58[12],stage1_57[24],stage1_56[38],stage1_55[47]}
   );
   gpc606_5 gpc537 (
      {stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55]},
      {stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5], stage0_58[6], stage0_58[7]},
      {stage1_60[0],stage1_59[7],stage1_58[13],stage1_57[25],stage1_56[39]}
   );
   gpc606_5 gpc538 (
      {stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11], stage0_58[12], stage0_58[13]},
      {stage1_60[1],stage1_59[8],stage1_58[14],stage1_57[26],stage1_56[40]}
   );
   gpc606_5 gpc539 (
      {stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67]},
      {stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17], stage0_58[18], stage0_58[19]},
      {stage1_60[2],stage1_59[9],stage1_58[15],stage1_57[27],stage1_56[41]}
   );
   gpc606_5 gpc540 (
      {stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73]},
      {stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23], stage0_58[24], stage0_58[25]},
      {stage1_60[3],stage1_59[10],stage1_58[16],stage1_57[28],stage1_56[42]}
   );
   gpc606_5 gpc541 (
      {stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79]},
      {stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29], stage0_58[30], stage0_58[31]},
      {stage1_60[4],stage1_59[11],stage1_58[17],stage1_57[29],stage1_56[43]}
   );
   gpc606_5 gpc542 (
      {stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85]},
      {stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35], stage0_58[36], stage0_58[37]},
      {stage1_60[5],stage1_59[12],stage1_58[18],stage1_57[30],stage1_56[44]}
   );
   gpc606_5 gpc543 (
      {stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91]},
      {stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41], stage0_58[42], stage0_58[43]},
      {stage1_60[6],stage1_59[13],stage1_58[19],stage1_57[31],stage1_56[45]}
   );
   gpc606_5 gpc544 (
      {stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97]},
      {stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47], stage0_58[48], stage0_58[49]},
      {stage1_60[7],stage1_59[14],stage1_58[20],stage1_57[32],stage1_56[46]}
   );
   gpc606_5 gpc545 (
      {stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103]},
      {stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53], stage0_58[54], stage0_58[55]},
      {stage1_60[8],stage1_59[15],stage1_58[21],stage1_57[33],stage1_56[47]}
   );
   gpc606_5 gpc546 (
      {stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109]},
      {stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59], stage0_58[60], stage0_58[61]},
      {stage1_60[9],stage1_59[16],stage1_58[22],stage1_57[34],stage1_56[48]}
   );
   gpc606_5 gpc547 (
      {stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115]},
      {stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65], stage0_58[66], stage0_58[67]},
      {stage1_60[10],stage1_59[17],stage1_58[23],stage1_57[35],stage1_56[49]}
   );
   gpc606_5 gpc548 (
      {stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121]},
      {stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71], stage0_58[72], stage0_58[73]},
      {stage1_60[11],stage1_59[18],stage1_58[24],stage1_57[36],stage1_56[50]}
   );
   gpc606_5 gpc549 (
      {stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35], stage0_57[36], stage0_57[37]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[12],stage1_59[19],stage1_58[25],stage1_57[37]}
   );
   gpc606_5 gpc550 (
      {stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41], stage0_57[42], stage0_57[43]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[13],stage1_59[20],stage1_58[26],stage1_57[38]}
   );
   gpc606_5 gpc551 (
      {stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47], stage0_57[48], stage0_57[49]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[14],stage1_59[21],stage1_58[27],stage1_57[39]}
   );
   gpc606_5 gpc552 (
      {stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53], stage0_57[54], stage0_57[55]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[15],stage1_59[22],stage1_58[28],stage1_57[40]}
   );
   gpc606_5 gpc553 (
      {stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59], stage0_57[60], stage0_57[61]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[16],stage1_59[23],stage1_58[29],stage1_57[41]}
   );
   gpc606_5 gpc554 (
      {stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65], stage0_57[66], stage0_57[67]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[17],stage1_59[24],stage1_58[30],stage1_57[42]}
   );
   gpc606_5 gpc555 (
      {stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71], stage0_57[72], stage0_57[73]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[18],stage1_59[25],stage1_58[31],stage1_57[43]}
   );
   gpc606_5 gpc556 (
      {stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77], stage0_57[78], stage0_57[79]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[19],stage1_59[26],stage1_58[32],stage1_57[44]}
   );
   gpc606_5 gpc557 (
      {stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83], stage0_57[84], stage0_57[85]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[20],stage1_59[27],stage1_58[33],stage1_57[45]}
   );
   gpc606_5 gpc558 (
      {stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89], stage0_57[90], stage0_57[91]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[21],stage1_59[28],stage1_58[34],stage1_57[46]}
   );
   gpc606_5 gpc559 (
      {stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95], stage0_57[96], stage0_57[97]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[22],stage1_59[29],stage1_58[35],stage1_57[47]}
   );
   gpc606_5 gpc560 (
      {stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101], stage0_57[102], stage0_57[103]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[23],stage1_59[30],stage1_58[36],stage1_57[48]}
   );
   gpc606_5 gpc561 (
      {stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107], stage0_57[108], stage0_57[109]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[24],stage1_59[31],stage1_58[37],stage1_57[49]}
   );
   gpc606_5 gpc562 (
      {stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113], stage0_57[114], stage0_57[115]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[25],stage1_59[32],stage1_58[38],stage1_57[50]}
   );
   gpc606_5 gpc563 (
      {stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119], stage0_57[120], stage0_57[121]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[26],stage1_59[33],stage1_58[39],stage1_57[51]}
   );
   gpc615_5 gpc564 (
      {stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77], stage0_58[78]},
      {stage0_59[90]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[15],stage1_60[27],stage1_59[34],stage1_58[40]}
   );
   gpc615_5 gpc565 (
      {stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage0_59[91]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[16],stage1_60[28],stage1_59[35],stage1_58[41]}
   );
   gpc615_5 gpc566 (
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88]},
      {stage0_59[92]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[17],stage1_60[29],stage1_59[36],stage1_58[42]}
   );
   gpc615_5 gpc567 (
      {stage0_58[89], stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93]},
      {stage0_59[93]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[18],stage1_60[30],stage1_59[37],stage1_58[43]}
   );
   gpc615_5 gpc568 (
      {stage0_58[94], stage0_58[95], stage0_58[96], stage0_58[97], stage0_58[98]},
      {stage0_59[94]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[19],stage1_60[31],stage1_59[38],stage1_58[44]}
   );
   gpc615_5 gpc569 (
      {stage0_58[99], stage0_58[100], stage0_58[101], stage0_58[102], stage0_58[103]},
      {stage0_59[95]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[20],stage1_60[32],stage1_59[39],stage1_58[45]}
   );
   gpc615_5 gpc570 (
      {stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107], stage0_58[108]},
      {stage0_59[96]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[21],stage1_60[33],stage1_59[40],stage1_58[46]}
   );
   gpc615_5 gpc571 (
      {stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage0_59[97]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[22],stage1_60[34],stage1_59[41],stage1_58[47]}
   );
   gpc623_5 gpc572 (
      {stage0_58[114], stage0_58[115], stage0_58[116]},
      {stage0_59[98], stage0_59[99]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[23],stage1_60[35],stage1_59[42],stage1_58[48]}
   );
   gpc606_5 gpc573 (
      {stage0_59[100], stage0_59[101], stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[9],stage1_61[24],stage1_60[36],stage1_59[43]}
   );
   gpc606_5 gpc574 (
      {stage0_59[106], stage0_59[107], stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111]},
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage1_63[1],stage1_62[10],stage1_61[25],stage1_60[37],stage1_59[44]}
   );
   gpc606_5 gpc575 (
      {stage0_59[112], stage0_59[113], stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117]},
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage1_63[2],stage1_62[11],stage1_61[26],stage1_60[38],stage1_59[45]}
   );
   gpc606_5 gpc576 (
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[3],stage1_62[12],stage1_61[27],stage1_60[39]}
   );
   gpc606_5 gpc577 (
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[4],stage1_62[13],stage1_61[28],stage1_60[40]}
   );
   gpc606_5 gpc578 (
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[5],stage1_62[14],stage1_61[29],stage1_60[41]}
   );
   gpc606_5 gpc579 (
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[6],stage1_62[15],stage1_61[30],stage1_60[42]}
   );
   gpc606_5 gpc580 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[7],stage1_62[16],stage1_61[31],stage1_60[43]}
   );
   gpc606_5 gpc581 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[8],stage1_62[17],stage1_61[32],stage1_60[44]}
   );
   gpc606_5 gpc582 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[9],stage1_62[18],stage1_61[33],stage1_60[45]}
   );
   gpc606_5 gpc583 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[10],stage1_62[19],stage1_61[34],stage1_60[46]}
   );
   gpc606_5 gpc584 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[11],stage1_62[20],stage1_61[35],stage1_60[47]}
   );
   gpc606_5 gpc585 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[12],stage1_62[21],stage1_61[36],stage1_60[48]}
   );
   gpc606_5 gpc586 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[13],stage1_62[22],stage1_61[37],stage1_60[49]}
   );
   gpc606_5 gpc587 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[14],stage1_62[23],stage1_61[38],stage1_60[50]}
   );
   gpc606_5 gpc588 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[12],stage1_63[15],stage1_62[24],stage1_61[39]}
   );
   gpc606_5 gpc589 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[13],stage1_63[16],stage1_62[25],stage1_61[40]}
   );
   gpc606_5 gpc590 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[14],stage1_63[17],stage1_62[26],stage1_61[41]}
   );
   gpc606_5 gpc591 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[15],stage1_63[18],stage1_62[27],stage1_61[42]}
   );
   gpc606_5 gpc592 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[16],stage1_63[19],stage1_62[28],stage1_61[43]}
   );
   gpc606_5 gpc593 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[17],stage1_63[20],stage1_62[29],stage1_61[44]}
   );
   gpc606_5 gpc594 (
      {stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58], stage0_61[59]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[18],stage1_63[21],stage1_62[30],stage1_61[45]}
   );
   gpc606_5 gpc595 (
      {stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64], stage0_61[65]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[19],stage1_63[22],stage1_62[31],stage1_61[46]}
   );
   gpc606_5 gpc596 (
      {stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70], stage0_61[71]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[20],stage1_63[23],stage1_62[32],stage1_61[47]}
   );
   gpc606_5 gpc597 (
      {stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76], stage0_61[77]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[21],stage1_63[24],stage1_62[33],stage1_61[48]}
   );
   gpc606_5 gpc598 (
      {stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82], stage0_61[83]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[22],stage1_63[25],stage1_62[34],stage1_61[49]}
   );
   gpc606_5 gpc599 (
      {stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88], stage0_61[89]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[23],stage1_63[26],stage1_62[35],stage1_61[50]}
   );
   gpc606_5 gpc600 (
      {stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94], stage0_61[95]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[24],stage1_63[27],stage1_62[36],stage1_61[51]}
   );
   gpc606_5 gpc601 (
      {stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100], stage0_61[101]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[25],stage1_63[28],stage1_62[37],stage1_61[52]}
   );
   gpc606_5 gpc602 (
      {stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106], stage0_61[107]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[26],stage1_63[29],stage1_62[38],stage1_61[53]}
   );
   gpc606_5 gpc603 (
      {stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112], stage0_61[113]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[27],stage1_63[30],stage1_62[39],stage1_61[54]}
   );
   gpc606_5 gpc604 (
      {stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118], stage0_61[119]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[28],stage1_63[31],stage1_62[40],stage1_61[55]}
   );
   gpc606_5 gpc605 (
      {stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124], stage0_61[125]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[29],stage1_63[32],stage1_62[41],stage1_61[56]}
   );
   gpc1_1 gpc606 (
      {stage0_2[121]},
      {stage1_2[40]}
   );
   gpc1_1 gpc607 (
      {stage0_2[122]},
      {stage1_2[41]}
   );
   gpc1_1 gpc608 (
      {stage0_2[123]},
      {stage1_2[42]}
   );
   gpc1_1 gpc609 (
      {stage0_2[124]},
      {stage1_2[43]}
   );
   gpc1_1 gpc610 (
      {stage0_2[125]},
      {stage1_2[44]}
   );
   gpc1_1 gpc611 (
      {stage0_2[126]},
      {stage1_2[45]}
   );
   gpc1_1 gpc612 (
      {stage0_2[127]},
      {stage1_2[46]}
   );
   gpc1_1 gpc613 (
      {stage0_3[117]},
      {stage1_3[56]}
   );
   gpc1_1 gpc614 (
      {stage0_3[118]},
      {stage1_3[57]}
   );
   gpc1_1 gpc615 (
      {stage0_3[119]},
      {stage1_3[58]}
   );
   gpc1_1 gpc616 (
      {stage0_3[120]},
      {stage1_3[59]}
   );
   gpc1_1 gpc617 (
      {stage0_3[121]},
      {stage1_3[60]}
   );
   gpc1_1 gpc618 (
      {stage0_3[122]},
      {stage1_3[61]}
   );
   gpc1_1 gpc619 (
      {stage0_3[123]},
      {stage1_3[62]}
   );
   gpc1_1 gpc620 (
      {stage0_3[124]},
      {stage1_3[63]}
   );
   gpc1_1 gpc621 (
      {stage0_3[125]},
      {stage1_3[64]}
   );
   gpc1_1 gpc622 (
      {stage0_3[126]},
      {stage1_3[65]}
   );
   gpc1_1 gpc623 (
      {stage0_3[127]},
      {stage1_3[66]}
   );
   gpc1_1 gpc624 (
      {stage0_5[118]},
      {stage1_5[42]}
   );
   gpc1_1 gpc625 (
      {stage0_5[119]},
      {stage1_5[43]}
   );
   gpc1_1 gpc626 (
      {stage0_5[120]},
      {stage1_5[44]}
   );
   gpc1_1 gpc627 (
      {stage0_5[121]},
      {stage1_5[45]}
   );
   gpc1_1 gpc628 (
      {stage0_5[122]},
      {stage1_5[46]}
   );
   gpc1_1 gpc629 (
      {stage0_5[123]},
      {stage1_5[47]}
   );
   gpc1_1 gpc630 (
      {stage0_5[124]},
      {stage1_5[48]}
   );
   gpc1_1 gpc631 (
      {stage0_5[125]},
      {stage1_5[49]}
   );
   gpc1_1 gpc632 (
      {stage0_5[126]},
      {stage1_5[50]}
   );
   gpc1_1 gpc633 (
      {stage0_5[127]},
      {stage1_5[51]}
   );
   gpc1_1 gpc634 (
      {stage0_6[79]},
      {stage1_6[40]}
   );
   gpc1_1 gpc635 (
      {stage0_6[80]},
      {stage1_6[41]}
   );
   gpc1_1 gpc636 (
      {stage0_6[81]},
      {stage1_6[42]}
   );
   gpc1_1 gpc637 (
      {stage0_6[82]},
      {stage1_6[43]}
   );
   gpc1_1 gpc638 (
      {stage0_6[83]},
      {stage1_6[44]}
   );
   gpc1_1 gpc639 (
      {stage0_6[84]},
      {stage1_6[45]}
   );
   gpc1_1 gpc640 (
      {stage0_6[85]},
      {stage1_6[46]}
   );
   gpc1_1 gpc641 (
      {stage0_6[86]},
      {stage1_6[47]}
   );
   gpc1_1 gpc642 (
      {stage0_6[87]},
      {stage1_6[48]}
   );
   gpc1_1 gpc643 (
      {stage0_6[88]},
      {stage1_6[49]}
   );
   gpc1_1 gpc644 (
      {stage0_6[89]},
      {stage1_6[50]}
   );
   gpc1_1 gpc645 (
      {stage0_6[90]},
      {stage1_6[51]}
   );
   gpc1_1 gpc646 (
      {stage0_6[91]},
      {stage1_6[52]}
   );
   gpc1_1 gpc647 (
      {stage0_6[92]},
      {stage1_6[53]}
   );
   gpc1_1 gpc648 (
      {stage0_6[93]},
      {stage1_6[54]}
   );
   gpc1_1 gpc649 (
      {stage0_6[94]},
      {stage1_6[55]}
   );
   gpc1_1 gpc650 (
      {stage0_6[95]},
      {stage1_6[56]}
   );
   gpc1_1 gpc651 (
      {stage0_6[96]},
      {stage1_6[57]}
   );
   gpc1_1 gpc652 (
      {stage0_6[97]},
      {stage1_6[58]}
   );
   gpc1_1 gpc653 (
      {stage0_6[98]},
      {stage1_6[59]}
   );
   gpc1_1 gpc654 (
      {stage0_6[99]},
      {stage1_6[60]}
   );
   gpc1_1 gpc655 (
      {stage0_6[100]},
      {stage1_6[61]}
   );
   gpc1_1 gpc656 (
      {stage0_6[101]},
      {stage1_6[62]}
   );
   gpc1_1 gpc657 (
      {stage0_6[102]},
      {stage1_6[63]}
   );
   gpc1_1 gpc658 (
      {stage0_6[103]},
      {stage1_6[64]}
   );
   gpc1_1 gpc659 (
      {stage0_6[104]},
      {stage1_6[65]}
   );
   gpc1_1 gpc660 (
      {stage0_6[105]},
      {stage1_6[66]}
   );
   gpc1_1 gpc661 (
      {stage0_6[106]},
      {stage1_6[67]}
   );
   gpc1_1 gpc662 (
      {stage0_6[107]},
      {stage1_6[68]}
   );
   gpc1_1 gpc663 (
      {stage0_6[108]},
      {stage1_6[69]}
   );
   gpc1_1 gpc664 (
      {stage0_6[109]},
      {stage1_6[70]}
   );
   gpc1_1 gpc665 (
      {stage0_6[110]},
      {stage1_6[71]}
   );
   gpc1_1 gpc666 (
      {stage0_6[111]},
      {stage1_6[72]}
   );
   gpc1_1 gpc667 (
      {stage0_6[112]},
      {stage1_6[73]}
   );
   gpc1_1 gpc668 (
      {stage0_6[113]},
      {stage1_6[74]}
   );
   gpc1_1 gpc669 (
      {stage0_6[114]},
      {stage1_6[75]}
   );
   gpc1_1 gpc670 (
      {stage0_6[115]},
      {stage1_6[76]}
   );
   gpc1_1 gpc671 (
      {stage0_6[116]},
      {stage1_6[77]}
   );
   gpc1_1 gpc672 (
      {stage0_6[117]},
      {stage1_6[78]}
   );
   gpc1_1 gpc673 (
      {stage0_6[118]},
      {stage1_6[79]}
   );
   gpc1_1 gpc674 (
      {stage0_6[119]},
      {stage1_6[80]}
   );
   gpc1_1 gpc675 (
      {stage0_6[120]},
      {stage1_6[81]}
   );
   gpc1_1 gpc676 (
      {stage0_6[121]},
      {stage1_6[82]}
   );
   gpc1_1 gpc677 (
      {stage0_6[122]},
      {stage1_6[83]}
   );
   gpc1_1 gpc678 (
      {stage0_6[123]},
      {stage1_6[84]}
   );
   gpc1_1 gpc679 (
      {stage0_6[124]},
      {stage1_6[85]}
   );
   gpc1_1 gpc680 (
      {stage0_6[125]},
      {stage1_6[86]}
   );
   gpc1_1 gpc681 (
      {stage0_6[126]},
      {stage1_6[87]}
   );
   gpc1_1 gpc682 (
      {stage0_6[127]},
      {stage1_6[88]}
   );
   gpc1_1 gpc683 (
      {stage0_7[103]},
      {stage1_7[46]}
   );
   gpc1_1 gpc684 (
      {stage0_7[104]},
      {stage1_7[47]}
   );
   gpc1_1 gpc685 (
      {stage0_7[105]},
      {stage1_7[48]}
   );
   gpc1_1 gpc686 (
      {stage0_7[106]},
      {stage1_7[49]}
   );
   gpc1_1 gpc687 (
      {stage0_7[107]},
      {stage1_7[50]}
   );
   gpc1_1 gpc688 (
      {stage0_7[108]},
      {stage1_7[51]}
   );
   gpc1_1 gpc689 (
      {stage0_7[109]},
      {stage1_7[52]}
   );
   gpc1_1 gpc690 (
      {stage0_7[110]},
      {stage1_7[53]}
   );
   gpc1_1 gpc691 (
      {stage0_7[111]},
      {stage1_7[54]}
   );
   gpc1_1 gpc692 (
      {stage0_7[112]},
      {stage1_7[55]}
   );
   gpc1_1 gpc693 (
      {stage0_7[113]},
      {stage1_7[56]}
   );
   gpc1_1 gpc694 (
      {stage0_7[114]},
      {stage1_7[57]}
   );
   gpc1_1 gpc695 (
      {stage0_7[115]},
      {stage1_7[58]}
   );
   gpc1_1 gpc696 (
      {stage0_7[116]},
      {stage1_7[59]}
   );
   gpc1_1 gpc697 (
      {stage0_7[117]},
      {stage1_7[60]}
   );
   gpc1_1 gpc698 (
      {stage0_7[118]},
      {stage1_7[61]}
   );
   gpc1_1 gpc699 (
      {stage0_7[119]},
      {stage1_7[62]}
   );
   gpc1_1 gpc700 (
      {stage0_7[120]},
      {stage1_7[63]}
   );
   gpc1_1 gpc701 (
      {stage0_7[121]},
      {stage1_7[64]}
   );
   gpc1_1 gpc702 (
      {stage0_7[122]},
      {stage1_7[65]}
   );
   gpc1_1 gpc703 (
      {stage0_7[123]},
      {stage1_7[66]}
   );
   gpc1_1 gpc704 (
      {stage0_7[124]},
      {stage1_7[67]}
   );
   gpc1_1 gpc705 (
      {stage0_7[125]},
      {stage1_7[68]}
   );
   gpc1_1 gpc706 (
      {stage0_7[126]},
      {stage1_7[69]}
   );
   gpc1_1 gpc707 (
      {stage0_7[127]},
      {stage1_7[70]}
   );
   gpc1_1 gpc708 (
      {stage0_8[109]},
      {stage1_8[47]}
   );
   gpc1_1 gpc709 (
      {stage0_8[110]},
      {stage1_8[48]}
   );
   gpc1_1 gpc710 (
      {stage0_8[111]},
      {stage1_8[49]}
   );
   gpc1_1 gpc711 (
      {stage0_8[112]},
      {stage1_8[50]}
   );
   gpc1_1 gpc712 (
      {stage0_8[113]},
      {stage1_8[51]}
   );
   gpc1_1 gpc713 (
      {stage0_8[114]},
      {stage1_8[52]}
   );
   gpc1_1 gpc714 (
      {stage0_8[115]},
      {stage1_8[53]}
   );
   gpc1_1 gpc715 (
      {stage0_8[116]},
      {stage1_8[54]}
   );
   gpc1_1 gpc716 (
      {stage0_8[117]},
      {stage1_8[55]}
   );
   gpc1_1 gpc717 (
      {stage0_8[118]},
      {stage1_8[56]}
   );
   gpc1_1 gpc718 (
      {stage0_8[119]},
      {stage1_8[57]}
   );
   gpc1_1 gpc719 (
      {stage0_8[120]},
      {stage1_8[58]}
   );
   gpc1_1 gpc720 (
      {stage0_8[121]},
      {stage1_8[59]}
   );
   gpc1_1 gpc721 (
      {stage0_8[122]},
      {stage1_8[60]}
   );
   gpc1_1 gpc722 (
      {stage0_8[123]},
      {stage1_8[61]}
   );
   gpc1_1 gpc723 (
      {stage0_8[124]},
      {stage1_8[62]}
   );
   gpc1_1 gpc724 (
      {stage0_8[125]},
      {stage1_8[63]}
   );
   gpc1_1 gpc725 (
      {stage0_8[126]},
      {stage1_8[64]}
   );
   gpc1_1 gpc726 (
      {stage0_8[127]},
      {stage1_8[65]}
   );
   gpc1_1 gpc727 (
      {stage0_9[108]},
      {stage1_9[41]}
   );
   gpc1_1 gpc728 (
      {stage0_9[109]},
      {stage1_9[42]}
   );
   gpc1_1 gpc729 (
      {stage0_9[110]},
      {stage1_9[43]}
   );
   gpc1_1 gpc730 (
      {stage0_9[111]},
      {stage1_9[44]}
   );
   gpc1_1 gpc731 (
      {stage0_9[112]},
      {stage1_9[45]}
   );
   gpc1_1 gpc732 (
      {stage0_9[113]},
      {stage1_9[46]}
   );
   gpc1_1 gpc733 (
      {stage0_9[114]},
      {stage1_9[47]}
   );
   gpc1_1 gpc734 (
      {stage0_9[115]},
      {stage1_9[48]}
   );
   gpc1_1 gpc735 (
      {stage0_9[116]},
      {stage1_9[49]}
   );
   gpc1_1 gpc736 (
      {stage0_9[117]},
      {stage1_9[50]}
   );
   gpc1_1 gpc737 (
      {stage0_9[118]},
      {stage1_9[51]}
   );
   gpc1_1 gpc738 (
      {stage0_9[119]},
      {stage1_9[52]}
   );
   gpc1_1 gpc739 (
      {stage0_9[120]},
      {stage1_9[53]}
   );
   gpc1_1 gpc740 (
      {stage0_9[121]},
      {stage1_9[54]}
   );
   gpc1_1 gpc741 (
      {stage0_9[122]},
      {stage1_9[55]}
   );
   gpc1_1 gpc742 (
      {stage0_9[123]},
      {stage1_9[56]}
   );
   gpc1_1 gpc743 (
      {stage0_9[124]},
      {stage1_9[57]}
   );
   gpc1_1 gpc744 (
      {stage0_9[125]},
      {stage1_9[58]}
   );
   gpc1_1 gpc745 (
      {stage0_9[126]},
      {stage1_9[59]}
   );
   gpc1_1 gpc746 (
      {stage0_9[127]},
      {stage1_9[60]}
   );
   gpc1_1 gpc747 (
      {stage0_11[118]},
      {stage1_11[54]}
   );
   gpc1_1 gpc748 (
      {stage0_11[119]},
      {stage1_11[55]}
   );
   gpc1_1 gpc749 (
      {stage0_11[120]},
      {stage1_11[56]}
   );
   gpc1_1 gpc750 (
      {stage0_11[121]},
      {stage1_11[57]}
   );
   gpc1_1 gpc751 (
      {stage0_11[122]},
      {stage1_11[58]}
   );
   gpc1_1 gpc752 (
      {stage0_11[123]},
      {stage1_11[59]}
   );
   gpc1_1 gpc753 (
      {stage0_11[124]},
      {stage1_11[60]}
   );
   gpc1_1 gpc754 (
      {stage0_11[125]},
      {stage1_11[61]}
   );
   gpc1_1 gpc755 (
      {stage0_11[126]},
      {stage1_11[62]}
   );
   gpc1_1 gpc756 (
      {stage0_11[127]},
      {stage1_11[63]}
   );
   gpc1_1 gpc757 (
      {stage0_13[124]},
      {stage1_13[50]}
   );
   gpc1_1 gpc758 (
      {stage0_13[125]},
      {stage1_13[51]}
   );
   gpc1_1 gpc759 (
      {stage0_13[126]},
      {stage1_13[52]}
   );
   gpc1_1 gpc760 (
      {stage0_13[127]},
      {stage1_13[53]}
   );
   gpc1_1 gpc761 (
      {stage0_14[109]},
      {stage1_14[47]}
   );
   gpc1_1 gpc762 (
      {stage0_14[110]},
      {stage1_14[48]}
   );
   gpc1_1 gpc763 (
      {stage0_14[111]},
      {stage1_14[49]}
   );
   gpc1_1 gpc764 (
      {stage0_14[112]},
      {stage1_14[50]}
   );
   gpc1_1 gpc765 (
      {stage0_14[113]},
      {stage1_14[51]}
   );
   gpc1_1 gpc766 (
      {stage0_14[114]},
      {stage1_14[52]}
   );
   gpc1_1 gpc767 (
      {stage0_14[115]},
      {stage1_14[53]}
   );
   gpc1_1 gpc768 (
      {stage0_14[116]},
      {stage1_14[54]}
   );
   gpc1_1 gpc769 (
      {stage0_14[117]},
      {stage1_14[55]}
   );
   gpc1_1 gpc770 (
      {stage0_14[118]},
      {stage1_14[56]}
   );
   gpc1_1 gpc771 (
      {stage0_14[119]},
      {stage1_14[57]}
   );
   gpc1_1 gpc772 (
      {stage0_14[120]},
      {stage1_14[58]}
   );
   gpc1_1 gpc773 (
      {stage0_14[121]},
      {stage1_14[59]}
   );
   gpc1_1 gpc774 (
      {stage0_14[122]},
      {stage1_14[60]}
   );
   gpc1_1 gpc775 (
      {stage0_14[123]},
      {stage1_14[61]}
   );
   gpc1_1 gpc776 (
      {stage0_14[124]},
      {stage1_14[62]}
   );
   gpc1_1 gpc777 (
      {stage0_14[125]},
      {stage1_14[63]}
   );
   gpc1_1 gpc778 (
      {stage0_14[126]},
      {stage1_14[64]}
   );
   gpc1_1 gpc779 (
      {stage0_14[127]},
      {stage1_14[65]}
   );
   gpc1_1 gpc780 (
      {stage0_15[106]},
      {stage1_15[46]}
   );
   gpc1_1 gpc781 (
      {stage0_15[107]},
      {stage1_15[47]}
   );
   gpc1_1 gpc782 (
      {stage0_15[108]},
      {stage1_15[48]}
   );
   gpc1_1 gpc783 (
      {stage0_15[109]},
      {stage1_15[49]}
   );
   gpc1_1 gpc784 (
      {stage0_15[110]},
      {stage1_15[50]}
   );
   gpc1_1 gpc785 (
      {stage0_15[111]},
      {stage1_15[51]}
   );
   gpc1_1 gpc786 (
      {stage0_15[112]},
      {stage1_15[52]}
   );
   gpc1_1 gpc787 (
      {stage0_15[113]},
      {stage1_15[53]}
   );
   gpc1_1 gpc788 (
      {stage0_15[114]},
      {stage1_15[54]}
   );
   gpc1_1 gpc789 (
      {stage0_15[115]},
      {stage1_15[55]}
   );
   gpc1_1 gpc790 (
      {stage0_15[116]},
      {stage1_15[56]}
   );
   gpc1_1 gpc791 (
      {stage0_15[117]},
      {stage1_15[57]}
   );
   gpc1_1 gpc792 (
      {stage0_15[118]},
      {stage1_15[58]}
   );
   gpc1_1 gpc793 (
      {stage0_15[119]},
      {stage1_15[59]}
   );
   gpc1_1 gpc794 (
      {stage0_15[120]},
      {stage1_15[60]}
   );
   gpc1_1 gpc795 (
      {stage0_15[121]},
      {stage1_15[61]}
   );
   gpc1_1 gpc796 (
      {stage0_15[122]},
      {stage1_15[62]}
   );
   gpc1_1 gpc797 (
      {stage0_15[123]},
      {stage1_15[63]}
   );
   gpc1_1 gpc798 (
      {stage0_15[124]},
      {stage1_15[64]}
   );
   gpc1_1 gpc799 (
      {stage0_15[125]},
      {stage1_15[65]}
   );
   gpc1_1 gpc800 (
      {stage0_15[126]},
      {stage1_15[66]}
   );
   gpc1_1 gpc801 (
      {stage0_15[127]},
      {stage1_15[67]}
   );
   gpc1_1 gpc802 (
      {stage0_16[85]},
      {stage1_16[46]}
   );
   gpc1_1 gpc803 (
      {stage0_16[86]},
      {stage1_16[47]}
   );
   gpc1_1 gpc804 (
      {stage0_16[87]},
      {stage1_16[48]}
   );
   gpc1_1 gpc805 (
      {stage0_16[88]},
      {stage1_16[49]}
   );
   gpc1_1 gpc806 (
      {stage0_16[89]},
      {stage1_16[50]}
   );
   gpc1_1 gpc807 (
      {stage0_16[90]},
      {stage1_16[51]}
   );
   gpc1_1 gpc808 (
      {stage0_16[91]},
      {stage1_16[52]}
   );
   gpc1_1 gpc809 (
      {stage0_16[92]},
      {stage1_16[53]}
   );
   gpc1_1 gpc810 (
      {stage0_16[93]},
      {stage1_16[54]}
   );
   gpc1_1 gpc811 (
      {stage0_16[94]},
      {stage1_16[55]}
   );
   gpc1_1 gpc812 (
      {stage0_16[95]},
      {stage1_16[56]}
   );
   gpc1_1 gpc813 (
      {stage0_16[96]},
      {stage1_16[57]}
   );
   gpc1_1 gpc814 (
      {stage0_16[97]},
      {stage1_16[58]}
   );
   gpc1_1 gpc815 (
      {stage0_16[98]},
      {stage1_16[59]}
   );
   gpc1_1 gpc816 (
      {stage0_16[99]},
      {stage1_16[60]}
   );
   gpc1_1 gpc817 (
      {stage0_16[100]},
      {stage1_16[61]}
   );
   gpc1_1 gpc818 (
      {stage0_16[101]},
      {stage1_16[62]}
   );
   gpc1_1 gpc819 (
      {stage0_16[102]},
      {stage1_16[63]}
   );
   gpc1_1 gpc820 (
      {stage0_16[103]},
      {stage1_16[64]}
   );
   gpc1_1 gpc821 (
      {stage0_16[104]},
      {stage1_16[65]}
   );
   gpc1_1 gpc822 (
      {stage0_16[105]},
      {stage1_16[66]}
   );
   gpc1_1 gpc823 (
      {stage0_16[106]},
      {stage1_16[67]}
   );
   gpc1_1 gpc824 (
      {stage0_16[107]},
      {stage1_16[68]}
   );
   gpc1_1 gpc825 (
      {stage0_16[108]},
      {stage1_16[69]}
   );
   gpc1_1 gpc826 (
      {stage0_16[109]},
      {stage1_16[70]}
   );
   gpc1_1 gpc827 (
      {stage0_16[110]},
      {stage1_16[71]}
   );
   gpc1_1 gpc828 (
      {stage0_16[111]},
      {stage1_16[72]}
   );
   gpc1_1 gpc829 (
      {stage0_16[112]},
      {stage1_16[73]}
   );
   gpc1_1 gpc830 (
      {stage0_16[113]},
      {stage1_16[74]}
   );
   gpc1_1 gpc831 (
      {stage0_16[114]},
      {stage1_16[75]}
   );
   gpc1_1 gpc832 (
      {stage0_16[115]},
      {stage1_16[76]}
   );
   gpc1_1 gpc833 (
      {stage0_16[116]},
      {stage1_16[77]}
   );
   gpc1_1 gpc834 (
      {stage0_16[117]},
      {stage1_16[78]}
   );
   gpc1_1 gpc835 (
      {stage0_16[118]},
      {stage1_16[79]}
   );
   gpc1_1 gpc836 (
      {stage0_16[119]},
      {stage1_16[80]}
   );
   gpc1_1 gpc837 (
      {stage0_16[120]},
      {stage1_16[81]}
   );
   gpc1_1 gpc838 (
      {stage0_16[121]},
      {stage1_16[82]}
   );
   gpc1_1 gpc839 (
      {stage0_16[122]},
      {stage1_16[83]}
   );
   gpc1_1 gpc840 (
      {stage0_16[123]},
      {stage1_16[84]}
   );
   gpc1_1 gpc841 (
      {stage0_16[124]},
      {stage1_16[85]}
   );
   gpc1_1 gpc842 (
      {stage0_16[125]},
      {stage1_16[86]}
   );
   gpc1_1 gpc843 (
      {stage0_16[126]},
      {stage1_16[87]}
   );
   gpc1_1 gpc844 (
      {stage0_16[127]},
      {stage1_16[88]}
   );
   gpc1_1 gpc845 (
      {stage0_17[103]},
      {stage1_17[42]}
   );
   gpc1_1 gpc846 (
      {stage0_17[104]},
      {stage1_17[43]}
   );
   gpc1_1 gpc847 (
      {stage0_17[105]},
      {stage1_17[44]}
   );
   gpc1_1 gpc848 (
      {stage0_17[106]},
      {stage1_17[45]}
   );
   gpc1_1 gpc849 (
      {stage0_17[107]},
      {stage1_17[46]}
   );
   gpc1_1 gpc850 (
      {stage0_17[108]},
      {stage1_17[47]}
   );
   gpc1_1 gpc851 (
      {stage0_17[109]},
      {stage1_17[48]}
   );
   gpc1_1 gpc852 (
      {stage0_17[110]},
      {stage1_17[49]}
   );
   gpc1_1 gpc853 (
      {stage0_17[111]},
      {stage1_17[50]}
   );
   gpc1_1 gpc854 (
      {stage0_17[112]},
      {stage1_17[51]}
   );
   gpc1_1 gpc855 (
      {stage0_17[113]},
      {stage1_17[52]}
   );
   gpc1_1 gpc856 (
      {stage0_17[114]},
      {stage1_17[53]}
   );
   gpc1_1 gpc857 (
      {stage0_17[115]},
      {stage1_17[54]}
   );
   gpc1_1 gpc858 (
      {stage0_17[116]},
      {stage1_17[55]}
   );
   gpc1_1 gpc859 (
      {stage0_17[117]},
      {stage1_17[56]}
   );
   gpc1_1 gpc860 (
      {stage0_17[118]},
      {stage1_17[57]}
   );
   gpc1_1 gpc861 (
      {stage0_17[119]},
      {stage1_17[58]}
   );
   gpc1_1 gpc862 (
      {stage0_17[120]},
      {stage1_17[59]}
   );
   gpc1_1 gpc863 (
      {stage0_17[121]},
      {stage1_17[60]}
   );
   gpc1_1 gpc864 (
      {stage0_17[122]},
      {stage1_17[61]}
   );
   gpc1_1 gpc865 (
      {stage0_17[123]},
      {stage1_17[62]}
   );
   gpc1_1 gpc866 (
      {stage0_17[124]},
      {stage1_17[63]}
   );
   gpc1_1 gpc867 (
      {stage0_17[125]},
      {stage1_17[64]}
   );
   gpc1_1 gpc868 (
      {stage0_17[126]},
      {stage1_17[65]}
   );
   gpc1_1 gpc869 (
      {stage0_17[127]},
      {stage1_17[66]}
   );
   gpc1_1 gpc870 (
      {stage0_19[123]},
      {stage1_19[50]}
   );
   gpc1_1 gpc871 (
      {stage0_19[124]},
      {stage1_19[51]}
   );
   gpc1_1 gpc872 (
      {stage0_19[125]},
      {stage1_19[52]}
   );
   gpc1_1 gpc873 (
      {stage0_19[126]},
      {stage1_19[53]}
   );
   gpc1_1 gpc874 (
      {stage0_19[127]},
      {stage1_19[54]}
   );
   gpc1_1 gpc875 (
      {stage0_20[104]},
      {stage1_20[48]}
   );
   gpc1_1 gpc876 (
      {stage0_20[105]},
      {stage1_20[49]}
   );
   gpc1_1 gpc877 (
      {stage0_20[106]},
      {stage1_20[50]}
   );
   gpc1_1 gpc878 (
      {stage0_20[107]},
      {stage1_20[51]}
   );
   gpc1_1 gpc879 (
      {stage0_20[108]},
      {stage1_20[52]}
   );
   gpc1_1 gpc880 (
      {stage0_20[109]},
      {stage1_20[53]}
   );
   gpc1_1 gpc881 (
      {stage0_20[110]},
      {stage1_20[54]}
   );
   gpc1_1 gpc882 (
      {stage0_20[111]},
      {stage1_20[55]}
   );
   gpc1_1 gpc883 (
      {stage0_20[112]},
      {stage1_20[56]}
   );
   gpc1_1 gpc884 (
      {stage0_20[113]},
      {stage1_20[57]}
   );
   gpc1_1 gpc885 (
      {stage0_20[114]},
      {stage1_20[58]}
   );
   gpc1_1 gpc886 (
      {stage0_20[115]},
      {stage1_20[59]}
   );
   gpc1_1 gpc887 (
      {stage0_20[116]},
      {stage1_20[60]}
   );
   gpc1_1 gpc888 (
      {stage0_20[117]},
      {stage1_20[61]}
   );
   gpc1_1 gpc889 (
      {stage0_20[118]},
      {stage1_20[62]}
   );
   gpc1_1 gpc890 (
      {stage0_20[119]},
      {stage1_20[63]}
   );
   gpc1_1 gpc891 (
      {stage0_20[120]},
      {stage1_20[64]}
   );
   gpc1_1 gpc892 (
      {stage0_20[121]},
      {stage1_20[65]}
   );
   gpc1_1 gpc893 (
      {stage0_20[122]},
      {stage1_20[66]}
   );
   gpc1_1 gpc894 (
      {stage0_20[123]},
      {stage1_20[67]}
   );
   gpc1_1 gpc895 (
      {stage0_20[124]},
      {stage1_20[68]}
   );
   gpc1_1 gpc896 (
      {stage0_20[125]},
      {stage1_20[69]}
   );
   gpc1_1 gpc897 (
      {stage0_20[126]},
      {stage1_20[70]}
   );
   gpc1_1 gpc898 (
      {stage0_20[127]},
      {stage1_20[71]}
   );
   gpc1_1 gpc899 (
      {stage0_21[121]},
      {stage1_21[48]}
   );
   gpc1_1 gpc900 (
      {stage0_21[122]},
      {stage1_21[49]}
   );
   gpc1_1 gpc901 (
      {stage0_21[123]},
      {stage1_21[50]}
   );
   gpc1_1 gpc902 (
      {stage0_21[124]},
      {stage1_21[51]}
   );
   gpc1_1 gpc903 (
      {stage0_21[125]},
      {stage1_21[52]}
   );
   gpc1_1 gpc904 (
      {stage0_21[126]},
      {stage1_21[53]}
   );
   gpc1_1 gpc905 (
      {stage0_21[127]},
      {stage1_21[54]}
   );
   gpc1_1 gpc906 (
      {stage0_22[106]},
      {stage1_22[49]}
   );
   gpc1_1 gpc907 (
      {stage0_22[107]},
      {stage1_22[50]}
   );
   gpc1_1 gpc908 (
      {stage0_22[108]},
      {stage1_22[51]}
   );
   gpc1_1 gpc909 (
      {stage0_22[109]},
      {stage1_22[52]}
   );
   gpc1_1 gpc910 (
      {stage0_22[110]},
      {stage1_22[53]}
   );
   gpc1_1 gpc911 (
      {stage0_22[111]},
      {stage1_22[54]}
   );
   gpc1_1 gpc912 (
      {stage0_22[112]},
      {stage1_22[55]}
   );
   gpc1_1 gpc913 (
      {stage0_22[113]},
      {stage1_22[56]}
   );
   gpc1_1 gpc914 (
      {stage0_22[114]},
      {stage1_22[57]}
   );
   gpc1_1 gpc915 (
      {stage0_22[115]},
      {stage1_22[58]}
   );
   gpc1_1 gpc916 (
      {stage0_22[116]},
      {stage1_22[59]}
   );
   gpc1_1 gpc917 (
      {stage0_22[117]},
      {stage1_22[60]}
   );
   gpc1_1 gpc918 (
      {stage0_22[118]},
      {stage1_22[61]}
   );
   gpc1_1 gpc919 (
      {stage0_22[119]},
      {stage1_22[62]}
   );
   gpc1_1 gpc920 (
      {stage0_22[120]},
      {stage1_22[63]}
   );
   gpc1_1 gpc921 (
      {stage0_22[121]},
      {stage1_22[64]}
   );
   gpc1_1 gpc922 (
      {stage0_22[122]},
      {stage1_22[65]}
   );
   gpc1_1 gpc923 (
      {stage0_22[123]},
      {stage1_22[66]}
   );
   gpc1_1 gpc924 (
      {stage0_22[124]},
      {stage1_22[67]}
   );
   gpc1_1 gpc925 (
      {stage0_22[125]},
      {stage1_22[68]}
   );
   gpc1_1 gpc926 (
      {stage0_22[126]},
      {stage1_22[69]}
   );
   gpc1_1 gpc927 (
      {stage0_22[127]},
      {stage1_22[70]}
   );
   gpc1_1 gpc928 (
      {stage0_23[122]},
      {stage1_23[48]}
   );
   gpc1_1 gpc929 (
      {stage0_23[123]},
      {stage1_23[49]}
   );
   gpc1_1 gpc930 (
      {stage0_23[124]},
      {stage1_23[50]}
   );
   gpc1_1 gpc931 (
      {stage0_23[125]},
      {stage1_23[51]}
   );
   gpc1_1 gpc932 (
      {stage0_23[126]},
      {stage1_23[52]}
   );
   gpc1_1 gpc933 (
      {stage0_23[127]},
      {stage1_23[53]}
   );
   gpc1_1 gpc934 (
      {stage0_24[109]},
      {stage1_24[43]}
   );
   gpc1_1 gpc935 (
      {stage0_24[110]},
      {stage1_24[44]}
   );
   gpc1_1 gpc936 (
      {stage0_24[111]},
      {stage1_24[45]}
   );
   gpc1_1 gpc937 (
      {stage0_24[112]},
      {stage1_24[46]}
   );
   gpc1_1 gpc938 (
      {stage0_24[113]},
      {stage1_24[47]}
   );
   gpc1_1 gpc939 (
      {stage0_24[114]},
      {stage1_24[48]}
   );
   gpc1_1 gpc940 (
      {stage0_24[115]},
      {stage1_24[49]}
   );
   gpc1_1 gpc941 (
      {stage0_24[116]},
      {stage1_24[50]}
   );
   gpc1_1 gpc942 (
      {stage0_24[117]},
      {stage1_24[51]}
   );
   gpc1_1 gpc943 (
      {stage0_24[118]},
      {stage1_24[52]}
   );
   gpc1_1 gpc944 (
      {stage0_24[119]},
      {stage1_24[53]}
   );
   gpc1_1 gpc945 (
      {stage0_24[120]},
      {stage1_24[54]}
   );
   gpc1_1 gpc946 (
      {stage0_24[121]},
      {stage1_24[55]}
   );
   gpc1_1 gpc947 (
      {stage0_24[122]},
      {stage1_24[56]}
   );
   gpc1_1 gpc948 (
      {stage0_24[123]},
      {stage1_24[57]}
   );
   gpc1_1 gpc949 (
      {stage0_24[124]},
      {stage1_24[58]}
   );
   gpc1_1 gpc950 (
      {stage0_24[125]},
      {stage1_24[59]}
   );
   gpc1_1 gpc951 (
      {stage0_24[126]},
      {stage1_24[60]}
   );
   gpc1_1 gpc952 (
      {stage0_24[127]},
      {stage1_24[61]}
   );
   gpc1_1 gpc953 (
      {stage0_25[114]},
      {stage1_25[47]}
   );
   gpc1_1 gpc954 (
      {stage0_25[115]},
      {stage1_25[48]}
   );
   gpc1_1 gpc955 (
      {stage0_25[116]},
      {stage1_25[49]}
   );
   gpc1_1 gpc956 (
      {stage0_25[117]},
      {stage1_25[50]}
   );
   gpc1_1 gpc957 (
      {stage0_25[118]},
      {stage1_25[51]}
   );
   gpc1_1 gpc958 (
      {stage0_25[119]},
      {stage1_25[52]}
   );
   gpc1_1 gpc959 (
      {stage0_25[120]},
      {stage1_25[53]}
   );
   gpc1_1 gpc960 (
      {stage0_25[121]},
      {stage1_25[54]}
   );
   gpc1_1 gpc961 (
      {stage0_25[122]},
      {stage1_25[55]}
   );
   gpc1_1 gpc962 (
      {stage0_25[123]},
      {stage1_25[56]}
   );
   gpc1_1 gpc963 (
      {stage0_25[124]},
      {stage1_25[57]}
   );
   gpc1_1 gpc964 (
      {stage0_25[125]},
      {stage1_25[58]}
   );
   gpc1_1 gpc965 (
      {stage0_25[126]},
      {stage1_25[59]}
   );
   gpc1_1 gpc966 (
      {stage0_25[127]},
      {stage1_25[60]}
   );
   gpc1_1 gpc967 (
      {stage0_26[93]},
      {stage1_26[49]}
   );
   gpc1_1 gpc968 (
      {stage0_26[94]},
      {stage1_26[50]}
   );
   gpc1_1 gpc969 (
      {stage0_26[95]},
      {stage1_26[51]}
   );
   gpc1_1 gpc970 (
      {stage0_26[96]},
      {stage1_26[52]}
   );
   gpc1_1 gpc971 (
      {stage0_26[97]},
      {stage1_26[53]}
   );
   gpc1_1 gpc972 (
      {stage0_26[98]},
      {stage1_26[54]}
   );
   gpc1_1 gpc973 (
      {stage0_26[99]},
      {stage1_26[55]}
   );
   gpc1_1 gpc974 (
      {stage0_26[100]},
      {stage1_26[56]}
   );
   gpc1_1 gpc975 (
      {stage0_26[101]},
      {stage1_26[57]}
   );
   gpc1_1 gpc976 (
      {stage0_26[102]},
      {stage1_26[58]}
   );
   gpc1_1 gpc977 (
      {stage0_26[103]},
      {stage1_26[59]}
   );
   gpc1_1 gpc978 (
      {stage0_26[104]},
      {stage1_26[60]}
   );
   gpc1_1 gpc979 (
      {stage0_26[105]},
      {stage1_26[61]}
   );
   gpc1_1 gpc980 (
      {stage0_26[106]},
      {stage1_26[62]}
   );
   gpc1_1 gpc981 (
      {stage0_26[107]},
      {stage1_26[63]}
   );
   gpc1_1 gpc982 (
      {stage0_26[108]},
      {stage1_26[64]}
   );
   gpc1_1 gpc983 (
      {stage0_26[109]},
      {stage1_26[65]}
   );
   gpc1_1 gpc984 (
      {stage0_26[110]},
      {stage1_26[66]}
   );
   gpc1_1 gpc985 (
      {stage0_26[111]},
      {stage1_26[67]}
   );
   gpc1_1 gpc986 (
      {stage0_26[112]},
      {stage1_26[68]}
   );
   gpc1_1 gpc987 (
      {stage0_26[113]},
      {stage1_26[69]}
   );
   gpc1_1 gpc988 (
      {stage0_26[114]},
      {stage1_26[70]}
   );
   gpc1_1 gpc989 (
      {stage0_26[115]},
      {stage1_26[71]}
   );
   gpc1_1 gpc990 (
      {stage0_26[116]},
      {stage1_26[72]}
   );
   gpc1_1 gpc991 (
      {stage0_26[117]},
      {stage1_26[73]}
   );
   gpc1_1 gpc992 (
      {stage0_26[118]},
      {stage1_26[74]}
   );
   gpc1_1 gpc993 (
      {stage0_26[119]},
      {stage1_26[75]}
   );
   gpc1_1 gpc994 (
      {stage0_26[120]},
      {stage1_26[76]}
   );
   gpc1_1 gpc995 (
      {stage0_26[121]},
      {stage1_26[77]}
   );
   gpc1_1 gpc996 (
      {stage0_26[122]},
      {stage1_26[78]}
   );
   gpc1_1 gpc997 (
      {stage0_26[123]},
      {stage1_26[79]}
   );
   gpc1_1 gpc998 (
      {stage0_26[124]},
      {stage1_26[80]}
   );
   gpc1_1 gpc999 (
      {stage0_26[125]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1000 (
      {stage0_26[126]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1001 (
      {stage0_26[127]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1002 (
      {stage0_27[114]},
      {stage1_27[42]}
   );
   gpc1_1 gpc1003 (
      {stage0_27[115]},
      {stage1_27[43]}
   );
   gpc1_1 gpc1004 (
      {stage0_27[116]},
      {stage1_27[44]}
   );
   gpc1_1 gpc1005 (
      {stage0_27[117]},
      {stage1_27[45]}
   );
   gpc1_1 gpc1006 (
      {stage0_27[118]},
      {stage1_27[46]}
   );
   gpc1_1 gpc1007 (
      {stage0_27[119]},
      {stage1_27[47]}
   );
   gpc1_1 gpc1008 (
      {stage0_27[120]},
      {stage1_27[48]}
   );
   gpc1_1 gpc1009 (
      {stage0_27[121]},
      {stage1_27[49]}
   );
   gpc1_1 gpc1010 (
      {stage0_27[122]},
      {stage1_27[50]}
   );
   gpc1_1 gpc1011 (
      {stage0_27[123]},
      {stage1_27[51]}
   );
   gpc1_1 gpc1012 (
      {stage0_27[124]},
      {stage1_27[52]}
   );
   gpc1_1 gpc1013 (
      {stage0_27[125]},
      {stage1_27[53]}
   );
   gpc1_1 gpc1014 (
      {stage0_27[126]},
      {stage1_27[54]}
   );
   gpc1_1 gpc1015 (
      {stage0_27[127]},
      {stage1_27[55]}
   );
   gpc1_1 gpc1016 (
      {stage0_28[126]},
      {stage1_28[46]}
   );
   gpc1_1 gpc1017 (
      {stage0_28[127]},
      {stage1_28[47]}
   );
   gpc1_1 gpc1018 (
      {stage0_29[99]},
      {stage1_29[51]}
   );
   gpc1_1 gpc1019 (
      {stage0_29[100]},
      {stage1_29[52]}
   );
   gpc1_1 gpc1020 (
      {stage0_29[101]},
      {stage1_29[53]}
   );
   gpc1_1 gpc1021 (
      {stage0_29[102]},
      {stage1_29[54]}
   );
   gpc1_1 gpc1022 (
      {stage0_29[103]},
      {stage1_29[55]}
   );
   gpc1_1 gpc1023 (
      {stage0_29[104]},
      {stage1_29[56]}
   );
   gpc1_1 gpc1024 (
      {stage0_29[105]},
      {stage1_29[57]}
   );
   gpc1_1 gpc1025 (
      {stage0_29[106]},
      {stage1_29[58]}
   );
   gpc1_1 gpc1026 (
      {stage0_29[107]},
      {stage1_29[59]}
   );
   gpc1_1 gpc1027 (
      {stage0_29[108]},
      {stage1_29[60]}
   );
   gpc1_1 gpc1028 (
      {stage0_29[109]},
      {stage1_29[61]}
   );
   gpc1_1 gpc1029 (
      {stage0_29[110]},
      {stage1_29[62]}
   );
   gpc1_1 gpc1030 (
      {stage0_29[111]},
      {stage1_29[63]}
   );
   gpc1_1 gpc1031 (
      {stage0_29[112]},
      {stage1_29[64]}
   );
   gpc1_1 gpc1032 (
      {stage0_29[113]},
      {stage1_29[65]}
   );
   gpc1_1 gpc1033 (
      {stage0_29[114]},
      {stage1_29[66]}
   );
   gpc1_1 gpc1034 (
      {stage0_29[115]},
      {stage1_29[67]}
   );
   gpc1_1 gpc1035 (
      {stage0_29[116]},
      {stage1_29[68]}
   );
   gpc1_1 gpc1036 (
      {stage0_29[117]},
      {stage1_29[69]}
   );
   gpc1_1 gpc1037 (
      {stage0_29[118]},
      {stage1_29[70]}
   );
   gpc1_1 gpc1038 (
      {stage0_29[119]},
      {stage1_29[71]}
   );
   gpc1_1 gpc1039 (
      {stage0_29[120]},
      {stage1_29[72]}
   );
   gpc1_1 gpc1040 (
      {stage0_29[121]},
      {stage1_29[73]}
   );
   gpc1_1 gpc1041 (
      {stage0_29[122]},
      {stage1_29[74]}
   );
   gpc1_1 gpc1042 (
      {stage0_29[123]},
      {stage1_29[75]}
   );
   gpc1_1 gpc1043 (
      {stage0_29[124]},
      {stage1_29[76]}
   );
   gpc1_1 gpc1044 (
      {stage0_29[125]},
      {stage1_29[77]}
   );
   gpc1_1 gpc1045 (
      {stage0_29[126]},
      {stage1_29[78]}
   );
   gpc1_1 gpc1046 (
      {stage0_29[127]},
      {stage1_29[79]}
   );
   gpc1_1 gpc1047 (
      {stage0_30[99]},
      {stage1_30[43]}
   );
   gpc1_1 gpc1048 (
      {stage0_30[100]},
      {stage1_30[44]}
   );
   gpc1_1 gpc1049 (
      {stage0_30[101]},
      {stage1_30[45]}
   );
   gpc1_1 gpc1050 (
      {stage0_30[102]},
      {stage1_30[46]}
   );
   gpc1_1 gpc1051 (
      {stage0_30[103]},
      {stage1_30[47]}
   );
   gpc1_1 gpc1052 (
      {stage0_30[104]},
      {stage1_30[48]}
   );
   gpc1_1 gpc1053 (
      {stage0_30[105]},
      {stage1_30[49]}
   );
   gpc1_1 gpc1054 (
      {stage0_30[106]},
      {stage1_30[50]}
   );
   gpc1_1 gpc1055 (
      {stage0_30[107]},
      {stage1_30[51]}
   );
   gpc1_1 gpc1056 (
      {stage0_30[108]},
      {stage1_30[52]}
   );
   gpc1_1 gpc1057 (
      {stage0_30[109]},
      {stage1_30[53]}
   );
   gpc1_1 gpc1058 (
      {stage0_30[110]},
      {stage1_30[54]}
   );
   gpc1_1 gpc1059 (
      {stage0_30[111]},
      {stage1_30[55]}
   );
   gpc1_1 gpc1060 (
      {stage0_30[112]},
      {stage1_30[56]}
   );
   gpc1_1 gpc1061 (
      {stage0_30[113]},
      {stage1_30[57]}
   );
   gpc1_1 gpc1062 (
      {stage0_30[114]},
      {stage1_30[58]}
   );
   gpc1_1 gpc1063 (
      {stage0_30[115]},
      {stage1_30[59]}
   );
   gpc1_1 gpc1064 (
      {stage0_30[116]},
      {stage1_30[60]}
   );
   gpc1_1 gpc1065 (
      {stage0_30[117]},
      {stage1_30[61]}
   );
   gpc1_1 gpc1066 (
      {stage0_30[118]},
      {stage1_30[62]}
   );
   gpc1_1 gpc1067 (
      {stage0_30[119]},
      {stage1_30[63]}
   );
   gpc1_1 gpc1068 (
      {stage0_30[120]},
      {stage1_30[64]}
   );
   gpc1_1 gpc1069 (
      {stage0_30[121]},
      {stage1_30[65]}
   );
   gpc1_1 gpc1070 (
      {stage0_30[122]},
      {stage1_30[66]}
   );
   gpc1_1 gpc1071 (
      {stage0_30[123]},
      {stage1_30[67]}
   );
   gpc1_1 gpc1072 (
      {stage0_30[124]},
      {stage1_30[68]}
   );
   gpc1_1 gpc1073 (
      {stage0_30[125]},
      {stage1_30[69]}
   );
   gpc1_1 gpc1074 (
      {stage0_30[126]},
      {stage1_30[70]}
   );
   gpc1_1 gpc1075 (
      {stage0_30[127]},
      {stage1_30[71]}
   );
   gpc1_1 gpc1076 (
      {stage0_31[109]},
      {stage1_31[41]}
   );
   gpc1_1 gpc1077 (
      {stage0_31[110]},
      {stage1_31[42]}
   );
   gpc1_1 gpc1078 (
      {stage0_31[111]},
      {stage1_31[43]}
   );
   gpc1_1 gpc1079 (
      {stage0_31[112]},
      {stage1_31[44]}
   );
   gpc1_1 gpc1080 (
      {stage0_31[113]},
      {stage1_31[45]}
   );
   gpc1_1 gpc1081 (
      {stage0_31[114]},
      {stage1_31[46]}
   );
   gpc1_1 gpc1082 (
      {stage0_31[115]},
      {stage1_31[47]}
   );
   gpc1_1 gpc1083 (
      {stage0_31[116]},
      {stage1_31[48]}
   );
   gpc1_1 gpc1084 (
      {stage0_31[117]},
      {stage1_31[49]}
   );
   gpc1_1 gpc1085 (
      {stage0_31[118]},
      {stage1_31[50]}
   );
   gpc1_1 gpc1086 (
      {stage0_31[119]},
      {stage1_31[51]}
   );
   gpc1_1 gpc1087 (
      {stage0_31[120]},
      {stage1_31[52]}
   );
   gpc1_1 gpc1088 (
      {stage0_31[121]},
      {stage1_31[53]}
   );
   gpc1_1 gpc1089 (
      {stage0_31[122]},
      {stage1_31[54]}
   );
   gpc1_1 gpc1090 (
      {stage0_31[123]},
      {stage1_31[55]}
   );
   gpc1_1 gpc1091 (
      {stage0_31[124]},
      {stage1_31[56]}
   );
   gpc1_1 gpc1092 (
      {stage0_31[125]},
      {stage1_31[57]}
   );
   gpc1_1 gpc1093 (
      {stage0_31[126]},
      {stage1_31[58]}
   );
   gpc1_1 gpc1094 (
      {stage0_31[127]},
      {stage1_31[59]}
   );
   gpc1_1 gpc1095 (
      {stage0_32[93]},
      {stage1_32[48]}
   );
   gpc1_1 gpc1096 (
      {stage0_32[94]},
      {stage1_32[49]}
   );
   gpc1_1 gpc1097 (
      {stage0_32[95]},
      {stage1_32[50]}
   );
   gpc1_1 gpc1098 (
      {stage0_32[96]},
      {stage1_32[51]}
   );
   gpc1_1 gpc1099 (
      {stage0_32[97]},
      {stage1_32[52]}
   );
   gpc1_1 gpc1100 (
      {stage0_32[98]},
      {stage1_32[53]}
   );
   gpc1_1 gpc1101 (
      {stage0_32[99]},
      {stage1_32[54]}
   );
   gpc1_1 gpc1102 (
      {stage0_32[100]},
      {stage1_32[55]}
   );
   gpc1_1 gpc1103 (
      {stage0_32[101]},
      {stage1_32[56]}
   );
   gpc1_1 gpc1104 (
      {stage0_32[102]},
      {stage1_32[57]}
   );
   gpc1_1 gpc1105 (
      {stage0_32[103]},
      {stage1_32[58]}
   );
   gpc1_1 gpc1106 (
      {stage0_32[104]},
      {stage1_32[59]}
   );
   gpc1_1 gpc1107 (
      {stage0_32[105]},
      {stage1_32[60]}
   );
   gpc1_1 gpc1108 (
      {stage0_32[106]},
      {stage1_32[61]}
   );
   gpc1_1 gpc1109 (
      {stage0_32[107]},
      {stage1_32[62]}
   );
   gpc1_1 gpc1110 (
      {stage0_32[108]},
      {stage1_32[63]}
   );
   gpc1_1 gpc1111 (
      {stage0_32[109]},
      {stage1_32[64]}
   );
   gpc1_1 gpc1112 (
      {stage0_32[110]},
      {stage1_32[65]}
   );
   gpc1_1 gpc1113 (
      {stage0_32[111]},
      {stage1_32[66]}
   );
   gpc1_1 gpc1114 (
      {stage0_32[112]},
      {stage1_32[67]}
   );
   gpc1_1 gpc1115 (
      {stage0_32[113]},
      {stage1_32[68]}
   );
   gpc1_1 gpc1116 (
      {stage0_32[114]},
      {stage1_32[69]}
   );
   gpc1_1 gpc1117 (
      {stage0_32[115]},
      {stage1_32[70]}
   );
   gpc1_1 gpc1118 (
      {stage0_32[116]},
      {stage1_32[71]}
   );
   gpc1_1 gpc1119 (
      {stage0_32[117]},
      {stage1_32[72]}
   );
   gpc1_1 gpc1120 (
      {stage0_32[118]},
      {stage1_32[73]}
   );
   gpc1_1 gpc1121 (
      {stage0_32[119]},
      {stage1_32[74]}
   );
   gpc1_1 gpc1122 (
      {stage0_32[120]},
      {stage1_32[75]}
   );
   gpc1_1 gpc1123 (
      {stage0_32[121]},
      {stage1_32[76]}
   );
   gpc1_1 gpc1124 (
      {stage0_32[122]},
      {stage1_32[77]}
   );
   gpc1_1 gpc1125 (
      {stage0_32[123]},
      {stage1_32[78]}
   );
   gpc1_1 gpc1126 (
      {stage0_32[124]},
      {stage1_32[79]}
   );
   gpc1_1 gpc1127 (
      {stage0_32[125]},
      {stage1_32[80]}
   );
   gpc1_1 gpc1128 (
      {stage0_32[126]},
      {stage1_32[81]}
   );
   gpc1_1 gpc1129 (
      {stage0_32[127]},
      {stage1_32[82]}
   );
   gpc1_1 gpc1130 (
      {stage0_33[109]},
      {stage1_33[44]}
   );
   gpc1_1 gpc1131 (
      {stage0_33[110]},
      {stage1_33[45]}
   );
   gpc1_1 gpc1132 (
      {stage0_33[111]},
      {stage1_33[46]}
   );
   gpc1_1 gpc1133 (
      {stage0_33[112]},
      {stage1_33[47]}
   );
   gpc1_1 gpc1134 (
      {stage0_33[113]},
      {stage1_33[48]}
   );
   gpc1_1 gpc1135 (
      {stage0_33[114]},
      {stage1_33[49]}
   );
   gpc1_1 gpc1136 (
      {stage0_33[115]},
      {stage1_33[50]}
   );
   gpc1_1 gpc1137 (
      {stage0_33[116]},
      {stage1_33[51]}
   );
   gpc1_1 gpc1138 (
      {stage0_33[117]},
      {stage1_33[52]}
   );
   gpc1_1 gpc1139 (
      {stage0_33[118]},
      {stage1_33[53]}
   );
   gpc1_1 gpc1140 (
      {stage0_33[119]},
      {stage1_33[54]}
   );
   gpc1_1 gpc1141 (
      {stage0_33[120]},
      {stage1_33[55]}
   );
   gpc1_1 gpc1142 (
      {stage0_33[121]},
      {stage1_33[56]}
   );
   gpc1_1 gpc1143 (
      {stage0_33[122]},
      {stage1_33[57]}
   );
   gpc1_1 gpc1144 (
      {stage0_33[123]},
      {stage1_33[58]}
   );
   gpc1_1 gpc1145 (
      {stage0_33[124]},
      {stage1_33[59]}
   );
   gpc1_1 gpc1146 (
      {stage0_33[125]},
      {stage1_33[60]}
   );
   gpc1_1 gpc1147 (
      {stage0_33[126]},
      {stage1_33[61]}
   );
   gpc1_1 gpc1148 (
      {stage0_33[127]},
      {stage1_33[62]}
   );
   gpc1_1 gpc1149 (
      {stage0_34[97]},
      {stage1_34[37]}
   );
   gpc1_1 gpc1150 (
      {stage0_34[98]},
      {stage1_34[38]}
   );
   gpc1_1 gpc1151 (
      {stage0_34[99]},
      {stage1_34[39]}
   );
   gpc1_1 gpc1152 (
      {stage0_34[100]},
      {stage1_34[40]}
   );
   gpc1_1 gpc1153 (
      {stage0_34[101]},
      {stage1_34[41]}
   );
   gpc1_1 gpc1154 (
      {stage0_34[102]},
      {stage1_34[42]}
   );
   gpc1_1 gpc1155 (
      {stage0_34[103]},
      {stage1_34[43]}
   );
   gpc1_1 gpc1156 (
      {stage0_34[104]},
      {stage1_34[44]}
   );
   gpc1_1 gpc1157 (
      {stage0_34[105]},
      {stage1_34[45]}
   );
   gpc1_1 gpc1158 (
      {stage0_34[106]},
      {stage1_34[46]}
   );
   gpc1_1 gpc1159 (
      {stage0_34[107]},
      {stage1_34[47]}
   );
   gpc1_1 gpc1160 (
      {stage0_34[108]},
      {stage1_34[48]}
   );
   gpc1_1 gpc1161 (
      {stage0_34[109]},
      {stage1_34[49]}
   );
   gpc1_1 gpc1162 (
      {stage0_34[110]},
      {stage1_34[50]}
   );
   gpc1_1 gpc1163 (
      {stage0_34[111]},
      {stage1_34[51]}
   );
   gpc1_1 gpc1164 (
      {stage0_34[112]},
      {stage1_34[52]}
   );
   gpc1_1 gpc1165 (
      {stage0_34[113]},
      {stage1_34[53]}
   );
   gpc1_1 gpc1166 (
      {stage0_34[114]},
      {stage1_34[54]}
   );
   gpc1_1 gpc1167 (
      {stage0_34[115]},
      {stage1_34[55]}
   );
   gpc1_1 gpc1168 (
      {stage0_34[116]},
      {stage1_34[56]}
   );
   gpc1_1 gpc1169 (
      {stage0_34[117]},
      {stage1_34[57]}
   );
   gpc1_1 gpc1170 (
      {stage0_34[118]},
      {stage1_34[58]}
   );
   gpc1_1 gpc1171 (
      {stage0_34[119]},
      {stage1_34[59]}
   );
   gpc1_1 gpc1172 (
      {stage0_34[120]},
      {stage1_34[60]}
   );
   gpc1_1 gpc1173 (
      {stage0_34[121]},
      {stage1_34[61]}
   );
   gpc1_1 gpc1174 (
      {stage0_34[122]},
      {stage1_34[62]}
   );
   gpc1_1 gpc1175 (
      {stage0_34[123]},
      {stage1_34[63]}
   );
   gpc1_1 gpc1176 (
      {stage0_34[124]},
      {stage1_34[64]}
   );
   gpc1_1 gpc1177 (
      {stage0_34[125]},
      {stage1_34[65]}
   );
   gpc1_1 gpc1178 (
      {stage0_34[126]},
      {stage1_34[66]}
   );
   gpc1_1 gpc1179 (
      {stage0_34[127]},
      {stage1_34[67]}
   );
   gpc1_1 gpc1180 (
      {stage0_35[127]},
      {stage1_35[47]}
   );
   gpc1_1 gpc1181 (
      {stage0_36[120]},
      {stage1_36[53]}
   );
   gpc1_1 gpc1182 (
      {stage0_36[121]},
      {stage1_36[54]}
   );
   gpc1_1 gpc1183 (
      {stage0_36[122]},
      {stage1_36[55]}
   );
   gpc1_1 gpc1184 (
      {stage0_36[123]},
      {stage1_36[56]}
   );
   gpc1_1 gpc1185 (
      {stage0_36[124]},
      {stage1_36[57]}
   );
   gpc1_1 gpc1186 (
      {stage0_36[125]},
      {stage1_36[58]}
   );
   gpc1_1 gpc1187 (
      {stage0_36[126]},
      {stage1_36[59]}
   );
   gpc1_1 gpc1188 (
      {stage0_36[127]},
      {stage1_36[60]}
   );
   gpc1_1 gpc1189 (
      {stage0_37[72]},
      {stage1_37[41]}
   );
   gpc1_1 gpc1190 (
      {stage0_37[73]},
      {stage1_37[42]}
   );
   gpc1_1 gpc1191 (
      {stage0_37[74]},
      {stage1_37[43]}
   );
   gpc1_1 gpc1192 (
      {stage0_37[75]},
      {stage1_37[44]}
   );
   gpc1_1 gpc1193 (
      {stage0_37[76]},
      {stage1_37[45]}
   );
   gpc1_1 gpc1194 (
      {stage0_37[77]},
      {stage1_37[46]}
   );
   gpc1_1 gpc1195 (
      {stage0_37[78]},
      {stage1_37[47]}
   );
   gpc1_1 gpc1196 (
      {stage0_37[79]},
      {stage1_37[48]}
   );
   gpc1_1 gpc1197 (
      {stage0_37[80]},
      {stage1_37[49]}
   );
   gpc1_1 gpc1198 (
      {stage0_37[81]},
      {stage1_37[50]}
   );
   gpc1_1 gpc1199 (
      {stage0_37[82]},
      {stage1_37[51]}
   );
   gpc1_1 gpc1200 (
      {stage0_37[83]},
      {stage1_37[52]}
   );
   gpc1_1 gpc1201 (
      {stage0_37[84]},
      {stage1_37[53]}
   );
   gpc1_1 gpc1202 (
      {stage0_37[85]},
      {stage1_37[54]}
   );
   gpc1_1 gpc1203 (
      {stage0_37[86]},
      {stage1_37[55]}
   );
   gpc1_1 gpc1204 (
      {stage0_37[87]},
      {stage1_37[56]}
   );
   gpc1_1 gpc1205 (
      {stage0_37[88]},
      {stage1_37[57]}
   );
   gpc1_1 gpc1206 (
      {stage0_37[89]},
      {stage1_37[58]}
   );
   gpc1_1 gpc1207 (
      {stage0_37[90]},
      {stage1_37[59]}
   );
   gpc1_1 gpc1208 (
      {stage0_37[91]},
      {stage1_37[60]}
   );
   gpc1_1 gpc1209 (
      {stage0_37[92]},
      {stage1_37[61]}
   );
   gpc1_1 gpc1210 (
      {stage0_37[93]},
      {stage1_37[62]}
   );
   gpc1_1 gpc1211 (
      {stage0_37[94]},
      {stage1_37[63]}
   );
   gpc1_1 gpc1212 (
      {stage0_37[95]},
      {stage1_37[64]}
   );
   gpc1_1 gpc1213 (
      {stage0_37[96]},
      {stage1_37[65]}
   );
   gpc1_1 gpc1214 (
      {stage0_37[97]},
      {stage1_37[66]}
   );
   gpc1_1 gpc1215 (
      {stage0_37[98]},
      {stage1_37[67]}
   );
   gpc1_1 gpc1216 (
      {stage0_37[99]},
      {stage1_37[68]}
   );
   gpc1_1 gpc1217 (
      {stage0_37[100]},
      {stage1_37[69]}
   );
   gpc1_1 gpc1218 (
      {stage0_37[101]},
      {stage1_37[70]}
   );
   gpc1_1 gpc1219 (
      {stage0_37[102]},
      {stage1_37[71]}
   );
   gpc1_1 gpc1220 (
      {stage0_37[103]},
      {stage1_37[72]}
   );
   gpc1_1 gpc1221 (
      {stage0_37[104]},
      {stage1_37[73]}
   );
   gpc1_1 gpc1222 (
      {stage0_37[105]},
      {stage1_37[74]}
   );
   gpc1_1 gpc1223 (
      {stage0_37[106]},
      {stage1_37[75]}
   );
   gpc1_1 gpc1224 (
      {stage0_37[107]},
      {stage1_37[76]}
   );
   gpc1_1 gpc1225 (
      {stage0_37[108]},
      {stage1_37[77]}
   );
   gpc1_1 gpc1226 (
      {stage0_37[109]},
      {stage1_37[78]}
   );
   gpc1_1 gpc1227 (
      {stage0_37[110]},
      {stage1_37[79]}
   );
   gpc1_1 gpc1228 (
      {stage0_37[111]},
      {stage1_37[80]}
   );
   gpc1_1 gpc1229 (
      {stage0_37[112]},
      {stage1_37[81]}
   );
   gpc1_1 gpc1230 (
      {stage0_37[113]},
      {stage1_37[82]}
   );
   gpc1_1 gpc1231 (
      {stage0_37[114]},
      {stage1_37[83]}
   );
   gpc1_1 gpc1232 (
      {stage0_37[115]},
      {stage1_37[84]}
   );
   gpc1_1 gpc1233 (
      {stage0_37[116]},
      {stage1_37[85]}
   );
   gpc1_1 gpc1234 (
      {stage0_37[117]},
      {stage1_37[86]}
   );
   gpc1_1 gpc1235 (
      {stage0_37[118]},
      {stage1_37[87]}
   );
   gpc1_1 gpc1236 (
      {stage0_37[119]},
      {stage1_37[88]}
   );
   gpc1_1 gpc1237 (
      {stage0_37[120]},
      {stage1_37[89]}
   );
   gpc1_1 gpc1238 (
      {stage0_37[121]},
      {stage1_37[90]}
   );
   gpc1_1 gpc1239 (
      {stage0_37[122]},
      {stage1_37[91]}
   );
   gpc1_1 gpc1240 (
      {stage0_37[123]},
      {stage1_37[92]}
   );
   gpc1_1 gpc1241 (
      {stage0_37[124]},
      {stage1_37[93]}
   );
   gpc1_1 gpc1242 (
      {stage0_37[125]},
      {stage1_37[94]}
   );
   gpc1_1 gpc1243 (
      {stage0_37[126]},
      {stage1_37[95]}
   );
   gpc1_1 gpc1244 (
      {stage0_37[127]},
      {stage1_37[96]}
   );
   gpc1_1 gpc1245 (
      {stage0_38[120]},
      {stage1_38[36]}
   );
   gpc1_1 gpc1246 (
      {stage0_38[121]},
      {stage1_38[37]}
   );
   gpc1_1 gpc1247 (
      {stage0_38[122]},
      {stage1_38[38]}
   );
   gpc1_1 gpc1248 (
      {stage0_38[123]},
      {stage1_38[39]}
   );
   gpc1_1 gpc1249 (
      {stage0_38[124]},
      {stage1_38[40]}
   );
   gpc1_1 gpc1250 (
      {stage0_38[125]},
      {stage1_38[41]}
   );
   gpc1_1 gpc1251 (
      {stage0_38[126]},
      {stage1_38[42]}
   );
   gpc1_1 gpc1252 (
      {stage0_38[127]},
      {stage1_38[43]}
   );
   gpc1_1 gpc1253 (
      {stage0_39[83]},
      {stage1_39[48]}
   );
   gpc1_1 gpc1254 (
      {stage0_39[84]},
      {stage1_39[49]}
   );
   gpc1_1 gpc1255 (
      {stage0_39[85]},
      {stage1_39[50]}
   );
   gpc1_1 gpc1256 (
      {stage0_39[86]},
      {stage1_39[51]}
   );
   gpc1_1 gpc1257 (
      {stage0_39[87]},
      {stage1_39[52]}
   );
   gpc1_1 gpc1258 (
      {stage0_39[88]},
      {stage1_39[53]}
   );
   gpc1_1 gpc1259 (
      {stage0_39[89]},
      {stage1_39[54]}
   );
   gpc1_1 gpc1260 (
      {stage0_39[90]},
      {stage1_39[55]}
   );
   gpc1_1 gpc1261 (
      {stage0_39[91]},
      {stage1_39[56]}
   );
   gpc1_1 gpc1262 (
      {stage0_39[92]},
      {stage1_39[57]}
   );
   gpc1_1 gpc1263 (
      {stage0_39[93]},
      {stage1_39[58]}
   );
   gpc1_1 gpc1264 (
      {stage0_39[94]},
      {stage1_39[59]}
   );
   gpc1_1 gpc1265 (
      {stage0_39[95]},
      {stage1_39[60]}
   );
   gpc1_1 gpc1266 (
      {stage0_39[96]},
      {stage1_39[61]}
   );
   gpc1_1 gpc1267 (
      {stage0_39[97]},
      {stage1_39[62]}
   );
   gpc1_1 gpc1268 (
      {stage0_39[98]},
      {stage1_39[63]}
   );
   gpc1_1 gpc1269 (
      {stage0_39[99]},
      {stage1_39[64]}
   );
   gpc1_1 gpc1270 (
      {stage0_39[100]},
      {stage1_39[65]}
   );
   gpc1_1 gpc1271 (
      {stage0_39[101]},
      {stage1_39[66]}
   );
   gpc1_1 gpc1272 (
      {stage0_39[102]},
      {stage1_39[67]}
   );
   gpc1_1 gpc1273 (
      {stage0_39[103]},
      {stage1_39[68]}
   );
   gpc1_1 gpc1274 (
      {stage0_39[104]},
      {stage1_39[69]}
   );
   gpc1_1 gpc1275 (
      {stage0_39[105]},
      {stage1_39[70]}
   );
   gpc1_1 gpc1276 (
      {stage0_39[106]},
      {stage1_39[71]}
   );
   gpc1_1 gpc1277 (
      {stage0_39[107]},
      {stage1_39[72]}
   );
   gpc1_1 gpc1278 (
      {stage0_39[108]},
      {stage1_39[73]}
   );
   gpc1_1 gpc1279 (
      {stage0_39[109]},
      {stage1_39[74]}
   );
   gpc1_1 gpc1280 (
      {stage0_39[110]},
      {stage1_39[75]}
   );
   gpc1_1 gpc1281 (
      {stage0_39[111]},
      {stage1_39[76]}
   );
   gpc1_1 gpc1282 (
      {stage0_39[112]},
      {stage1_39[77]}
   );
   gpc1_1 gpc1283 (
      {stage0_39[113]},
      {stage1_39[78]}
   );
   gpc1_1 gpc1284 (
      {stage0_39[114]},
      {stage1_39[79]}
   );
   gpc1_1 gpc1285 (
      {stage0_39[115]},
      {stage1_39[80]}
   );
   gpc1_1 gpc1286 (
      {stage0_39[116]},
      {stage1_39[81]}
   );
   gpc1_1 gpc1287 (
      {stage0_39[117]},
      {stage1_39[82]}
   );
   gpc1_1 gpc1288 (
      {stage0_39[118]},
      {stage1_39[83]}
   );
   gpc1_1 gpc1289 (
      {stage0_39[119]},
      {stage1_39[84]}
   );
   gpc1_1 gpc1290 (
      {stage0_39[120]},
      {stage1_39[85]}
   );
   gpc1_1 gpc1291 (
      {stage0_39[121]},
      {stage1_39[86]}
   );
   gpc1_1 gpc1292 (
      {stage0_39[122]},
      {stage1_39[87]}
   );
   gpc1_1 gpc1293 (
      {stage0_39[123]},
      {stage1_39[88]}
   );
   gpc1_1 gpc1294 (
      {stage0_39[124]},
      {stage1_39[89]}
   );
   gpc1_1 gpc1295 (
      {stage0_39[125]},
      {stage1_39[90]}
   );
   gpc1_1 gpc1296 (
      {stage0_39[126]},
      {stage1_39[91]}
   );
   gpc1_1 gpc1297 (
      {stage0_39[127]},
      {stage1_39[92]}
   );
   gpc1_1 gpc1298 (
      {stage0_40[112]},
      {stage1_40[47]}
   );
   gpc1_1 gpc1299 (
      {stage0_40[113]},
      {stage1_40[48]}
   );
   gpc1_1 gpc1300 (
      {stage0_40[114]},
      {stage1_40[49]}
   );
   gpc1_1 gpc1301 (
      {stage0_40[115]},
      {stage1_40[50]}
   );
   gpc1_1 gpc1302 (
      {stage0_40[116]},
      {stage1_40[51]}
   );
   gpc1_1 gpc1303 (
      {stage0_40[117]},
      {stage1_40[52]}
   );
   gpc1_1 gpc1304 (
      {stage0_40[118]},
      {stage1_40[53]}
   );
   gpc1_1 gpc1305 (
      {stage0_40[119]},
      {stage1_40[54]}
   );
   gpc1_1 gpc1306 (
      {stage0_40[120]},
      {stage1_40[55]}
   );
   gpc1_1 gpc1307 (
      {stage0_40[121]},
      {stage1_40[56]}
   );
   gpc1_1 gpc1308 (
      {stage0_40[122]},
      {stage1_40[57]}
   );
   gpc1_1 gpc1309 (
      {stage0_40[123]},
      {stage1_40[58]}
   );
   gpc1_1 gpc1310 (
      {stage0_40[124]},
      {stage1_40[59]}
   );
   gpc1_1 gpc1311 (
      {stage0_40[125]},
      {stage1_40[60]}
   );
   gpc1_1 gpc1312 (
      {stage0_40[126]},
      {stage1_40[61]}
   );
   gpc1_1 gpc1313 (
      {stage0_40[127]},
      {stage1_40[62]}
   );
   gpc1_1 gpc1314 (
      {stage0_41[126]},
      {stage1_41[38]}
   );
   gpc1_1 gpc1315 (
      {stage0_41[127]},
      {stage1_41[39]}
   );
   gpc1_1 gpc1316 (
      {stage0_42[127]},
      {stage1_42[50]}
   );
   gpc1_1 gpc1317 (
      {stage0_43[104]},
      {stage1_43[55]}
   );
   gpc1_1 gpc1318 (
      {stage0_43[105]},
      {stage1_43[56]}
   );
   gpc1_1 gpc1319 (
      {stage0_43[106]},
      {stage1_43[57]}
   );
   gpc1_1 gpc1320 (
      {stage0_43[107]},
      {stage1_43[58]}
   );
   gpc1_1 gpc1321 (
      {stage0_43[108]},
      {stage1_43[59]}
   );
   gpc1_1 gpc1322 (
      {stage0_43[109]},
      {stage1_43[60]}
   );
   gpc1_1 gpc1323 (
      {stage0_43[110]},
      {stage1_43[61]}
   );
   gpc1_1 gpc1324 (
      {stage0_43[111]},
      {stage1_43[62]}
   );
   gpc1_1 gpc1325 (
      {stage0_43[112]},
      {stage1_43[63]}
   );
   gpc1_1 gpc1326 (
      {stage0_43[113]},
      {stage1_43[64]}
   );
   gpc1_1 gpc1327 (
      {stage0_43[114]},
      {stage1_43[65]}
   );
   gpc1_1 gpc1328 (
      {stage0_43[115]},
      {stage1_43[66]}
   );
   gpc1_1 gpc1329 (
      {stage0_43[116]},
      {stage1_43[67]}
   );
   gpc1_1 gpc1330 (
      {stage0_43[117]},
      {stage1_43[68]}
   );
   gpc1_1 gpc1331 (
      {stage0_43[118]},
      {stage1_43[69]}
   );
   gpc1_1 gpc1332 (
      {stage0_43[119]},
      {stage1_43[70]}
   );
   gpc1_1 gpc1333 (
      {stage0_43[120]},
      {stage1_43[71]}
   );
   gpc1_1 gpc1334 (
      {stage0_43[121]},
      {stage1_43[72]}
   );
   gpc1_1 gpc1335 (
      {stage0_43[122]},
      {stage1_43[73]}
   );
   gpc1_1 gpc1336 (
      {stage0_43[123]},
      {stage1_43[74]}
   );
   gpc1_1 gpc1337 (
      {stage0_43[124]},
      {stage1_43[75]}
   );
   gpc1_1 gpc1338 (
      {stage0_43[125]},
      {stage1_43[76]}
   );
   gpc1_1 gpc1339 (
      {stage0_43[126]},
      {stage1_43[77]}
   );
   gpc1_1 gpc1340 (
      {stage0_43[127]},
      {stage1_43[78]}
   );
   gpc1_1 gpc1341 (
      {stage0_44[125]},
      {stage1_44[47]}
   );
   gpc1_1 gpc1342 (
      {stage0_44[126]},
      {stage1_44[48]}
   );
   gpc1_1 gpc1343 (
      {stage0_44[127]},
      {stage1_44[49]}
   );
   gpc1_1 gpc1344 (
      {stage0_45[114]},
      {stage1_45[44]}
   );
   gpc1_1 gpc1345 (
      {stage0_45[115]},
      {stage1_45[45]}
   );
   gpc1_1 gpc1346 (
      {stage0_45[116]},
      {stage1_45[46]}
   );
   gpc1_1 gpc1347 (
      {stage0_45[117]},
      {stage1_45[47]}
   );
   gpc1_1 gpc1348 (
      {stage0_45[118]},
      {stage1_45[48]}
   );
   gpc1_1 gpc1349 (
      {stage0_45[119]},
      {stage1_45[49]}
   );
   gpc1_1 gpc1350 (
      {stage0_45[120]},
      {stage1_45[50]}
   );
   gpc1_1 gpc1351 (
      {stage0_45[121]},
      {stage1_45[51]}
   );
   gpc1_1 gpc1352 (
      {stage0_45[122]},
      {stage1_45[52]}
   );
   gpc1_1 gpc1353 (
      {stage0_45[123]},
      {stage1_45[53]}
   );
   gpc1_1 gpc1354 (
      {stage0_45[124]},
      {stage1_45[54]}
   );
   gpc1_1 gpc1355 (
      {stage0_45[125]},
      {stage1_45[55]}
   );
   gpc1_1 gpc1356 (
      {stage0_45[126]},
      {stage1_45[56]}
   );
   gpc1_1 gpc1357 (
      {stage0_45[127]},
      {stage1_45[57]}
   );
   gpc1_1 gpc1358 (
      {stage0_46[96]},
      {stage1_46[48]}
   );
   gpc1_1 gpc1359 (
      {stage0_46[97]},
      {stage1_46[49]}
   );
   gpc1_1 gpc1360 (
      {stage0_46[98]},
      {stage1_46[50]}
   );
   gpc1_1 gpc1361 (
      {stage0_46[99]},
      {stage1_46[51]}
   );
   gpc1_1 gpc1362 (
      {stage0_46[100]},
      {stage1_46[52]}
   );
   gpc1_1 gpc1363 (
      {stage0_46[101]},
      {stage1_46[53]}
   );
   gpc1_1 gpc1364 (
      {stage0_46[102]},
      {stage1_46[54]}
   );
   gpc1_1 gpc1365 (
      {stage0_46[103]},
      {stage1_46[55]}
   );
   gpc1_1 gpc1366 (
      {stage0_46[104]},
      {stage1_46[56]}
   );
   gpc1_1 gpc1367 (
      {stage0_46[105]},
      {stage1_46[57]}
   );
   gpc1_1 gpc1368 (
      {stage0_46[106]},
      {stage1_46[58]}
   );
   gpc1_1 gpc1369 (
      {stage0_46[107]},
      {stage1_46[59]}
   );
   gpc1_1 gpc1370 (
      {stage0_46[108]},
      {stage1_46[60]}
   );
   gpc1_1 gpc1371 (
      {stage0_46[109]},
      {stage1_46[61]}
   );
   gpc1_1 gpc1372 (
      {stage0_46[110]},
      {stage1_46[62]}
   );
   gpc1_1 gpc1373 (
      {stage0_46[111]},
      {stage1_46[63]}
   );
   gpc1_1 gpc1374 (
      {stage0_46[112]},
      {stage1_46[64]}
   );
   gpc1_1 gpc1375 (
      {stage0_46[113]},
      {stage1_46[65]}
   );
   gpc1_1 gpc1376 (
      {stage0_46[114]},
      {stage1_46[66]}
   );
   gpc1_1 gpc1377 (
      {stage0_46[115]},
      {stage1_46[67]}
   );
   gpc1_1 gpc1378 (
      {stage0_46[116]},
      {stage1_46[68]}
   );
   gpc1_1 gpc1379 (
      {stage0_46[117]},
      {stage1_46[69]}
   );
   gpc1_1 gpc1380 (
      {stage0_46[118]},
      {stage1_46[70]}
   );
   gpc1_1 gpc1381 (
      {stage0_46[119]},
      {stage1_46[71]}
   );
   gpc1_1 gpc1382 (
      {stage0_46[120]},
      {stage1_46[72]}
   );
   gpc1_1 gpc1383 (
      {stage0_46[121]},
      {stage1_46[73]}
   );
   gpc1_1 gpc1384 (
      {stage0_46[122]},
      {stage1_46[74]}
   );
   gpc1_1 gpc1385 (
      {stage0_46[123]},
      {stage1_46[75]}
   );
   gpc1_1 gpc1386 (
      {stage0_46[124]},
      {stage1_46[76]}
   );
   gpc1_1 gpc1387 (
      {stage0_46[125]},
      {stage1_46[77]}
   );
   gpc1_1 gpc1388 (
      {stage0_46[126]},
      {stage1_46[78]}
   );
   gpc1_1 gpc1389 (
      {stage0_46[127]},
      {stage1_46[79]}
   );
   gpc1_1 gpc1390 (
      {stage0_47[103]},
      {stage1_47[45]}
   );
   gpc1_1 gpc1391 (
      {stage0_47[104]},
      {stage1_47[46]}
   );
   gpc1_1 gpc1392 (
      {stage0_47[105]},
      {stage1_47[47]}
   );
   gpc1_1 gpc1393 (
      {stage0_47[106]},
      {stage1_47[48]}
   );
   gpc1_1 gpc1394 (
      {stage0_47[107]},
      {stage1_47[49]}
   );
   gpc1_1 gpc1395 (
      {stage0_47[108]},
      {stage1_47[50]}
   );
   gpc1_1 gpc1396 (
      {stage0_47[109]},
      {stage1_47[51]}
   );
   gpc1_1 gpc1397 (
      {stage0_47[110]},
      {stage1_47[52]}
   );
   gpc1_1 gpc1398 (
      {stage0_47[111]},
      {stage1_47[53]}
   );
   gpc1_1 gpc1399 (
      {stage0_47[112]},
      {stage1_47[54]}
   );
   gpc1_1 gpc1400 (
      {stage0_47[113]},
      {stage1_47[55]}
   );
   gpc1_1 gpc1401 (
      {stage0_47[114]},
      {stage1_47[56]}
   );
   gpc1_1 gpc1402 (
      {stage0_47[115]},
      {stage1_47[57]}
   );
   gpc1_1 gpc1403 (
      {stage0_47[116]},
      {stage1_47[58]}
   );
   gpc1_1 gpc1404 (
      {stage0_47[117]},
      {stage1_47[59]}
   );
   gpc1_1 gpc1405 (
      {stage0_47[118]},
      {stage1_47[60]}
   );
   gpc1_1 gpc1406 (
      {stage0_47[119]},
      {stage1_47[61]}
   );
   gpc1_1 gpc1407 (
      {stage0_47[120]},
      {stage1_47[62]}
   );
   gpc1_1 gpc1408 (
      {stage0_47[121]},
      {stage1_47[63]}
   );
   gpc1_1 gpc1409 (
      {stage0_47[122]},
      {stage1_47[64]}
   );
   gpc1_1 gpc1410 (
      {stage0_47[123]},
      {stage1_47[65]}
   );
   gpc1_1 gpc1411 (
      {stage0_47[124]},
      {stage1_47[66]}
   );
   gpc1_1 gpc1412 (
      {stage0_47[125]},
      {stage1_47[67]}
   );
   gpc1_1 gpc1413 (
      {stage0_47[126]},
      {stage1_47[68]}
   );
   gpc1_1 gpc1414 (
      {stage0_47[127]},
      {stage1_47[69]}
   );
   gpc1_1 gpc1415 (
      {stage0_48[127]},
      {stage1_48[45]}
   );
   gpc1_1 gpc1416 (
      {stage0_50[106]},
      {stage1_50[49]}
   );
   gpc1_1 gpc1417 (
      {stage0_50[107]},
      {stage1_50[50]}
   );
   gpc1_1 gpc1418 (
      {stage0_50[108]},
      {stage1_50[51]}
   );
   gpc1_1 gpc1419 (
      {stage0_50[109]},
      {stage1_50[52]}
   );
   gpc1_1 gpc1420 (
      {stage0_50[110]},
      {stage1_50[53]}
   );
   gpc1_1 gpc1421 (
      {stage0_50[111]},
      {stage1_50[54]}
   );
   gpc1_1 gpc1422 (
      {stage0_50[112]},
      {stage1_50[55]}
   );
   gpc1_1 gpc1423 (
      {stage0_50[113]},
      {stage1_50[56]}
   );
   gpc1_1 gpc1424 (
      {stage0_50[114]},
      {stage1_50[57]}
   );
   gpc1_1 gpc1425 (
      {stage0_50[115]},
      {stage1_50[58]}
   );
   gpc1_1 gpc1426 (
      {stage0_50[116]},
      {stage1_50[59]}
   );
   gpc1_1 gpc1427 (
      {stage0_50[117]},
      {stage1_50[60]}
   );
   gpc1_1 gpc1428 (
      {stage0_50[118]},
      {stage1_50[61]}
   );
   gpc1_1 gpc1429 (
      {stage0_50[119]},
      {stage1_50[62]}
   );
   gpc1_1 gpc1430 (
      {stage0_50[120]},
      {stage1_50[63]}
   );
   gpc1_1 gpc1431 (
      {stage0_50[121]},
      {stage1_50[64]}
   );
   gpc1_1 gpc1432 (
      {stage0_50[122]},
      {stage1_50[65]}
   );
   gpc1_1 gpc1433 (
      {stage0_50[123]},
      {stage1_50[66]}
   );
   gpc1_1 gpc1434 (
      {stage0_50[124]},
      {stage1_50[67]}
   );
   gpc1_1 gpc1435 (
      {stage0_50[125]},
      {stage1_50[68]}
   );
   gpc1_1 gpc1436 (
      {stage0_50[126]},
      {stage1_50[69]}
   );
   gpc1_1 gpc1437 (
      {stage0_50[127]},
      {stage1_50[70]}
   );
   gpc1_1 gpc1438 (
      {stage0_52[120]},
      {stage1_52[53]}
   );
   gpc1_1 gpc1439 (
      {stage0_52[121]},
      {stage1_52[54]}
   );
   gpc1_1 gpc1440 (
      {stage0_52[122]},
      {stage1_52[55]}
   );
   gpc1_1 gpc1441 (
      {stage0_52[123]},
      {stage1_52[56]}
   );
   gpc1_1 gpc1442 (
      {stage0_52[124]},
      {stage1_52[57]}
   );
   gpc1_1 gpc1443 (
      {stage0_52[125]},
      {stage1_52[58]}
   );
   gpc1_1 gpc1444 (
      {stage0_52[126]},
      {stage1_52[59]}
   );
   gpc1_1 gpc1445 (
      {stage0_52[127]},
      {stage1_52[60]}
   );
   gpc1_1 gpc1446 (
      {stage0_53[120]},
      {stage1_53[54]}
   );
   gpc1_1 gpc1447 (
      {stage0_53[121]},
      {stage1_53[55]}
   );
   gpc1_1 gpc1448 (
      {stage0_53[122]},
      {stage1_53[56]}
   );
   gpc1_1 gpc1449 (
      {stage0_53[123]},
      {stage1_53[57]}
   );
   gpc1_1 gpc1450 (
      {stage0_53[124]},
      {stage1_53[58]}
   );
   gpc1_1 gpc1451 (
      {stage0_53[125]},
      {stage1_53[59]}
   );
   gpc1_1 gpc1452 (
      {stage0_53[126]},
      {stage1_53[60]}
   );
   gpc1_1 gpc1453 (
      {stage0_53[127]},
      {stage1_53[61]}
   );
   gpc1_1 gpc1454 (
      {stage0_54[123]},
      {stage1_54[47]}
   );
   gpc1_1 gpc1455 (
      {stage0_54[124]},
      {stage1_54[48]}
   );
   gpc1_1 gpc1456 (
      {stage0_54[125]},
      {stage1_54[49]}
   );
   gpc1_1 gpc1457 (
      {stage0_54[126]},
      {stage1_54[50]}
   );
   gpc1_1 gpc1458 (
      {stage0_54[127]},
      {stage1_54[51]}
   );
   gpc1_1 gpc1459 (
      {stage0_55[108]},
      {stage1_55[48]}
   );
   gpc1_1 gpc1460 (
      {stage0_55[109]},
      {stage1_55[49]}
   );
   gpc1_1 gpc1461 (
      {stage0_55[110]},
      {stage1_55[50]}
   );
   gpc1_1 gpc1462 (
      {stage0_55[111]},
      {stage1_55[51]}
   );
   gpc1_1 gpc1463 (
      {stage0_55[112]},
      {stage1_55[52]}
   );
   gpc1_1 gpc1464 (
      {stage0_55[113]},
      {stage1_55[53]}
   );
   gpc1_1 gpc1465 (
      {stage0_55[114]},
      {stage1_55[54]}
   );
   gpc1_1 gpc1466 (
      {stage0_55[115]},
      {stage1_55[55]}
   );
   gpc1_1 gpc1467 (
      {stage0_55[116]},
      {stage1_55[56]}
   );
   gpc1_1 gpc1468 (
      {stage0_55[117]},
      {stage1_55[57]}
   );
   gpc1_1 gpc1469 (
      {stage0_55[118]},
      {stage1_55[58]}
   );
   gpc1_1 gpc1470 (
      {stage0_55[119]},
      {stage1_55[59]}
   );
   gpc1_1 gpc1471 (
      {stage0_55[120]},
      {stage1_55[60]}
   );
   gpc1_1 gpc1472 (
      {stage0_55[121]},
      {stage1_55[61]}
   );
   gpc1_1 gpc1473 (
      {stage0_55[122]},
      {stage1_55[62]}
   );
   gpc1_1 gpc1474 (
      {stage0_55[123]},
      {stage1_55[63]}
   );
   gpc1_1 gpc1475 (
      {stage0_55[124]},
      {stage1_55[64]}
   );
   gpc1_1 gpc1476 (
      {stage0_55[125]},
      {stage1_55[65]}
   );
   gpc1_1 gpc1477 (
      {stage0_55[126]},
      {stage1_55[66]}
   );
   gpc1_1 gpc1478 (
      {stage0_55[127]},
      {stage1_55[67]}
   );
   gpc1_1 gpc1479 (
      {stage0_56[122]},
      {stage1_56[51]}
   );
   gpc1_1 gpc1480 (
      {stage0_56[123]},
      {stage1_56[52]}
   );
   gpc1_1 gpc1481 (
      {stage0_56[124]},
      {stage1_56[53]}
   );
   gpc1_1 gpc1482 (
      {stage0_56[125]},
      {stage1_56[54]}
   );
   gpc1_1 gpc1483 (
      {stage0_56[126]},
      {stage1_56[55]}
   );
   gpc1_1 gpc1484 (
      {stage0_56[127]},
      {stage1_56[56]}
   );
   gpc1_1 gpc1485 (
      {stage0_57[122]},
      {stage1_57[52]}
   );
   gpc1_1 gpc1486 (
      {stage0_57[123]},
      {stage1_57[53]}
   );
   gpc1_1 gpc1487 (
      {stage0_57[124]},
      {stage1_57[54]}
   );
   gpc1_1 gpc1488 (
      {stage0_57[125]},
      {stage1_57[55]}
   );
   gpc1_1 gpc1489 (
      {stage0_57[126]},
      {stage1_57[56]}
   );
   gpc1_1 gpc1490 (
      {stage0_57[127]},
      {stage1_57[57]}
   );
   gpc1_1 gpc1491 (
      {stage0_58[117]},
      {stage1_58[49]}
   );
   gpc1_1 gpc1492 (
      {stage0_58[118]},
      {stage1_58[50]}
   );
   gpc1_1 gpc1493 (
      {stage0_58[119]},
      {stage1_58[51]}
   );
   gpc1_1 gpc1494 (
      {stage0_58[120]},
      {stage1_58[52]}
   );
   gpc1_1 gpc1495 (
      {stage0_58[121]},
      {stage1_58[53]}
   );
   gpc1_1 gpc1496 (
      {stage0_58[122]},
      {stage1_58[54]}
   );
   gpc1_1 gpc1497 (
      {stage0_58[123]},
      {stage1_58[55]}
   );
   gpc1_1 gpc1498 (
      {stage0_58[124]},
      {stage1_58[56]}
   );
   gpc1_1 gpc1499 (
      {stage0_58[125]},
      {stage1_58[57]}
   );
   gpc1_1 gpc1500 (
      {stage0_58[126]},
      {stage1_58[58]}
   );
   gpc1_1 gpc1501 (
      {stage0_58[127]},
      {stage1_58[59]}
   );
   gpc1_1 gpc1502 (
      {stage0_59[118]},
      {stage1_59[46]}
   );
   gpc1_1 gpc1503 (
      {stage0_59[119]},
      {stage1_59[47]}
   );
   gpc1_1 gpc1504 (
      {stage0_59[120]},
      {stage1_59[48]}
   );
   gpc1_1 gpc1505 (
      {stage0_59[121]},
      {stage1_59[49]}
   );
   gpc1_1 gpc1506 (
      {stage0_59[122]},
      {stage1_59[50]}
   );
   gpc1_1 gpc1507 (
      {stage0_59[123]},
      {stage1_59[51]}
   );
   gpc1_1 gpc1508 (
      {stage0_59[124]},
      {stage1_59[52]}
   );
   gpc1_1 gpc1509 (
      {stage0_59[125]},
      {stage1_59[53]}
   );
   gpc1_1 gpc1510 (
      {stage0_59[126]},
      {stage1_59[54]}
   );
   gpc1_1 gpc1511 (
      {stage0_59[127]},
      {stage1_59[55]}
   );
   gpc1_1 gpc1512 (
      {stage0_60[126]},
      {stage1_60[51]}
   );
   gpc1_1 gpc1513 (
      {stage0_60[127]},
      {stage1_60[52]}
   );
   gpc1_1 gpc1514 (
      {stage0_61[126]},
      {stage1_61[57]}
   );
   gpc1_1 gpc1515 (
      {stage0_61[127]},
      {stage1_61[58]}
   );
   gpc1_1 gpc1516 (
      {stage0_62[72]},
      {stage1_62[42]}
   );
   gpc1_1 gpc1517 (
      {stage0_62[73]},
      {stage1_62[43]}
   );
   gpc1_1 gpc1518 (
      {stage0_62[74]},
      {stage1_62[44]}
   );
   gpc1_1 gpc1519 (
      {stage0_62[75]},
      {stage1_62[45]}
   );
   gpc1_1 gpc1520 (
      {stage0_62[76]},
      {stage1_62[46]}
   );
   gpc1_1 gpc1521 (
      {stage0_62[77]},
      {stage1_62[47]}
   );
   gpc1_1 gpc1522 (
      {stage0_62[78]},
      {stage1_62[48]}
   );
   gpc1_1 gpc1523 (
      {stage0_62[79]},
      {stage1_62[49]}
   );
   gpc1_1 gpc1524 (
      {stage0_62[80]},
      {stage1_62[50]}
   );
   gpc1_1 gpc1525 (
      {stage0_62[81]},
      {stage1_62[51]}
   );
   gpc1_1 gpc1526 (
      {stage0_62[82]},
      {stage1_62[52]}
   );
   gpc1_1 gpc1527 (
      {stage0_62[83]},
      {stage1_62[53]}
   );
   gpc1_1 gpc1528 (
      {stage0_62[84]},
      {stage1_62[54]}
   );
   gpc1_1 gpc1529 (
      {stage0_62[85]},
      {stage1_62[55]}
   );
   gpc1_1 gpc1530 (
      {stage0_62[86]},
      {stage1_62[56]}
   );
   gpc1_1 gpc1531 (
      {stage0_62[87]},
      {stage1_62[57]}
   );
   gpc1_1 gpc1532 (
      {stage0_62[88]},
      {stage1_62[58]}
   );
   gpc1_1 gpc1533 (
      {stage0_62[89]},
      {stage1_62[59]}
   );
   gpc1_1 gpc1534 (
      {stage0_62[90]},
      {stage1_62[60]}
   );
   gpc1_1 gpc1535 (
      {stage0_62[91]},
      {stage1_62[61]}
   );
   gpc1_1 gpc1536 (
      {stage0_62[92]},
      {stage1_62[62]}
   );
   gpc1_1 gpc1537 (
      {stage0_62[93]},
      {stage1_62[63]}
   );
   gpc1_1 gpc1538 (
      {stage0_62[94]},
      {stage1_62[64]}
   );
   gpc1_1 gpc1539 (
      {stage0_62[95]},
      {stage1_62[65]}
   );
   gpc1_1 gpc1540 (
      {stage0_62[96]},
      {stage1_62[66]}
   );
   gpc1_1 gpc1541 (
      {stage0_62[97]},
      {stage1_62[67]}
   );
   gpc1_1 gpc1542 (
      {stage0_62[98]},
      {stage1_62[68]}
   );
   gpc1_1 gpc1543 (
      {stage0_62[99]},
      {stage1_62[69]}
   );
   gpc1_1 gpc1544 (
      {stage0_62[100]},
      {stage1_62[70]}
   );
   gpc1_1 gpc1545 (
      {stage0_62[101]},
      {stage1_62[71]}
   );
   gpc1_1 gpc1546 (
      {stage0_62[102]},
      {stage1_62[72]}
   );
   gpc1_1 gpc1547 (
      {stage0_62[103]},
      {stage1_62[73]}
   );
   gpc1_1 gpc1548 (
      {stage0_62[104]},
      {stage1_62[74]}
   );
   gpc1_1 gpc1549 (
      {stage0_62[105]},
      {stage1_62[75]}
   );
   gpc1_1 gpc1550 (
      {stage0_62[106]},
      {stage1_62[76]}
   );
   gpc1_1 gpc1551 (
      {stage0_62[107]},
      {stage1_62[77]}
   );
   gpc1_1 gpc1552 (
      {stage0_62[108]},
      {stage1_62[78]}
   );
   gpc1_1 gpc1553 (
      {stage0_62[109]},
      {stage1_62[79]}
   );
   gpc1_1 gpc1554 (
      {stage0_62[110]},
      {stage1_62[80]}
   );
   gpc1_1 gpc1555 (
      {stage0_62[111]},
      {stage1_62[81]}
   );
   gpc1_1 gpc1556 (
      {stage0_62[112]},
      {stage1_62[82]}
   );
   gpc1_1 gpc1557 (
      {stage0_62[113]},
      {stage1_62[83]}
   );
   gpc1_1 gpc1558 (
      {stage0_62[114]},
      {stage1_62[84]}
   );
   gpc1_1 gpc1559 (
      {stage0_62[115]},
      {stage1_62[85]}
   );
   gpc1_1 gpc1560 (
      {stage0_62[116]},
      {stage1_62[86]}
   );
   gpc1_1 gpc1561 (
      {stage0_62[117]},
      {stage1_62[87]}
   );
   gpc1_1 gpc1562 (
      {stage0_62[118]},
      {stage1_62[88]}
   );
   gpc1_1 gpc1563 (
      {stage0_62[119]},
      {stage1_62[89]}
   );
   gpc1_1 gpc1564 (
      {stage0_62[120]},
      {stage1_62[90]}
   );
   gpc1_1 gpc1565 (
      {stage0_62[121]},
      {stage1_62[91]}
   );
   gpc1_1 gpc1566 (
      {stage0_62[122]},
      {stage1_62[92]}
   );
   gpc1_1 gpc1567 (
      {stage0_62[123]},
      {stage1_62[93]}
   );
   gpc1_1 gpc1568 (
      {stage0_62[124]},
      {stage1_62[94]}
   );
   gpc1_1 gpc1569 (
      {stage0_62[125]},
      {stage1_62[95]}
   );
   gpc1_1 gpc1570 (
      {stage0_62[126]},
      {stage1_62[96]}
   );
   gpc1_1 gpc1571 (
      {stage0_62[127]},
      {stage1_62[97]}
   );
   gpc1_1 gpc1572 (
      {stage0_63[108]},
      {stage1_63[33]}
   );
   gpc1_1 gpc1573 (
      {stage0_63[109]},
      {stage1_63[34]}
   );
   gpc1_1 gpc1574 (
      {stage0_63[110]},
      {stage1_63[35]}
   );
   gpc1_1 gpc1575 (
      {stage0_63[111]},
      {stage1_63[36]}
   );
   gpc1_1 gpc1576 (
      {stage0_63[112]},
      {stage1_63[37]}
   );
   gpc1_1 gpc1577 (
      {stage0_63[113]},
      {stage1_63[38]}
   );
   gpc1_1 gpc1578 (
      {stage0_63[114]},
      {stage1_63[39]}
   );
   gpc1_1 gpc1579 (
      {stage0_63[115]},
      {stage1_63[40]}
   );
   gpc1_1 gpc1580 (
      {stage0_63[116]},
      {stage1_63[41]}
   );
   gpc1_1 gpc1581 (
      {stage0_63[117]},
      {stage1_63[42]}
   );
   gpc1_1 gpc1582 (
      {stage0_63[118]},
      {stage1_63[43]}
   );
   gpc1_1 gpc1583 (
      {stage0_63[119]},
      {stage1_63[44]}
   );
   gpc1_1 gpc1584 (
      {stage0_63[120]},
      {stage1_63[45]}
   );
   gpc1_1 gpc1585 (
      {stage0_63[121]},
      {stage1_63[46]}
   );
   gpc1_1 gpc1586 (
      {stage0_63[122]},
      {stage1_63[47]}
   );
   gpc1_1 gpc1587 (
      {stage0_63[123]},
      {stage1_63[48]}
   );
   gpc1_1 gpc1588 (
      {stage0_63[124]},
      {stage1_63[49]}
   );
   gpc1_1 gpc1589 (
      {stage0_63[125]},
      {stage1_63[50]}
   );
   gpc1_1 gpc1590 (
      {stage0_63[126]},
      {stage1_63[51]}
   );
   gpc1_1 gpc1591 (
      {stage0_63[127]},
      {stage1_63[52]}
   );
   gpc1163_5 gpc1592 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc1593 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[6]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc1594 (
      {stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[7]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc1595 (
      {stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc1596 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc606_5 gpc1597 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18]},
      {stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc1598 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc1599 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc1600 (
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[5],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc1163_5 gpc1601 (
      {stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_5[0]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[3],stage2_5[6],stage2_4[9],stage2_3[9]}
   );
   gpc606_5 gpc1602 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[1],stage2_6[4],stage2_5[7],stage2_4[10],stage2_3[10]}
   );
   gpc606_5 gpc1603 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[2],stage2_6[5],stage2_5[8],stage2_4[11],stage2_3[11]}
   );
   gpc606_5 gpc1604 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[3],stage2_6[6],stage2_5[9],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc1605 (
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44]},
      {stage1_4[24]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[4],stage2_6[7],stage2_5[10],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc1606 (
      {stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage1_4[25]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[5],stage2_6[8],stage2_5[11],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc1607 (
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54]},
      {stage1_4[26]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[6],stage2_6[9],stage2_5[12],stage2_4[15],stage2_3[15]}
   );
   gpc606_5 gpc1608 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[0],stage2_7[7],stage2_6[10],stage2_5[13],stage2_4[16]}
   );
   gpc615_5 gpc1609 (
      {stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36], stage1_4[37]},
      {stage1_5[37]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[1],stage2_7[8],stage2_6[11],stage2_5[14],stage2_4[17]}
   );
   gpc615_5 gpc1610 (
      {stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42]},
      {stage1_5[38]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[2],stage2_7[9],stage2_6[12],stage2_5[15],stage2_4[18]}
   );
   gpc615_5 gpc1611 (
      {stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_5[39]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[3],stage2_7[10],stage2_6[13],stage2_5[16],stage2_4[19]}
   );
   gpc615_5 gpc1612 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52]},
      {stage1_5[40]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[4],stage2_7[11],stage2_6[14],stage2_5[17],stage2_4[20]}
   );
   gpc615_5 gpc1613 (
      {stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_5[41]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[5],stage2_7[12],stage2_6[15],stage2_5[18],stage2_4[21]}
   );
   gpc615_5 gpc1614 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_5[42]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[6],stage2_7[13],stage2_6[16],stage2_5[19],stage2_4[22]}
   );
   gpc606_5 gpc1615 (
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[7],stage2_7[14],stage2_6[17]}
   );
   gpc606_5 gpc1616 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[8],stage2_7[15],stage2_6[18]}
   );
   gpc615_5 gpc1617 (
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage1_7[0]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[9],stage2_7[16],stage2_6[19]}
   );
   gpc615_5 gpc1618 (
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64]},
      {stage1_7[1]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[3],stage2_8[10],stage2_7[17],stage2_6[20]}
   );
   gpc615_5 gpc1619 (
      {stage1_6[65], stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69]},
      {stage1_7[2]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[4],stage2_8[11],stage2_7[18],stage2_6[21]}
   );
   gpc615_5 gpc1620 (
      {stage1_6[70], stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74]},
      {stage1_7[3]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[5],stage2_8[12],stage2_7[19],stage2_6[22]}
   );
   gpc615_5 gpc1621 (
      {stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79]},
      {stage1_7[4]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[6],stage2_8[13],stage2_7[20],stage2_6[23]}
   );
   gpc615_5 gpc1622 (
      {stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage1_7[5]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[7],stage2_8[14],stage2_7[21],stage2_6[24]}
   );
   gpc615_5 gpc1623 (
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], 1'b0},
      {stage1_7[6]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[8],stage2_8[15],stage2_7[22],stage2_6[25]}
   );
   gpc1406_5 gpc1624 (
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[9],stage2_9[9],stage2_8[16],stage2_7[23]}
   );
   gpc117_4 gpc1625 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage1_8[54]},
      {stage1_9[4]},
      {stage2_10[10],stage2_9[10],stage2_8[17],stage2_7[24]}
   );
   gpc117_4 gpc1626 (
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26]},
      {stage1_8[55]},
      {stage1_9[5]},
      {stage2_10[11],stage2_9[11],stage2_8[18],stage2_7[25]}
   );
   gpc117_4 gpc1627 (
      {stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[56]},
      {stage1_9[6]},
      {stage2_10[12],stage2_9[12],stage2_8[19],stage2_7[26]}
   );
   gpc117_4 gpc1628 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40]},
      {stage1_8[57]},
      {stage1_9[7]},
      {stage2_10[13],stage2_9[13],stage2_8[20],stage2_7[27]}
   );
   gpc606_5 gpc1629 (
      {stage1_7[41], stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13]},
      {stage2_11[1],stage2_10[14],stage2_9[14],stage2_8[21],stage2_7[28]}
   );
   gpc606_5 gpc1630 (
      {stage1_7[47], stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52]},
      {stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage2_11[2],stage2_10[15],stage2_9[15],stage2_8[22],stage2_7[29]}
   );
   gpc606_5 gpc1631 (
      {stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24], stage1_9[25]},
      {stage2_11[3],stage2_10[16],stage2_9[16],stage2_8[23],stage2_7[30]}
   );
   gpc615_5 gpc1632 (
      {stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63]},
      {stage1_8[58]},
      {stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30], stage1_9[31]},
      {stage2_11[4],stage2_10[17],stage2_9[17],stage2_8[24],stage2_7[31]}
   );
   gpc606_5 gpc1633 (
      {stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35], stage1_9[36], stage1_9[37]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[5],stage2_10[18],stage2_9[18]}
   );
   gpc615_5 gpc1634 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[6],stage2_10[19]}
   );
   gpc615_5 gpc1635 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10]},
      {stage1_11[7]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[7],stage2_10[20]}
   );
   gpc615_5 gpc1636 (
      {stage1_10[11], stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[8]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[8],stage2_10[21]}
   );
   gpc615_5 gpc1637 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20]},
      {stage1_11[9]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[9],stage2_10[22]}
   );
   gpc615_5 gpc1638 (
      {stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_11[10]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[10],stage2_10[23]}
   );
   gpc615_5 gpc1639 (
      {stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_11[11]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[11],stage2_10[24]}
   );
   gpc615_5 gpc1640 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_11[12]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[12],stage2_10[25]}
   );
   gpc606_5 gpc1641 (
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[8],stage2_12[8],stage2_11[13]}
   );
   gpc606_5 gpc1642 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[9],stage2_12[9],stage2_11[14]}
   );
   gpc606_5 gpc1643 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[10],stage2_12[10],stage2_11[15]}
   );
   gpc606_5 gpc1644 (
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[11],stage2_12[11],stage2_11[16]}
   );
   gpc606_5 gpc1645 (
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[12],stage2_12[12],stage2_11[17]}
   );
   gpc606_5 gpc1646 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[12],stage2_13[13],stage2_12[13],stage2_11[18]}
   );
   gpc615_5 gpc1647 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[42]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[13],stage2_13[14],stage2_12[14],stage2_11[19]}
   );
   gpc615_5 gpc1648 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[43]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[14],stage2_13[15],stage2_12[15],stage2_11[20]}
   );
   gpc615_5 gpc1649 (
      {stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63]},
      {stage1_12[44]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[15],stage2_13[16],stage2_12[16],stage2_11[21]}
   );
   gpc606_5 gpc1650 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[0],stage2_16[0],stage2_15[9],stage2_14[16]}
   );
   gpc606_5 gpc1651 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[1],stage2_16[1],stage2_15[10],stage2_14[17]}
   );
   gpc606_5 gpc1652 (
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[2],stage2_16[2],stage2_15[11],stage2_14[18]}
   );
   gpc615_5 gpc1653 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22]},
      {stage1_15[0]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[3],stage2_16[3],stage2_15[12],stage2_14[19]}
   );
   gpc615_5 gpc1654 (
      {stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27]},
      {stage1_15[1]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[4],stage2_16[4],stage2_15[13],stage2_14[20]}
   );
   gpc615_5 gpc1655 (
      {stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31], stage1_14[32]},
      {stage1_15[2]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[5],stage2_16[5],stage2_15[14],stage2_14[21]}
   );
   gpc615_5 gpc1656 (
      {stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_15[3]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[6],stage2_16[6],stage2_15[15],stage2_14[22]}
   );
   gpc615_5 gpc1657 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_15[4]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[7],stage2_16[7],stage2_15[16],stage2_14[23]}
   );
   gpc615_5 gpc1658 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_15[5]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[8],stage2_16[8],stage2_15[17],stage2_14[24]}
   );
   gpc615_5 gpc1659 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52]},
      {stage1_15[6]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[9],stage2_16[9],stage2_15[18],stage2_14[25]}
   );
   gpc1415_5 gpc1660 (
      {stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[60]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[10],stage2_17[10],stage2_16[10],stage2_15[19]}
   );
   gpc2116_5 gpc1661 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[61]},
      {stage1_17[4]},
      {stage1_18[1], stage1_18[2]},
      {stage2_19[1],stage2_18[11],stage2_17[11],stage2_16[11],stage2_15[20]}
   );
   gpc2116_5 gpc1662 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[62]},
      {stage1_17[5]},
      {stage1_18[3], stage1_18[4]},
      {stage2_19[2],stage2_18[12],stage2_17[12],stage2_16[12],stage2_15[21]}
   );
   gpc2116_5 gpc1663 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[63]},
      {stage1_17[6]},
      {stage1_18[5], stage1_18[6]},
      {stage2_19[3],stage2_18[13],stage2_17[13],stage2_16[13],stage2_15[22]}
   );
   gpc2116_5 gpc1664 (
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[64]},
      {stage1_17[7]},
      {stage1_18[7], stage1_18[8]},
      {stage2_19[4],stage2_18[14],stage2_17[14],stage2_16[14],stage2_15[23]}
   );
   gpc2116_5 gpc1665 (
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage1_16[65]},
      {stage1_17[8]},
      {stage1_18[9], stage1_18[10]},
      {stage2_19[5],stage2_18[15],stage2_17[15],stage2_16[15],stage2_15[24]}
   );
   gpc615_5 gpc1666 (
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46]},
      {stage1_16[66]},
      {stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12], stage1_17[13], stage1_17[14]},
      {stage2_19[6],stage2_18[16],stage2_17[16],stage2_16[16],stage2_15[25]}
   );
   gpc615_5 gpc1667 (
      {stage1_15[47], stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51]},
      {stage1_16[67]},
      {stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18], stage1_17[19], stage1_17[20]},
      {stage2_19[7],stage2_18[17],stage2_17[17],stage2_16[17],stage2_15[26]}
   );
   gpc615_5 gpc1668 (
      {stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55], stage1_15[56]},
      {stage1_16[68]},
      {stage1_17[21], stage1_17[22], stage1_17[23], stage1_17[24], stage1_17[25], stage1_17[26]},
      {stage2_19[8],stage2_18[18],stage2_17[18],stage2_16[18],stage2_15[27]}
   );
   gpc615_5 gpc1669 (
      {stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage1_16[69]},
      {stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30], stage1_17[31], stage1_17[32]},
      {stage2_19[9],stage2_18[19],stage2_17[19],stage2_16[19],stage2_15[28]}
   );
   gpc615_5 gpc1670 (
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66]},
      {stage1_16[70]},
      {stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36], stage1_17[37], stage1_17[38]},
      {stage2_19[10],stage2_18[20],stage2_17[20],stage2_16[20],stage2_15[29]}
   );
   gpc606_5 gpc1671 (
      {stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76]},
      {stage1_18[11], stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16]},
      {stage2_20[0],stage2_19[11],stage2_18[21],stage2_17[21],stage2_16[21]}
   );
   gpc606_5 gpc1672 (
      {stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82]},
      {stage1_18[17], stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage2_20[1],stage2_19[12],stage2_18[22],stage2_17[22],stage2_16[22]}
   );
   gpc606_5 gpc1673 (
      {stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88]},
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28]},
      {stage2_20[2],stage2_19[13],stage2_18[23],stage2_17[23],stage2_16[23]}
   );
   gpc135_4 gpc1674 (
      {stage1_17[39], stage1_17[40], stage1_17[41], stage1_17[42], stage1_17[43]},
      {stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage1_19[0]},
      {stage2_20[3],stage2_19[14],stage2_18[24],stage2_17[24]}
   );
   gpc1343_5 gpc1675 (
      {stage1_17[44], stage1_17[45], stage1_17[46]},
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage1_19[1], stage1_19[2], stage1_19[3]},
      {stage1_20[0]},
      {stage2_21[0],stage2_20[4],stage2_19[15],stage2_18[25],stage2_17[25]}
   );
   gpc1343_5 gpc1676 (
      {stage1_17[47], stage1_17[48], stage1_17[49]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39]},
      {stage1_19[4], stage1_19[5], stage1_19[6]},
      {stage1_20[1]},
      {stage2_21[1],stage2_20[5],stage2_19[16],stage2_18[26],stage2_17[26]}
   );
   gpc606_5 gpc1677 (
      {stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53], stage1_17[54], stage1_17[55]},
      {stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11], stage1_19[12]},
      {stage2_21[2],stage2_20[6],stage2_19[17],stage2_18[27],stage2_17[27]}
   );
   gpc606_5 gpc1678 (
      {stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59], stage1_17[60], stage1_17[61]},
      {stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17], stage1_19[18]},
      {stage2_21[3],stage2_20[7],stage2_19[18],stage2_18[28],stage2_17[28]}
   );
   gpc615_5 gpc1679 (
      {stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage1_20[2]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[4],stage2_20[8],stage2_19[19]}
   );
   gpc615_5 gpc1680 (
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28]},
      {stage1_20[3]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[5],stage2_20[9],stage2_19[20]}
   );
   gpc615_5 gpc1681 (
      {stage1_19[29], stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33]},
      {stage1_20[4]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[6],stage2_20[10],stage2_19[21]}
   );
   gpc615_5 gpc1682 (
      {stage1_19[34], stage1_19[35], stage1_19[36], stage1_19[37], stage1_19[38]},
      {stage1_20[5]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[7],stage2_20[11],stage2_19[22]}
   );
   gpc615_5 gpc1683 (
      {stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42], stage1_19[43]},
      {stage1_20[6]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[8],stage2_20[12],stage2_19[23]}
   );
   gpc615_5 gpc1684 (
      {stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47], stage1_19[48]},
      {stage1_20[7]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[9],stage2_20[13],stage2_19[24]}
   );
   gpc615_5 gpc1685 (
      {stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage1_20[8]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[6],stage2_21[10],stage2_20[14],stage2_19[25]}
   );
   gpc606_5 gpc1686 (
      {stage1_20[9], stage1_20[10], stage1_20[11], stage1_20[12], stage1_20[13], stage1_20[14]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[7],stage2_22[7],stage2_21[11],stage2_20[15]}
   );
   gpc606_5 gpc1687 (
      {stage1_20[15], stage1_20[16], stage1_20[17], stage1_20[18], stage1_20[19], stage1_20[20]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[8],stage2_22[8],stage2_21[12],stage2_20[16]}
   );
   gpc606_5 gpc1688 (
      {stage1_20[21], stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[9],stage2_22[9],stage2_21[13],stage2_20[17]}
   );
   gpc606_5 gpc1689 (
      {stage1_20[27], stage1_20[28], stage1_20[29], stage1_20[30], stage1_20[31], stage1_20[32]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[10],stage2_22[10],stage2_21[14],stage2_20[18]}
   );
   gpc606_5 gpc1690 (
      {stage1_20[33], stage1_20[34], stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[11],stage2_22[11],stage2_21[15],stage2_20[19]}
   );
   gpc606_5 gpc1691 (
      {stage1_20[39], stage1_20[40], stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[12],stage2_22[12],stage2_21[16],stage2_20[20]}
   );
   gpc606_5 gpc1692 (
      {stage1_20[45], stage1_20[46], stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[13],stage2_22[13],stage2_21[17],stage2_20[21]}
   );
   gpc606_5 gpc1693 (
      {stage1_20[51], stage1_20[52], stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[14],stage2_22[14],stage2_21[18],stage2_20[22]}
   );
   gpc615_5 gpc1694 (
      {stage1_20[57], stage1_20[58], stage1_20[59], stage1_20[60], stage1_20[61]},
      {stage1_21[42]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[15],stage2_22[15],stage2_21[19],stage2_20[23]}
   );
   gpc606_5 gpc1695 (
      {stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[9],stage2_23[16],stage2_22[16],stage2_21[20]}
   );
   gpc606_5 gpc1696 (
      {stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[10],stage2_23[17],stage2_22[17],stage2_21[21]}
   );
   gpc615_5 gpc1697 (
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[0],stage2_25[2],stage2_24[11],stage2_23[18]}
   );
   gpc615_5 gpc1698 (
      {stage1_23[17], stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21]},
      {stage1_24[1]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[1],stage2_25[3],stage2_24[12],stage2_23[19]}
   );
   gpc615_5 gpc1699 (
      {stage1_23[22], stage1_23[23], stage1_23[24], stage1_23[25], stage1_23[26]},
      {stage1_24[2]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[2],stage2_25[4],stage2_24[13],stage2_23[20]}
   );
   gpc615_5 gpc1700 (
      {stage1_23[27], stage1_23[28], stage1_23[29], stage1_23[30], stage1_23[31]},
      {stage1_24[3]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[3],stage2_25[5],stage2_24[14],stage2_23[21]}
   );
   gpc615_5 gpc1701 (
      {stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36]},
      {stage1_24[4]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[4],stage2_25[6],stage2_24[15],stage2_23[22]}
   );
   gpc615_5 gpc1702 (
      {stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage1_24[5]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[5],stage2_25[7],stage2_24[16],stage2_23[23]}
   );
   gpc615_5 gpc1703 (
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46]},
      {stage1_24[6]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[6],stage2_25[8],stage2_24[17],stage2_23[24]}
   );
   gpc615_5 gpc1704 (
      {stage1_23[47], stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51]},
      {stage1_24[7]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[7],stage2_25[9],stage2_24[18],stage2_23[25]}
   );
   gpc606_5 gpc1705 (
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[8],stage2_25[10],stage2_24[19]}
   );
   gpc606_5 gpc1706 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[9],stage2_25[11],stage2_24[20]}
   );
   gpc606_5 gpc1707 (
      {stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[10],stage2_25[12],stage2_24[21]}
   );
   gpc606_5 gpc1708 (
      {stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30], stage1_24[31]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[11],stage2_25[13],stage2_24[22]}
   );
   gpc606_5 gpc1709 (
      {stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36], stage1_24[37]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[12],stage2_26[12],stage2_25[14],stage2_24[23]}
   );
   gpc606_5 gpc1710 (
      {stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42], stage1_24[43]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[13],stage2_26[13],stage2_25[15],stage2_24[24]}
   );
   gpc606_5 gpc1711 (
      {stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48], stage1_24[49]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[14],stage2_26[14],stage2_25[16],stage2_24[25]}
   );
   gpc606_5 gpc1712 (
      {stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54], stage1_24[55]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[15],stage2_26[15],stage2_25[17],stage2_24[26]}
   );
   gpc606_5 gpc1713 (
      {stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59], stage1_24[60], stage1_24[61]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[16],stage2_26[16],stage2_25[18],stage2_24[27]}
   );
   gpc615_5 gpc1714 (
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58]},
      {stage1_27[0]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[0],stage2_28[9],stage2_27[17],stage2_26[17]}
   );
   gpc615_5 gpc1715 (
      {stage1_26[59], stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63]},
      {stage1_27[1]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[1],stage2_28[10],stage2_27[18],stage2_26[18]}
   );
   gpc615_5 gpc1716 (
      {stage1_26[64], stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68]},
      {stage1_27[2]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[2],stage2_28[11],stage2_27[19],stage2_26[19]}
   );
   gpc615_5 gpc1717 (
      {stage1_26[69], stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73]},
      {stage1_27[3]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[3],stage2_28[12],stage2_27[20],stage2_26[20]}
   );
   gpc615_5 gpc1718 (
      {stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77], stage1_26[78]},
      {stage1_27[4]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[4],stage2_28[13],stage2_27[21],stage2_26[21]}
   );
   gpc615_5 gpc1719 (
      {stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage1_28[30]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[5],stage2_29[5],stage2_28[14],stage2_27[22]}
   );
   gpc615_5 gpc1720 (
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14]},
      {stage1_28[31]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[6],stage2_29[6],stage2_28[15],stage2_27[23]}
   );
   gpc615_5 gpc1721 (
      {stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19]},
      {stage1_28[32]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[7],stage2_29[7],stage2_28[16],stage2_27[24]}
   );
   gpc615_5 gpc1722 (
      {stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23], stage1_27[24]},
      {stage1_28[33]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[8],stage2_29[8],stage2_28[17],stage2_27[25]}
   );
   gpc615_5 gpc1723 (
      {stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage1_28[34]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[9],stage2_29[9],stage2_28[18],stage2_27[26]}
   );
   gpc615_5 gpc1724 (
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34]},
      {stage1_28[35]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[10],stage2_29[10],stage2_28[19],stage2_27[27]}
   );
   gpc615_5 gpc1725 (
      {stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39]},
      {stage1_28[36]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[11],stage2_29[11],stage2_28[20],stage2_27[28]}
   );
   gpc615_5 gpc1726 (
      {stage1_27[40], stage1_27[41], stage1_27[42], stage1_27[43], stage1_27[44]},
      {stage1_28[37]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[12],stage2_29[12],stage2_28[21],stage2_27[29]}
   );
   gpc615_5 gpc1727 (
      {stage1_27[45], stage1_27[46], stage1_27[47], stage1_27[48], stage1_27[49]},
      {stage1_28[38]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[13],stage2_29[13],stage2_28[22],stage2_27[30]}
   );
   gpc615_5 gpc1728 (
      {stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53], stage1_27[54]},
      {stage1_28[39]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[14],stage2_29[14],stage2_28[23],stage2_27[31]}
   );
   gpc606_5 gpc1729 (
      {stage1_28[40], stage1_28[41], stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[10],stage2_30[15],stage2_29[15],stage2_28[24]}
   );
   gpc606_5 gpc1730 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[11],stage2_30[16],stage2_29[16]}
   );
   gpc606_5 gpc1731 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[12],stage2_30[17],stage2_29[17]}
   );
   gpc606_5 gpc1732 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[3],stage2_31[13],stage2_30[18],stage2_29[18]}
   );
   gpc1406_5 gpc1733 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3]},
      {stage1_33[0]},
      {stage2_34[0],stage2_33[3],stage2_32[4],stage2_31[14],stage2_30[19]}
   );
   gpc615_5 gpc1734 (
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16]},
      {stage1_31[18]},
      {stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9]},
      {stage2_34[1],stage2_33[4],stage2_32[5],stage2_31[15],stage2_30[20]}
   );
   gpc615_5 gpc1735 (
      {stage1_30[17], stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21]},
      {stage1_31[19]},
      {stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15]},
      {stage2_34[2],stage2_33[5],stage2_32[6],stage2_31[16],stage2_30[21]}
   );
   gpc615_5 gpc1736 (
      {stage1_30[22], stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26]},
      {stage1_31[20]},
      {stage1_32[16], stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21]},
      {stage2_34[3],stage2_33[6],stage2_32[7],stage2_31[17],stage2_30[22]}
   );
   gpc615_5 gpc1737 (
      {stage1_30[27], stage1_30[28], stage1_30[29], stage1_30[30], stage1_30[31]},
      {stage1_31[21]},
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage2_34[4],stage2_33[7],stage2_32[8],stage2_31[18],stage2_30[23]}
   );
   gpc615_5 gpc1738 (
      {stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35], stage1_30[36]},
      {stage1_31[22]},
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage2_34[5],stage2_33[8],stage2_32[9],stage2_31[19],stage2_30[24]}
   );
   gpc615_5 gpc1739 (
      {stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage1_31[23]},
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage2_34[6],stage2_33[9],stage2_32[10],stage2_31[20],stage2_30[25]}
   );
   gpc615_5 gpc1740 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46]},
      {stage1_31[24]},
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage2_34[7],stage2_33[10],stage2_32[11],stage2_31[21],stage2_30[26]}
   );
   gpc606_5 gpc1741 (
      {stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29], stage1_31[30]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[0],stage2_34[8],stage2_33[11],stage2_32[12],stage2_31[22]}
   );
   gpc606_5 gpc1742 (
      {stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35], stage1_31[36]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[1],stage2_34[9],stage2_33[12],stage2_32[13],stage2_31[23]}
   );
   gpc606_5 gpc1743 (
      {stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42]},
      {stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18]},
      {stage2_35[2],stage2_34[10],stage2_33[13],stage2_32[14],stage2_31[24]}
   );
   gpc606_5 gpc1744 (
      {stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48]},
      {stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24]},
      {stage2_35[3],stage2_34[11],stage2_33[14],stage2_32[15],stage2_31[25]}
   );
   gpc606_5 gpc1745 (
      {stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54]},
      {stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30]},
      {stage2_35[4],stage2_34[12],stage2_33[15],stage2_32[16],stage2_31[26]}
   );
   gpc606_5 gpc1746 (
      {stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59], 1'b0},
      {stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36]},
      {stage2_35[5],stage2_34[13],stage2_33[16],stage2_32[17],stage2_31[27]}
   );
   gpc606_5 gpc1747 (
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[6],stage2_34[14],stage2_33[17],stage2_32[18]}
   );
   gpc606_5 gpc1748 (
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[7],stage2_34[15],stage2_33[18],stage2_32[19]}
   );
   gpc606_5 gpc1749 (
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[8],stage2_34[16],stage2_33[19],stage2_32[20]}
   );
   gpc606_5 gpc1750 (
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[9],stage2_34[17],stage2_33[20],stage2_32[21]}
   );
   gpc606_5 gpc1751 (
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[10],stage2_34[18],stage2_33[21],stage2_32[22]}
   );
   gpc606_5 gpc1752 (
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[11],stage2_34[19],stage2_33[22],stage2_32[23]}
   );
   gpc606_5 gpc1753 (
      {stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[6],stage2_35[12],stage2_34[20],stage2_33[23]}
   );
   gpc606_5 gpc1754 (
      {stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[7],stage2_35[13],stage2_34[21],stage2_33[24]}
   );
   gpc606_5 gpc1755 (
      {stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[8],stage2_35[14],stage2_34[22],stage2_33[25]}
   );
   gpc606_5 gpc1756 (
      {stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[9],stage2_35[15],stage2_34[23],stage2_33[26]}
   );
   gpc615_5 gpc1757 (
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40]},
      {stage1_35[24]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[4],stage2_36[10],stage2_35[16],stage2_34[24]}
   );
   gpc615_5 gpc1758 (
      {stage1_34[41], stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45]},
      {stage1_35[25]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[5],stage2_36[11],stage2_35[17],stage2_34[25]}
   );
   gpc615_5 gpc1759 (
      {stage1_34[46], stage1_34[47], stage1_34[48], stage1_34[49], stage1_34[50]},
      {stage1_35[26]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[6],stage2_36[12],stage2_35[18],stage2_34[26]}
   );
   gpc615_5 gpc1760 (
      {stage1_34[51], stage1_34[52], stage1_34[53], stage1_34[54], stage1_34[55]},
      {stage1_35[27]},
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23]},
      {stage2_38[3],stage2_37[7],stage2_36[13],stage2_35[19],stage2_34[27]}
   );
   gpc615_5 gpc1761 (
      {stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59], stage1_34[60]},
      {stage1_35[28]},
      {stage1_36[24], stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29]},
      {stage2_38[4],stage2_37[8],stage2_36[14],stage2_35[20],stage2_34[28]}
   );
   gpc615_5 gpc1762 (
      {stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage1_35[29]},
      {stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35]},
      {stage2_38[5],stage2_37[9],stage2_36[15],stage2_35[21],stage2_34[29]}
   );
   gpc606_5 gpc1763 (
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[6],stage2_37[10],stage2_36[16],stage2_35[22]}
   );
   gpc606_5 gpc1764 (
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[7],stage2_37[11],stage2_36[17],stage2_35[23]}
   );
   gpc606_5 gpc1765 (
      {stage1_36[36], stage1_36[37], stage1_36[38], stage1_36[39], stage1_36[40], stage1_36[41]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[2],stage2_38[8],stage2_37[12],stage2_36[18]}
   );
   gpc606_5 gpc1766 (
      {stage1_36[42], stage1_36[43], stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47]},
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11]},
      {stage2_40[1],stage2_39[3],stage2_38[9],stage2_37[13],stage2_36[19]}
   );
   gpc606_5 gpc1767 (
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[2],stage2_39[4],stage2_38[10],stage2_37[14]}
   );
   gpc606_5 gpc1768 (
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[3],stage2_39[5],stage2_38[11],stage2_37[15]}
   );
   gpc615_5 gpc1769 (
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28]},
      {stage1_38[12]},
      {stage1_39[12], stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17]},
      {stage2_41[2],stage2_40[4],stage2_39[6],stage2_38[12],stage2_37[16]}
   );
   gpc615_5 gpc1770 (
      {stage1_37[29], stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33]},
      {stage1_38[13]},
      {stage1_39[18], stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23]},
      {stage2_41[3],stage2_40[5],stage2_39[7],stage2_38[13],stage2_37[17]}
   );
   gpc615_5 gpc1771 (
      {stage1_37[34], stage1_37[35], stage1_37[36], stage1_37[37], stage1_37[38]},
      {stage1_38[14]},
      {stage1_39[24], stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29]},
      {stage2_41[4],stage2_40[6],stage2_39[8],stage2_38[14],stage2_37[18]}
   );
   gpc615_5 gpc1772 (
      {stage1_37[39], stage1_37[40], stage1_37[41], stage1_37[42], stage1_37[43]},
      {stage1_38[15]},
      {stage1_39[30], stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35]},
      {stage2_41[5],stage2_40[7],stage2_39[9],stage2_38[15],stage2_37[19]}
   );
   gpc615_5 gpc1773 (
      {stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47], stage1_37[48]},
      {stage1_38[16]},
      {stage1_39[36], stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41]},
      {stage2_41[6],stage2_40[8],stage2_39[10],stage2_38[16],stage2_37[20]}
   );
   gpc615_5 gpc1774 (
      {stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage1_38[17]},
      {stage1_39[42], stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47]},
      {stage2_41[7],stage2_40[9],stage2_39[11],stage2_38[17],stage2_37[21]}
   );
   gpc615_5 gpc1775 (
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58]},
      {stage1_38[18]},
      {stage1_39[48], stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53]},
      {stage2_41[8],stage2_40[10],stage2_39[12],stage2_38[18],stage2_37[22]}
   );
   gpc615_5 gpc1776 (
      {stage1_37[59], stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63]},
      {stage1_38[19]},
      {stage1_39[54], stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59]},
      {stage2_41[9],stage2_40[11],stage2_39[13],stage2_38[19],stage2_37[23]}
   );
   gpc615_5 gpc1777 (
      {stage1_37[64], stage1_37[65], stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_38[20]},
      {stage1_39[60], stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65]},
      {stage2_41[10],stage2_40[12],stage2_39[14],stage2_38[20],stage2_37[24]}
   );
   gpc615_5 gpc1778 (
      {stage1_37[69], stage1_37[70], stage1_37[71], stage1_37[72], stage1_37[73]},
      {stage1_38[21]},
      {stage1_39[66], stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71]},
      {stage2_41[11],stage2_40[13],stage2_39[15],stage2_38[21],stage2_37[25]}
   );
   gpc615_5 gpc1779 (
      {stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77], stage1_37[78]},
      {stage1_38[22]},
      {stage1_39[72], stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77]},
      {stage2_41[12],stage2_40[14],stage2_39[16],stage2_38[22],stage2_37[26]}
   );
   gpc615_5 gpc1780 (
      {stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage1_38[23]},
      {stage1_39[78], stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83]},
      {stage2_41[13],stage2_40[15],stage2_39[17],stage2_38[23],stage2_37[27]}
   );
   gpc615_5 gpc1781 (
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88]},
      {stage1_38[24]},
      {stage1_39[84], stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89]},
      {stage2_41[14],stage2_40[16],stage2_39[18],stage2_38[24],stage2_37[28]}
   );
   gpc615_5 gpc1782 (
      {stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28], stage1_38[29]},
      {stage1_39[90]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[15],stage2_40[17],stage2_39[19],stage2_38[25]}
   );
   gpc615_5 gpc1783 (
      {stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34]},
      {stage1_39[91]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[16],stage2_40[18],stage2_39[20],stage2_38[26]}
   );
   gpc606_5 gpc1784 (
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[2],stage2_41[17],stage2_40[19]}
   );
   gpc606_5 gpc1785 (
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[3],stage2_41[18],stage2_40[20]}
   );
   gpc606_5 gpc1786 (
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[4],stage2_41[19],stage2_40[21]}
   );
   gpc606_5 gpc1787 (
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[5],stage2_41[20],stage2_40[22]}
   );
   gpc606_5 gpc1788 (
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[6],stage2_41[21],stage2_40[23]}
   );
   gpc606_5 gpc1789 (
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[7],stage2_41[22],stage2_40[24]}
   );
   gpc606_5 gpc1790 (
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[8],stage2_41[23],stage2_40[25]}
   );
   gpc615_5 gpc1791 (
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4]},
      {stage1_42[42]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[7],stage2_43[7],stage2_42[9],stage2_41[24]}
   );
   gpc615_5 gpc1792 (
      {stage1_41[5], stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9]},
      {stage1_42[43]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[8],stage2_43[8],stage2_42[10],stage2_41[25]}
   );
   gpc615_5 gpc1793 (
      {stage1_41[10], stage1_41[11], stage1_41[12], stage1_41[13], stage1_41[14]},
      {stage1_42[44]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[9],stage2_43[9],stage2_42[11],stage2_41[26]}
   );
   gpc615_5 gpc1794 (
      {stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19]},
      {stage1_42[45]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[10],stage2_43[10],stage2_42[12],stage2_41[27]}
   );
   gpc615_5 gpc1795 (
      {stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24]},
      {stage1_42[46]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[11],stage2_43[11],stage2_42[13],stage2_41[28]}
   );
   gpc615_5 gpc1796 (
      {stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage1_42[47]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[12],stage2_43[12],stage2_42[14],stage2_41[29]}
   );
   gpc615_5 gpc1797 (
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34]},
      {stage1_42[48]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[13],stage2_43[13],stage2_42[15],stage2_41[30]}
   );
   gpc615_5 gpc1798 (
      {stage1_41[35], stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39]},
      {stage1_42[49]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[14],stage2_43[14],stage2_42[16],stage2_41[31]}
   );
   gpc606_5 gpc1799 (
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[8],stage2_44[15],stage2_43[15]}
   );
   gpc606_5 gpc1800 (
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[9],stage2_44[16],stage2_43[16]}
   );
   gpc606_5 gpc1801 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[10],stage2_44[17],stage2_43[17]}
   );
   gpc606_5 gpc1802 (
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[3],stage2_45[11],stage2_44[18],stage2_43[18]}
   );
   gpc606_5 gpc1803 (
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[4],stage2_45[12],stage2_44[19],stage2_43[19]}
   );
   gpc615_5 gpc1804 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[30]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[5],stage2_46[5],stage2_45[13],stage2_44[20]}
   );
   gpc615_5 gpc1805 (
      {stage1_44[5], stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9]},
      {stage1_45[31]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[6],stage2_46[6],stage2_45[14],stage2_44[21]}
   );
   gpc615_5 gpc1806 (
      {stage1_44[10], stage1_44[11], stage1_44[12], stage1_44[13], stage1_44[14]},
      {stage1_45[32]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[7],stage2_46[7],stage2_45[15],stage2_44[22]}
   );
   gpc615_5 gpc1807 (
      {stage1_44[15], stage1_44[16], stage1_44[17], stage1_44[18], stage1_44[19]},
      {stage1_45[33]},
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage2_48[3],stage2_47[8],stage2_46[8],stage2_45[16],stage2_44[23]}
   );
   gpc615_5 gpc1808 (
      {stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23], stage1_44[24]},
      {stage1_45[34]},
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage2_48[4],stage2_47[9],stage2_46[9],stage2_45[17],stage2_44[24]}
   );
   gpc615_5 gpc1809 (
      {stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage1_45[35]},
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage2_48[5],stage2_47[10],stage2_46[10],stage2_45[18],stage2_44[25]}
   );
   gpc615_5 gpc1810 (
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34]},
      {stage1_45[36]},
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage2_48[6],stage2_47[11],stage2_46[11],stage2_45[19],stage2_44[26]}
   );
   gpc615_5 gpc1811 (
      {stage1_44[35], stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39]},
      {stage1_45[37]},
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage2_48[7],stage2_47[12],stage2_46[12],stage2_45[20],stage2_44[27]}
   );
   gpc615_5 gpc1812 (
      {stage1_44[40], stage1_44[41], stage1_44[42], stage1_44[43], stage1_44[44]},
      {stage1_45[38]},
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage2_48[8],stage2_47[13],stage2_46[13],stage2_45[21],stage2_44[28]}
   );
   gpc615_5 gpc1813 (
      {stage1_44[45], stage1_44[46], stage1_44[47], stage1_44[48], stage1_44[49]},
      {stage1_45[39]},
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage2_48[9],stage2_47[14],stage2_46[14],stage2_45[22],stage2_44[29]}
   );
   gpc117_4 gpc1814 (
      {stage1_45[40], stage1_45[41], stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46]},
      {stage1_46[60]},
      {stage1_47[0]},
      {stage2_48[10],stage2_47[15],stage2_46[15],stage2_45[23]}
   );
   gpc615_5 gpc1815 (
      {stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage1_47[1]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[0],stage2_48[11],stage2_47[16],stage2_46[16]}
   );
   gpc615_5 gpc1816 (
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70]},
      {stage1_47[2]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[1],stage2_48[12],stage2_47[17],stage2_46[17]}
   );
   gpc615_5 gpc1817 (
      {stage1_46[71], stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75]},
      {stage1_47[3]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[2],stage2_48[13],stage2_47[18],stage2_46[18]}
   );
   gpc2135_5 gpc1818 (
      {stage1_47[4], stage1_47[5], stage1_47[6], stage1_47[7], stage1_47[8]},
      {stage1_48[18], stage1_48[19], stage1_48[20]},
      {stage1_49[0]},
      {stage1_50[0], stage1_50[1]},
      {stage2_51[0],stage2_50[3],stage2_49[3],stage2_48[14],stage2_47[19]}
   );
   gpc2135_5 gpc1819 (
      {stage1_47[9], stage1_47[10], stage1_47[11], stage1_47[12], stage1_47[13]},
      {stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage1_49[1]},
      {stage1_50[2], stage1_50[3]},
      {stage2_51[1],stage2_50[4],stage2_49[4],stage2_48[15],stage2_47[20]}
   );
   gpc2135_5 gpc1820 (
      {stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17], stage1_47[18]},
      {stage1_48[24], stage1_48[25], stage1_48[26]},
      {stage1_49[2]},
      {stage1_50[4], stage1_50[5]},
      {stage2_51[2],stage2_50[5],stage2_49[5],stage2_48[16],stage2_47[21]}
   );
   gpc606_5 gpc1821 (
      {stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23], stage1_47[24]},
      {stage1_49[3], stage1_49[4], stage1_49[5], stage1_49[6], stage1_49[7], stage1_49[8]},
      {stage2_51[3],stage2_50[6],stage2_49[6],stage2_48[17],stage2_47[22]}
   );
   gpc606_5 gpc1822 (
      {stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29], stage1_47[30]},
      {stage1_49[9], stage1_49[10], stage1_49[11], stage1_49[12], stage1_49[13], stage1_49[14]},
      {stage2_51[4],stage2_50[7],stage2_49[7],stage2_48[18],stage2_47[23]}
   );
   gpc606_5 gpc1823 (
      {stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35], stage1_47[36]},
      {stage1_49[15], stage1_49[16], stage1_49[17], stage1_49[18], stage1_49[19], stage1_49[20]},
      {stage2_51[5],stage2_50[8],stage2_49[8],stage2_48[19],stage2_47[24]}
   );
   gpc606_5 gpc1824 (
      {stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41], stage1_47[42]},
      {stage1_49[21], stage1_49[22], stage1_49[23], stage1_49[24], stage1_49[25], stage1_49[26]},
      {stage2_51[6],stage2_50[9],stage2_49[9],stage2_48[20],stage2_47[25]}
   );
   gpc606_5 gpc1825 (
      {stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47], stage1_47[48]},
      {stage1_49[27], stage1_49[28], stage1_49[29], stage1_49[30], stage1_49[31], stage1_49[32]},
      {stage2_51[7],stage2_50[10],stage2_49[10],stage2_48[21],stage2_47[26]}
   );
   gpc615_5 gpc1826 (
      {stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage1_48[27]},
      {stage1_49[33], stage1_49[34], stage1_49[35], stage1_49[36], stage1_49[37], stage1_49[38]},
      {stage2_51[8],stage2_50[11],stage2_49[11],stage2_48[22],stage2_47[27]}
   );
   gpc615_5 gpc1827 (
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58]},
      {stage1_48[28]},
      {stage1_49[39], stage1_49[40], stage1_49[41], stage1_49[42], stage1_49[43], stage1_49[44]},
      {stage2_51[9],stage2_50[12],stage2_49[12],stage2_48[23],stage2_47[28]}
   );
   gpc615_5 gpc1828 (
      {stage1_47[59], stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63]},
      {stage1_48[29]},
      {stage1_49[45], stage1_49[46], stage1_49[47], stage1_49[48], stage1_49[49], stage1_49[50]},
      {stage2_51[10],stage2_50[13],stage2_49[13],stage2_48[24],stage2_47[29]}
   );
   gpc606_5 gpc1829 (
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[0],stage2_51[11],stage2_50[14],stage2_49[14],stage2_48[25]}
   );
   gpc606_5 gpc1830 (
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[1],stage2_51[12],stage2_50[15],stage2_49[15],stage2_48[26]}
   );
   gpc1163_5 gpc1831 (
      {stage1_50[18], stage1_50[19], stage1_50[20]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[0]},
      {stage1_53[0]},
      {stage2_54[0],stage2_53[0],stage2_52[2],stage2_51[13],stage2_50[16]}
   );
   gpc1163_5 gpc1832 (
      {stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage1_52[1]},
      {stage1_53[1]},
      {stage2_54[1],stage2_53[1],stage2_52[3],stage2_51[14],stage2_50[17]}
   );
   gpc1163_5 gpc1833 (
      {stage1_50[24], stage1_50[25], stage1_50[26]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage1_52[2]},
      {stage1_53[2]},
      {stage2_54[2],stage2_53[2],stage2_52[4],stage2_51[15],stage2_50[18]}
   );
   gpc1163_5 gpc1834 (
      {stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage1_52[3]},
      {stage1_53[3]},
      {stage2_54[3],stage2_53[3],stage2_52[5],stage2_51[16],stage2_50[19]}
   );
   gpc1163_5 gpc1835 (
      {stage1_50[30], stage1_50[31], stage1_50[32]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage1_52[4]},
      {stage1_53[4]},
      {stage2_54[4],stage2_53[4],stage2_52[6],stage2_51[17],stage2_50[20]}
   );
   gpc1163_5 gpc1836 (
      {stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage1_52[5]},
      {stage1_53[5]},
      {stage2_54[5],stage2_53[5],stage2_52[7],stage2_51[18],stage2_50[21]}
   );
   gpc615_5 gpc1837 (
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40]},
      {stage1_51[36]},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage2_54[6],stage2_53[6],stage2_52[8],stage2_51[19],stage2_50[22]}
   );
   gpc615_5 gpc1838 (
      {stage1_50[41], stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45]},
      {stage1_51[37]},
      {stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17]},
      {stage2_54[7],stage2_53[7],stage2_52[9],stage2_51[20],stage2_50[23]}
   );
   gpc615_5 gpc1839 (
      {stage1_50[46], stage1_50[47], stage1_50[48], stage1_50[49], stage1_50[50]},
      {stage1_51[38]},
      {stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23]},
      {stage2_54[8],stage2_53[8],stage2_52[10],stage2_51[21],stage2_50[24]}
   );
   gpc615_5 gpc1840 (
      {stage1_50[51], stage1_50[52], stage1_50[53], stage1_50[54], stage1_50[55]},
      {stage1_51[39]},
      {stage1_52[24], stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29]},
      {stage2_54[9],stage2_53[9],stage2_52[11],stage2_51[22],stage2_50[25]}
   );
   gpc615_5 gpc1841 (
      {stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59], stage1_50[60]},
      {stage1_51[40]},
      {stage1_52[30], stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35]},
      {stage2_54[10],stage2_53[10],stage2_52[12],stage2_51[23],stage2_50[26]}
   );
   gpc615_5 gpc1842 (
      {stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage1_51[41]},
      {stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41]},
      {stage2_54[11],stage2_53[11],stage2_52[13],stage2_51[24],stage2_50[27]}
   );
   gpc606_5 gpc1843 (
      {stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[0],stage2_54[12],stage2_53[12],stage2_52[14]}
   );
   gpc606_5 gpc1844 (
      {stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[1],stage2_54[13],stage2_53[13],stage2_52[15]}
   );
   gpc606_5 gpc1845 (
      {stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[2],stage2_54[14],stage2_53[14],stage2_52[16]}
   );
   gpc606_5 gpc1846 (
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[3],stage2_55[3],stage2_54[15],stage2_53[15]}
   );
   gpc606_5 gpc1847 (
      {stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16], stage1_53[17]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[4],stage2_55[4],stage2_54[16],stage2_53[16]}
   );
   gpc606_5 gpc1848 (
      {stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[5],stage2_55[5],stage2_54[17],stage2_53[17]}
   );
   gpc606_5 gpc1849 (
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[6],stage2_55[6],stage2_54[18],stage2_53[18]}
   );
   gpc615_5 gpc1850 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage1_54[18]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[7],stage2_55[7],stage2_54[19],stage2_53[19]}
   );
   gpc615_5 gpc1851 (
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage1_54[19]},
      {stage1_55[30], stage1_55[31], stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35]},
      {stage2_57[5],stage2_56[8],stage2_55[8],stage2_54[20],stage2_53[20]}
   );
   gpc615_5 gpc1852 (
      {stage1_53[40], stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44]},
      {stage1_54[20]},
      {stage1_55[36], stage1_55[37], stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41]},
      {stage2_57[6],stage2_56[9],stage2_55[9],stage2_54[21],stage2_53[21]}
   );
   gpc615_5 gpc1853 (
      {stage1_54[21], stage1_54[22], stage1_54[23], stage1_54[24], stage1_54[25]},
      {stage1_55[42]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[7],stage2_56[10],stage2_55[10],stage2_54[22]}
   );
   gpc615_5 gpc1854 (
      {stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29], stage1_54[30]},
      {stage1_55[43]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[8],stage2_56[11],stage2_55[11],stage2_54[23]}
   );
   gpc615_5 gpc1855 (
      {stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage1_55[44]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[9],stage2_56[12],stage2_55[12],stage2_54[24]}
   );
   gpc615_5 gpc1856 (
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40]},
      {stage1_55[45]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[10],stage2_56[13],stage2_55[13],stage2_54[25]}
   );
   gpc615_5 gpc1857 (
      {stage1_54[41], stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45]},
      {stage1_55[46]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[11],stage2_56[14],stage2_55[14],stage2_54[26]}
   );
   gpc615_5 gpc1858 (
      {stage1_54[46], stage1_54[47], stage1_54[48], stage1_54[49], stage1_54[50]},
      {stage1_55[47]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[12],stage2_56[15],stage2_55[15],stage2_54[27]}
   );
   gpc615_5 gpc1859 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[36]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[6],stage2_57[13],stage2_56[16],stage2_55[16]}
   );
   gpc615_5 gpc1860 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[37]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[7],stage2_57[14],stage2_56[17],stage2_55[17]}
   );
   gpc615_5 gpc1861 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[38]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[8],stage2_57[15],stage2_56[18],stage2_55[18]}
   );
   gpc615_5 gpc1862 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[39]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[9],stage2_57[16],stage2_56[19],stage2_55[19]}
   );
   gpc606_5 gpc1863 (
      {stage1_56[40], stage1_56[41], stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[4],stage2_58[10],stage2_57[17],stage2_56[20]}
   );
   gpc606_5 gpc1864 (
      {stage1_56[46], stage1_56[47], stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[5],stage2_58[11],stage2_57[18],stage2_56[21]}
   );
   gpc606_5 gpc1865 (
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[2],stage2_59[6],stage2_58[12],stage2_57[19]}
   );
   gpc606_5 gpc1866 (
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[3],stage2_59[7],stage2_58[13],stage2_57[20]}
   );
   gpc606_5 gpc1867 (
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[4],stage2_59[8],stage2_58[14],stage2_57[21]}
   );
   gpc606_5 gpc1868 (
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[5],stage2_59[9],stage2_58[15],stage2_57[22]}
   );
   gpc606_5 gpc1869 (
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[4],stage2_60[6],stage2_59[10],stage2_58[16]}
   );
   gpc606_5 gpc1870 (
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[5],stage2_60[7],stage2_59[11],stage2_58[17]}
   );
   gpc606_5 gpc1871 (
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[6],stage2_60[8],stage2_59[12],stage2_58[18]}
   );
   gpc606_5 gpc1872 (
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[7],stage2_60[9],stage2_59[13],stage2_58[19]}
   );
   gpc606_5 gpc1873 (
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[8],stage2_60[10],stage2_59[14],stage2_58[20]}
   );
   gpc606_5 gpc1874 (
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage2_62[5],stage2_61[9],stage2_60[11],stage2_59[15],stage2_58[21]}
   );
   gpc606_5 gpc1875 (
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage2_62[6],stage2_61[10],stage2_60[12],stage2_59[16],stage2_58[22]}
   );
   gpc606_5 gpc1876 (
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage2_62[7],stage2_61[11],stage2_60[13],stage2_59[17],stage2_58[23]}
   );
   gpc606_5 gpc1877 (
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[8],stage2_61[12],stage2_60[14],stage2_59[18]}
   );
   gpc606_5 gpc1878 (
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[9],stage2_61[13],stage2_60[15],stage2_59[19]}
   );
   gpc606_5 gpc1879 (
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[10],stage2_61[14],stage2_60[16],stage2_59[20]}
   );
   gpc1163_5 gpc1880 (
      {stage1_61[18], stage1_61[19], stage1_61[20]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage1_63[0]},
      {stage1_64[0]},
      {stage2_65[0],stage2_64[0],stage2_63[3],stage2_62[11],stage2_61[15]}
   );
   gpc1163_5 gpc1881 (
      {stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage1_63[1]},
      {stage1_64[1]},
      {stage2_65[1],stage2_64[1],stage2_63[4],stage2_62[12],stage2_61[16]}
   );
   gpc1163_5 gpc1882 (
      {stage1_61[24], stage1_61[25], stage1_61[26]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage1_63[2]},
      {stage1_64[2]},
      {stage2_65[2],stage2_64[2],stage2_63[5],stage2_62[13],stage2_61[17]}
   );
   gpc1163_5 gpc1883 (
      {stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage1_63[3]},
      {stage1_64[3]},
      {stage2_65[3],stage2_64[3],stage2_63[6],stage2_62[14],stage2_61[18]}
   );
   gpc1163_5 gpc1884 (
      {stage1_61[30], stage1_61[31], stage1_61[32]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage1_63[4]},
      {stage1_64[4]},
      {stage2_65[4],stage2_64[4],stage2_63[7],stage2_62[15],stage2_61[19]}
   );
   gpc1163_5 gpc1885 (
      {stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage1_63[5]},
      {stage1_64[5]},
      {stage2_65[5],stage2_64[5],stage2_63[8],stage2_62[16],stage2_61[20]}
   );
   gpc1163_5 gpc1886 (
      {stage1_61[36], stage1_61[37], stage1_61[38]},
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41]},
      {stage1_63[6]},
      {stage1_64[6]},
      {stage2_65[6],stage2_64[6],stage2_63[9],stage2_62[17],stage2_61[21]}
   );
   gpc1163_5 gpc1887 (
      {stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47]},
      {stage1_63[7]},
      {stage1_64[7]},
      {stage2_65[7],stage2_64[7],stage2_63[10],stage2_62[18],stage2_61[22]}
   );
   gpc1163_5 gpc1888 (
      {stage1_61[42], stage1_61[43], stage1_61[44]},
      {stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53]},
      {stage1_63[8]},
      {stage1_64[8]},
      {stage2_65[8],stage2_64[8],stage2_63[11],stage2_62[19],stage2_61[23]}
   );
   gpc1163_5 gpc1889 (
      {stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59]},
      {stage1_63[9]},
      {stage1_64[9]},
      {stage2_65[9],stage2_64[9],stage2_63[12],stage2_62[20],stage2_61[24]}
   );
   gpc1163_5 gpc1890 (
      {stage1_61[48], stage1_61[49], stage1_61[50]},
      {stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage1_63[10]},
      {stage1_64[10]},
      {stage2_65[10],stage2_64[10],stage2_63[13],stage2_62[21],stage2_61[25]}
   );
   gpc606_5 gpc1891 (
      {stage1_61[51], stage1_61[52], stage1_61[53], stage1_61[54], stage1_61[55], stage1_61[56]},
      {stage1_63[11], stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16]},
      {stage2_65[11],stage2_64[11],stage2_63[14],stage2_62[22],stage2_61[26]}
   );
   gpc2135_5 gpc1892 (
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70]},
      {stage1_63[17], stage1_63[18], stage1_63[19]},
      {stage1_64[11]},
      {stage1_65[0], stage1_65[1]},
      {stage2_66[0],stage2_65[12],stage2_64[12],stage2_63[15],stage2_62[23]}
   );
   gpc2135_5 gpc1893 (
      {stage1_62[71], stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75]},
      {stage1_63[20], stage1_63[21], stage1_63[22]},
      {stage1_64[12]},
      {stage1_65[2], stage1_65[3]},
      {stage2_66[1],stage2_65[13],stage2_64[13],stage2_63[16],stage2_62[24]}
   );
   gpc2135_5 gpc1894 (
      {stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79], stage1_62[80]},
      {stage1_63[23], stage1_63[24], stage1_63[25]},
      {stage1_64[13]},
      {stage1_65[4], stage1_65[5]},
      {stage2_66[2],stage2_65[14],stage2_64[14],stage2_63[17],stage2_62[25]}
   );
   gpc606_5 gpc1895 (
      {stage1_62[81], stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85], stage1_62[86]},
      {stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17], stage1_64[18], stage1_64[19]},
      {stage2_66[3],stage2_65[15],stage2_64[15],stage2_63[18],stage2_62[26]}
   );
   gpc615_5 gpc1896 (
      {stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29], stage1_63[30]},
      {stage1_64[20]},
      {stage1_65[6], stage1_65[7], stage1_65[8], stage1_65[9], stage1_65[10], stage1_65[11]},
      {stage2_67[0],stage2_66[4],stage2_65[16],stage2_64[16],stage2_63[19]}
   );
   gpc615_5 gpc1897 (
      {stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_64[21]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[1],stage2_66[5],stage2_65[17],stage2_64[17],stage2_63[20]}
   );
   gpc1_1 gpc1898 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc1899 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc1900 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc1901 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc1902 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc1903 (
      {stage1_0[18]},
      {stage2_0[8]}
   );
   gpc1_1 gpc1904 (
      {stage1_0[19]},
      {stage2_0[9]}
   );
   gpc1_1 gpc1905 (
      {stage1_0[20]},
      {stage2_0[10]}
   );
   gpc1_1 gpc1906 (
      {stage1_0[21]},
      {stage2_0[11]}
   );
   gpc1_1 gpc1907 (
      {stage1_0[22]},
      {stage2_0[12]}
   );
   gpc1_1 gpc1908 (
      {stage1_0[23]},
      {stage2_0[13]}
   );
   gpc1_1 gpc1909 (
      {stage1_0[24]},
      {stage2_0[14]}
   );
   gpc1_1 gpc1910 (
      {stage1_0[25]},
      {stage2_0[15]}
   );
   gpc1_1 gpc1911 (
      {stage1_0[26]},
      {stage2_0[16]}
   );
   gpc1_1 gpc1912 (
      {stage1_0[27]},
      {stage2_0[17]}
   );
   gpc1_1 gpc1913 (
      {stage1_0[28]},
      {stage2_0[18]}
   );
   gpc1_1 gpc1914 (
      {stage1_0[29]},
      {stage2_0[19]}
   );
   gpc1_1 gpc1915 (
      {stage1_1[26]},
      {stage2_1[6]}
   );
   gpc1_1 gpc1916 (
      {stage1_1[27]},
      {stage2_1[7]}
   );
   gpc1_1 gpc1917 (
      {stage1_1[28]},
      {stage2_1[8]}
   );
   gpc1_1 gpc1918 (
      {stage1_1[29]},
      {stage2_1[9]}
   );
   gpc1_1 gpc1919 (
      {stage1_1[30]},
      {stage2_1[10]}
   );
   gpc1_1 gpc1920 (
      {stage1_1[31]},
      {stage2_1[11]}
   );
   gpc1_1 gpc1921 (
      {stage1_1[32]},
      {stage2_1[12]}
   );
   gpc1_1 gpc1922 (
      {stage1_2[31]},
      {stage2_2[9]}
   );
   gpc1_1 gpc1923 (
      {stage1_2[32]},
      {stage2_2[10]}
   );
   gpc1_1 gpc1924 (
      {stage1_2[33]},
      {stage2_2[11]}
   );
   gpc1_1 gpc1925 (
      {stage1_2[34]},
      {stage2_2[12]}
   );
   gpc1_1 gpc1926 (
      {stage1_2[35]},
      {stage2_2[13]}
   );
   gpc1_1 gpc1927 (
      {stage1_2[36]},
      {stage2_2[14]}
   );
   gpc1_1 gpc1928 (
      {stage1_2[37]},
      {stage2_2[15]}
   );
   gpc1_1 gpc1929 (
      {stage1_2[38]},
      {stage2_2[16]}
   );
   gpc1_1 gpc1930 (
      {stage1_2[39]},
      {stage2_2[17]}
   );
   gpc1_1 gpc1931 (
      {stage1_2[40]},
      {stage2_2[18]}
   );
   gpc1_1 gpc1932 (
      {stage1_2[41]},
      {stage2_2[19]}
   );
   gpc1_1 gpc1933 (
      {stage1_2[42]},
      {stage2_2[20]}
   );
   gpc1_1 gpc1934 (
      {stage1_2[43]},
      {stage2_2[21]}
   );
   gpc1_1 gpc1935 (
      {stage1_2[44]},
      {stage2_2[22]}
   );
   gpc1_1 gpc1936 (
      {stage1_2[45]},
      {stage2_2[23]}
   );
   gpc1_1 gpc1937 (
      {stage1_2[46]},
      {stage2_2[24]}
   );
   gpc1_1 gpc1938 (
      {stage1_3[55]},
      {stage2_3[16]}
   );
   gpc1_1 gpc1939 (
      {stage1_3[56]},
      {stage2_3[17]}
   );
   gpc1_1 gpc1940 (
      {stage1_3[57]},
      {stage2_3[18]}
   );
   gpc1_1 gpc1941 (
      {stage1_3[58]},
      {stage2_3[19]}
   );
   gpc1_1 gpc1942 (
      {stage1_3[59]},
      {stage2_3[20]}
   );
   gpc1_1 gpc1943 (
      {stage1_3[60]},
      {stage2_3[21]}
   );
   gpc1_1 gpc1944 (
      {stage1_3[61]},
      {stage2_3[22]}
   );
   gpc1_1 gpc1945 (
      {stage1_3[62]},
      {stage2_3[23]}
   );
   gpc1_1 gpc1946 (
      {stage1_3[63]},
      {stage2_3[24]}
   );
   gpc1_1 gpc1947 (
      {stage1_3[64]},
      {stage2_3[25]}
   );
   gpc1_1 gpc1948 (
      {stage1_3[65]},
      {stage2_3[26]}
   );
   gpc1_1 gpc1949 (
      {stage1_3[66]},
      {stage2_3[27]}
   );
   gpc1_1 gpc1950 (
      {stage1_4[63]},
      {stage2_4[23]}
   );
   gpc1_1 gpc1951 (
      {stage1_4[64]},
      {stage2_4[24]}
   );
   gpc1_1 gpc1952 (
      {stage1_4[65]},
      {stage2_4[25]}
   );
   gpc1_1 gpc1953 (
      {stage1_5[43]},
      {stage2_5[20]}
   );
   gpc1_1 gpc1954 (
      {stage1_5[44]},
      {stage2_5[21]}
   );
   gpc1_1 gpc1955 (
      {stage1_5[45]},
      {stage2_5[22]}
   );
   gpc1_1 gpc1956 (
      {stage1_5[46]},
      {stage2_5[23]}
   );
   gpc1_1 gpc1957 (
      {stage1_5[47]},
      {stage2_5[24]}
   );
   gpc1_1 gpc1958 (
      {stage1_5[48]},
      {stage2_5[25]}
   );
   gpc1_1 gpc1959 (
      {stage1_5[49]},
      {stage2_5[26]}
   );
   gpc1_1 gpc1960 (
      {stage1_5[50]},
      {stage2_5[27]}
   );
   gpc1_1 gpc1961 (
      {stage1_5[51]},
      {stage2_5[28]}
   );
   gpc1_1 gpc1962 (
      {stage1_7[64]},
      {stage2_7[32]}
   );
   gpc1_1 gpc1963 (
      {stage1_7[65]},
      {stage2_7[33]}
   );
   gpc1_1 gpc1964 (
      {stage1_7[66]},
      {stage2_7[34]}
   );
   gpc1_1 gpc1965 (
      {stage1_7[67]},
      {stage2_7[35]}
   );
   gpc1_1 gpc1966 (
      {stage1_7[68]},
      {stage2_7[36]}
   );
   gpc1_1 gpc1967 (
      {stage1_7[69]},
      {stage2_7[37]}
   );
   gpc1_1 gpc1968 (
      {stage1_7[70]},
      {stage2_7[38]}
   );
   gpc1_1 gpc1969 (
      {stage1_8[59]},
      {stage2_8[25]}
   );
   gpc1_1 gpc1970 (
      {stage1_8[60]},
      {stage2_8[26]}
   );
   gpc1_1 gpc1971 (
      {stage1_8[61]},
      {stage2_8[27]}
   );
   gpc1_1 gpc1972 (
      {stage1_8[62]},
      {stage2_8[28]}
   );
   gpc1_1 gpc1973 (
      {stage1_8[63]},
      {stage2_8[29]}
   );
   gpc1_1 gpc1974 (
      {stage1_8[64]},
      {stage2_8[30]}
   );
   gpc1_1 gpc1975 (
      {stage1_8[65]},
      {stage2_8[31]}
   );
   gpc1_1 gpc1976 (
      {stage1_9[38]},
      {stage2_9[19]}
   );
   gpc1_1 gpc1977 (
      {stage1_9[39]},
      {stage2_9[20]}
   );
   gpc1_1 gpc1978 (
      {stage1_9[40]},
      {stage2_9[21]}
   );
   gpc1_1 gpc1979 (
      {stage1_9[41]},
      {stage2_9[22]}
   );
   gpc1_1 gpc1980 (
      {stage1_9[42]},
      {stage2_9[23]}
   );
   gpc1_1 gpc1981 (
      {stage1_9[43]},
      {stage2_9[24]}
   );
   gpc1_1 gpc1982 (
      {stage1_9[44]},
      {stage2_9[25]}
   );
   gpc1_1 gpc1983 (
      {stage1_9[45]},
      {stage2_9[26]}
   );
   gpc1_1 gpc1984 (
      {stage1_9[46]},
      {stage2_9[27]}
   );
   gpc1_1 gpc1985 (
      {stage1_9[47]},
      {stage2_9[28]}
   );
   gpc1_1 gpc1986 (
      {stage1_9[48]},
      {stage2_9[29]}
   );
   gpc1_1 gpc1987 (
      {stage1_9[49]},
      {stage2_9[30]}
   );
   gpc1_1 gpc1988 (
      {stage1_9[50]},
      {stage2_9[31]}
   );
   gpc1_1 gpc1989 (
      {stage1_9[51]},
      {stage2_9[32]}
   );
   gpc1_1 gpc1990 (
      {stage1_9[52]},
      {stage2_9[33]}
   );
   gpc1_1 gpc1991 (
      {stage1_9[53]},
      {stage2_9[34]}
   );
   gpc1_1 gpc1992 (
      {stage1_9[54]},
      {stage2_9[35]}
   );
   gpc1_1 gpc1993 (
      {stage1_9[55]},
      {stage2_9[36]}
   );
   gpc1_1 gpc1994 (
      {stage1_9[56]},
      {stage2_9[37]}
   );
   gpc1_1 gpc1995 (
      {stage1_9[57]},
      {stage2_9[38]}
   );
   gpc1_1 gpc1996 (
      {stage1_9[58]},
      {stage2_9[39]}
   );
   gpc1_1 gpc1997 (
      {stage1_9[59]},
      {stage2_9[40]}
   );
   gpc1_1 gpc1998 (
      {stage1_9[60]},
      {stage2_9[41]}
   );
   gpc1_1 gpc1999 (
      {stage1_10[36]},
      {stage2_10[26]}
   );
   gpc1_1 gpc2000 (
      {stage1_10[37]},
      {stage2_10[27]}
   );
   gpc1_1 gpc2001 (
      {stage1_10[38]},
      {stage2_10[28]}
   );
   gpc1_1 gpc2002 (
      {stage1_10[39]},
      {stage2_10[29]}
   );
   gpc1_1 gpc2003 (
      {stage1_10[40]},
      {stage2_10[30]}
   );
   gpc1_1 gpc2004 (
      {stage1_12[45]},
      {stage2_12[17]}
   );
   gpc1_1 gpc2005 (
      {stage1_12[46]},
      {stage2_12[18]}
   );
   gpc1_1 gpc2006 (
      {stage1_12[47]},
      {stage2_12[19]}
   );
   gpc1_1 gpc2007 (
      {stage1_12[48]},
      {stage2_12[20]}
   );
   gpc1_1 gpc2008 (
      {stage1_12[49]},
      {stage2_12[21]}
   );
   gpc1_1 gpc2009 (
      {stage1_12[50]},
      {stage2_12[22]}
   );
   gpc1_1 gpc2010 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc2011 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc2012 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc2013 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc2014 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc2015 (
      {stage1_14[53]},
      {stage2_14[26]}
   );
   gpc1_1 gpc2016 (
      {stage1_14[54]},
      {stage2_14[27]}
   );
   gpc1_1 gpc2017 (
      {stage1_14[55]},
      {stage2_14[28]}
   );
   gpc1_1 gpc2018 (
      {stage1_14[56]},
      {stage2_14[29]}
   );
   gpc1_1 gpc2019 (
      {stage1_14[57]},
      {stage2_14[30]}
   );
   gpc1_1 gpc2020 (
      {stage1_14[58]},
      {stage2_14[31]}
   );
   gpc1_1 gpc2021 (
      {stage1_14[59]},
      {stage2_14[32]}
   );
   gpc1_1 gpc2022 (
      {stage1_14[60]},
      {stage2_14[33]}
   );
   gpc1_1 gpc2023 (
      {stage1_14[61]},
      {stage2_14[34]}
   );
   gpc1_1 gpc2024 (
      {stage1_14[62]},
      {stage2_14[35]}
   );
   gpc1_1 gpc2025 (
      {stage1_14[63]},
      {stage2_14[36]}
   );
   gpc1_1 gpc2026 (
      {stage1_14[64]},
      {stage2_14[37]}
   );
   gpc1_1 gpc2027 (
      {stage1_14[65]},
      {stage2_14[38]}
   );
   gpc1_1 gpc2028 (
      {stage1_15[67]},
      {stage2_15[30]}
   );
   gpc1_1 gpc2029 (
      {stage1_17[62]},
      {stage2_17[29]}
   );
   gpc1_1 gpc2030 (
      {stage1_17[63]},
      {stage2_17[30]}
   );
   gpc1_1 gpc2031 (
      {stage1_17[64]},
      {stage2_17[31]}
   );
   gpc1_1 gpc2032 (
      {stage1_17[65]},
      {stage2_17[32]}
   );
   gpc1_1 gpc2033 (
      {stage1_17[66]},
      {stage2_17[33]}
   );
   gpc1_1 gpc2034 (
      {stage1_18[40]},
      {stage2_18[29]}
   );
   gpc1_1 gpc2035 (
      {stage1_18[41]},
      {stage2_18[30]}
   );
   gpc1_1 gpc2036 (
      {stage1_19[54]},
      {stage2_19[26]}
   );
   gpc1_1 gpc2037 (
      {stage1_20[62]},
      {stage2_20[24]}
   );
   gpc1_1 gpc2038 (
      {stage1_20[63]},
      {stage2_20[25]}
   );
   gpc1_1 gpc2039 (
      {stage1_20[64]},
      {stage2_20[26]}
   );
   gpc1_1 gpc2040 (
      {stage1_20[65]},
      {stage2_20[27]}
   );
   gpc1_1 gpc2041 (
      {stage1_20[66]},
      {stage2_20[28]}
   );
   gpc1_1 gpc2042 (
      {stage1_20[67]},
      {stage2_20[29]}
   );
   gpc1_1 gpc2043 (
      {stage1_20[68]},
      {stage2_20[30]}
   );
   gpc1_1 gpc2044 (
      {stage1_20[69]},
      {stage2_20[31]}
   );
   gpc1_1 gpc2045 (
      {stage1_20[70]},
      {stage2_20[32]}
   );
   gpc1_1 gpc2046 (
      {stage1_20[71]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2047 (
      {stage1_22[54]},
      {stage2_22[18]}
   );
   gpc1_1 gpc2048 (
      {stage1_22[55]},
      {stage2_22[19]}
   );
   gpc1_1 gpc2049 (
      {stage1_22[56]},
      {stage2_22[20]}
   );
   gpc1_1 gpc2050 (
      {stage1_22[57]},
      {stage2_22[21]}
   );
   gpc1_1 gpc2051 (
      {stage1_22[58]},
      {stage2_22[22]}
   );
   gpc1_1 gpc2052 (
      {stage1_22[59]},
      {stage2_22[23]}
   );
   gpc1_1 gpc2053 (
      {stage1_22[60]},
      {stage2_22[24]}
   );
   gpc1_1 gpc2054 (
      {stage1_22[61]},
      {stage2_22[25]}
   );
   gpc1_1 gpc2055 (
      {stage1_22[62]},
      {stage2_22[26]}
   );
   gpc1_1 gpc2056 (
      {stage1_22[63]},
      {stage2_22[27]}
   );
   gpc1_1 gpc2057 (
      {stage1_22[64]},
      {stage2_22[28]}
   );
   gpc1_1 gpc2058 (
      {stage1_22[65]},
      {stage2_22[29]}
   );
   gpc1_1 gpc2059 (
      {stage1_22[66]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2060 (
      {stage1_22[67]},
      {stage2_22[31]}
   );
   gpc1_1 gpc2061 (
      {stage1_22[68]},
      {stage2_22[32]}
   );
   gpc1_1 gpc2062 (
      {stage1_22[69]},
      {stage2_22[33]}
   );
   gpc1_1 gpc2063 (
      {stage1_22[70]},
      {stage2_22[34]}
   );
   gpc1_1 gpc2064 (
      {stage1_23[52]},
      {stage2_23[26]}
   );
   gpc1_1 gpc2065 (
      {stage1_23[53]},
      {stage2_23[27]}
   );
   gpc1_1 gpc2066 (
      {stage1_25[48]},
      {stage2_25[19]}
   );
   gpc1_1 gpc2067 (
      {stage1_25[49]},
      {stage2_25[20]}
   );
   gpc1_1 gpc2068 (
      {stage1_25[50]},
      {stage2_25[21]}
   );
   gpc1_1 gpc2069 (
      {stage1_25[51]},
      {stage2_25[22]}
   );
   gpc1_1 gpc2070 (
      {stage1_25[52]},
      {stage2_25[23]}
   );
   gpc1_1 gpc2071 (
      {stage1_25[53]},
      {stage2_25[24]}
   );
   gpc1_1 gpc2072 (
      {stage1_25[54]},
      {stage2_25[25]}
   );
   gpc1_1 gpc2073 (
      {stage1_25[55]},
      {stage2_25[26]}
   );
   gpc1_1 gpc2074 (
      {stage1_25[56]},
      {stage2_25[27]}
   );
   gpc1_1 gpc2075 (
      {stage1_25[57]},
      {stage2_25[28]}
   );
   gpc1_1 gpc2076 (
      {stage1_25[58]},
      {stage2_25[29]}
   );
   gpc1_1 gpc2077 (
      {stage1_25[59]},
      {stage2_25[30]}
   );
   gpc1_1 gpc2078 (
      {stage1_25[60]},
      {stage2_25[31]}
   );
   gpc1_1 gpc2079 (
      {stage1_26[79]},
      {stage2_26[22]}
   );
   gpc1_1 gpc2080 (
      {stage1_26[80]},
      {stage2_26[23]}
   );
   gpc1_1 gpc2081 (
      {stage1_26[81]},
      {stage2_26[24]}
   );
   gpc1_1 gpc2082 (
      {stage1_26[82]},
      {stage2_26[25]}
   );
   gpc1_1 gpc2083 (
      {stage1_26[83]},
      {stage2_26[26]}
   );
   gpc1_1 gpc2084 (
      {stage1_27[55]},
      {stage2_27[32]}
   );
   gpc1_1 gpc2085 (
      {stage1_28[46]},
      {stage2_28[25]}
   );
   gpc1_1 gpc2086 (
      {stage1_28[47]},
      {stage2_28[26]}
   );
   gpc1_1 gpc2087 (
      {stage1_29[78]},
      {stage2_29[19]}
   );
   gpc1_1 gpc2088 (
      {stage1_29[79]},
      {stage2_29[20]}
   );
   gpc1_1 gpc2089 (
      {stage1_30[47]},
      {stage2_30[27]}
   );
   gpc1_1 gpc2090 (
      {stage1_30[48]},
      {stage2_30[28]}
   );
   gpc1_1 gpc2091 (
      {stage1_30[49]},
      {stage2_30[29]}
   );
   gpc1_1 gpc2092 (
      {stage1_30[50]},
      {stage2_30[30]}
   );
   gpc1_1 gpc2093 (
      {stage1_30[51]},
      {stage2_30[31]}
   );
   gpc1_1 gpc2094 (
      {stage1_30[52]},
      {stage2_30[32]}
   );
   gpc1_1 gpc2095 (
      {stage1_30[53]},
      {stage2_30[33]}
   );
   gpc1_1 gpc2096 (
      {stage1_30[54]},
      {stage2_30[34]}
   );
   gpc1_1 gpc2097 (
      {stage1_30[55]},
      {stage2_30[35]}
   );
   gpc1_1 gpc2098 (
      {stage1_30[56]},
      {stage2_30[36]}
   );
   gpc1_1 gpc2099 (
      {stage1_30[57]},
      {stage2_30[37]}
   );
   gpc1_1 gpc2100 (
      {stage1_30[58]},
      {stage2_30[38]}
   );
   gpc1_1 gpc2101 (
      {stage1_30[59]},
      {stage2_30[39]}
   );
   gpc1_1 gpc2102 (
      {stage1_30[60]},
      {stage2_30[40]}
   );
   gpc1_1 gpc2103 (
      {stage1_30[61]},
      {stage2_30[41]}
   );
   gpc1_1 gpc2104 (
      {stage1_30[62]},
      {stage2_30[42]}
   );
   gpc1_1 gpc2105 (
      {stage1_30[63]},
      {stage2_30[43]}
   );
   gpc1_1 gpc2106 (
      {stage1_30[64]},
      {stage2_30[44]}
   );
   gpc1_1 gpc2107 (
      {stage1_30[65]},
      {stage2_30[45]}
   );
   gpc1_1 gpc2108 (
      {stage1_30[66]},
      {stage2_30[46]}
   );
   gpc1_1 gpc2109 (
      {stage1_30[67]},
      {stage2_30[47]}
   );
   gpc1_1 gpc2110 (
      {stage1_30[68]},
      {stage2_30[48]}
   );
   gpc1_1 gpc2111 (
      {stage1_30[69]},
      {stage2_30[49]}
   );
   gpc1_1 gpc2112 (
      {stage1_30[70]},
      {stage2_30[50]}
   );
   gpc1_1 gpc2113 (
      {stage1_30[71]},
      {stage2_30[51]}
   );
   gpc1_1 gpc2114 (
      {stage1_32[82]},
      {stage2_32[24]}
   );
   gpc1_1 gpc2115 (
      {stage1_33[61]},
      {stage2_33[27]}
   );
   gpc1_1 gpc2116 (
      {stage1_33[62]},
      {stage2_33[28]}
   );
   gpc1_1 gpc2117 (
      {stage1_34[66]},
      {stage2_34[30]}
   );
   gpc1_1 gpc2118 (
      {stage1_34[67]},
      {stage2_34[31]}
   );
   gpc1_1 gpc2119 (
      {stage1_35[42]},
      {stage2_35[24]}
   );
   gpc1_1 gpc2120 (
      {stage1_35[43]},
      {stage2_35[25]}
   );
   gpc1_1 gpc2121 (
      {stage1_35[44]},
      {stage2_35[26]}
   );
   gpc1_1 gpc2122 (
      {stage1_35[45]},
      {stage2_35[27]}
   );
   gpc1_1 gpc2123 (
      {stage1_35[46]},
      {stage2_35[28]}
   );
   gpc1_1 gpc2124 (
      {stage1_35[47]},
      {stage2_35[29]}
   );
   gpc1_1 gpc2125 (
      {stage1_36[48]},
      {stage2_36[20]}
   );
   gpc1_1 gpc2126 (
      {stage1_36[49]},
      {stage2_36[21]}
   );
   gpc1_1 gpc2127 (
      {stage1_36[50]},
      {stage2_36[22]}
   );
   gpc1_1 gpc2128 (
      {stage1_36[51]},
      {stage2_36[23]}
   );
   gpc1_1 gpc2129 (
      {stage1_36[52]},
      {stage2_36[24]}
   );
   gpc1_1 gpc2130 (
      {stage1_36[53]},
      {stage2_36[25]}
   );
   gpc1_1 gpc2131 (
      {stage1_36[54]},
      {stage2_36[26]}
   );
   gpc1_1 gpc2132 (
      {stage1_36[55]},
      {stage2_36[27]}
   );
   gpc1_1 gpc2133 (
      {stage1_36[56]},
      {stage2_36[28]}
   );
   gpc1_1 gpc2134 (
      {stage1_36[57]},
      {stage2_36[29]}
   );
   gpc1_1 gpc2135 (
      {stage1_36[58]},
      {stage2_36[30]}
   );
   gpc1_1 gpc2136 (
      {stage1_36[59]},
      {stage2_36[31]}
   );
   gpc1_1 gpc2137 (
      {stage1_36[60]},
      {stage2_36[32]}
   );
   gpc1_1 gpc2138 (
      {stage1_37[89]},
      {stage2_37[29]}
   );
   gpc1_1 gpc2139 (
      {stage1_37[90]},
      {stage2_37[30]}
   );
   gpc1_1 gpc2140 (
      {stage1_37[91]},
      {stage2_37[31]}
   );
   gpc1_1 gpc2141 (
      {stage1_37[92]},
      {stage2_37[32]}
   );
   gpc1_1 gpc2142 (
      {stage1_37[93]},
      {stage2_37[33]}
   );
   gpc1_1 gpc2143 (
      {stage1_37[94]},
      {stage2_37[34]}
   );
   gpc1_1 gpc2144 (
      {stage1_37[95]},
      {stage2_37[35]}
   );
   gpc1_1 gpc2145 (
      {stage1_37[96]},
      {stage2_37[36]}
   );
   gpc1_1 gpc2146 (
      {stage1_38[35]},
      {stage2_38[27]}
   );
   gpc1_1 gpc2147 (
      {stage1_38[36]},
      {stage2_38[28]}
   );
   gpc1_1 gpc2148 (
      {stage1_38[37]},
      {stage2_38[29]}
   );
   gpc1_1 gpc2149 (
      {stage1_38[38]},
      {stage2_38[30]}
   );
   gpc1_1 gpc2150 (
      {stage1_38[39]},
      {stage2_38[31]}
   );
   gpc1_1 gpc2151 (
      {stage1_38[40]},
      {stage2_38[32]}
   );
   gpc1_1 gpc2152 (
      {stage1_38[41]},
      {stage2_38[33]}
   );
   gpc1_1 gpc2153 (
      {stage1_38[42]},
      {stage2_38[34]}
   );
   gpc1_1 gpc2154 (
      {stage1_38[43]},
      {stage2_38[35]}
   );
   gpc1_1 gpc2155 (
      {stage1_39[92]},
      {stage2_39[21]}
   );
   gpc1_1 gpc2156 (
      {stage1_40[54]},
      {stage2_40[26]}
   );
   gpc1_1 gpc2157 (
      {stage1_40[55]},
      {stage2_40[27]}
   );
   gpc1_1 gpc2158 (
      {stage1_40[56]},
      {stage2_40[28]}
   );
   gpc1_1 gpc2159 (
      {stage1_40[57]},
      {stage2_40[29]}
   );
   gpc1_1 gpc2160 (
      {stage1_40[58]},
      {stage2_40[30]}
   );
   gpc1_1 gpc2161 (
      {stage1_40[59]},
      {stage2_40[31]}
   );
   gpc1_1 gpc2162 (
      {stage1_40[60]},
      {stage2_40[32]}
   );
   gpc1_1 gpc2163 (
      {stage1_40[61]},
      {stage2_40[33]}
   );
   gpc1_1 gpc2164 (
      {stage1_40[62]},
      {stage2_40[34]}
   );
   gpc1_1 gpc2165 (
      {stage1_42[50]},
      {stage2_42[17]}
   );
   gpc1_1 gpc2166 (
      {stage1_43[78]},
      {stage2_43[20]}
   );
   gpc1_1 gpc2167 (
      {stage1_45[47]},
      {stage2_45[24]}
   );
   gpc1_1 gpc2168 (
      {stage1_45[48]},
      {stage2_45[25]}
   );
   gpc1_1 gpc2169 (
      {stage1_45[49]},
      {stage2_45[26]}
   );
   gpc1_1 gpc2170 (
      {stage1_45[50]},
      {stage2_45[27]}
   );
   gpc1_1 gpc2171 (
      {stage1_45[51]},
      {stage2_45[28]}
   );
   gpc1_1 gpc2172 (
      {stage1_45[52]},
      {stage2_45[29]}
   );
   gpc1_1 gpc2173 (
      {stage1_45[53]},
      {stage2_45[30]}
   );
   gpc1_1 gpc2174 (
      {stage1_45[54]},
      {stage2_45[31]}
   );
   gpc1_1 gpc2175 (
      {stage1_45[55]},
      {stage2_45[32]}
   );
   gpc1_1 gpc2176 (
      {stage1_45[56]},
      {stage2_45[33]}
   );
   gpc1_1 gpc2177 (
      {stage1_45[57]},
      {stage2_45[34]}
   );
   gpc1_1 gpc2178 (
      {stage1_46[76]},
      {stage2_46[19]}
   );
   gpc1_1 gpc2179 (
      {stage1_46[77]},
      {stage2_46[20]}
   );
   gpc1_1 gpc2180 (
      {stage1_46[78]},
      {stage2_46[21]}
   );
   gpc1_1 gpc2181 (
      {stage1_46[79]},
      {stage2_46[22]}
   );
   gpc1_1 gpc2182 (
      {stage1_47[64]},
      {stage2_47[30]}
   );
   gpc1_1 gpc2183 (
      {stage1_47[65]},
      {stage2_47[31]}
   );
   gpc1_1 gpc2184 (
      {stage1_47[66]},
      {stage2_47[32]}
   );
   gpc1_1 gpc2185 (
      {stage1_47[67]},
      {stage2_47[33]}
   );
   gpc1_1 gpc2186 (
      {stage1_47[68]},
      {stage2_47[34]}
   );
   gpc1_1 gpc2187 (
      {stage1_47[69]},
      {stage2_47[35]}
   );
   gpc1_1 gpc2188 (
      {stage1_48[42]},
      {stage2_48[27]}
   );
   gpc1_1 gpc2189 (
      {stage1_48[43]},
      {stage2_48[28]}
   );
   gpc1_1 gpc2190 (
      {stage1_48[44]},
      {stage2_48[29]}
   );
   gpc1_1 gpc2191 (
      {stage1_48[45]},
      {stage2_48[30]}
   );
   gpc1_1 gpc2192 (
      {stage1_50[66]},
      {stage2_50[28]}
   );
   gpc1_1 gpc2193 (
      {stage1_50[67]},
      {stage2_50[29]}
   );
   gpc1_1 gpc2194 (
      {stage1_50[68]},
      {stage2_50[30]}
   );
   gpc1_1 gpc2195 (
      {stage1_50[69]},
      {stage2_50[31]}
   );
   gpc1_1 gpc2196 (
      {stage1_50[70]},
      {stage2_50[32]}
   );
   gpc1_1 gpc2197 (
      {stage1_51[42]},
      {stage2_51[25]}
   );
   gpc1_1 gpc2198 (
      {stage1_51[43]},
      {stage2_51[26]}
   );
   gpc1_1 gpc2199 (
      {stage1_51[44]},
      {stage2_51[27]}
   );
   gpc1_1 gpc2200 (
      {stage1_51[45]},
      {stage2_51[28]}
   );
   gpc1_1 gpc2201 (
      {stage1_51[46]},
      {stage2_51[29]}
   );
   gpc1_1 gpc2202 (
      {stage1_51[47]},
      {stage2_51[30]}
   );
   gpc1_1 gpc2203 (
      {stage1_52[60]},
      {stage2_52[17]}
   );
   gpc1_1 gpc2204 (
      {stage1_53[45]},
      {stage2_53[22]}
   );
   gpc1_1 gpc2205 (
      {stage1_53[46]},
      {stage2_53[23]}
   );
   gpc1_1 gpc2206 (
      {stage1_53[47]},
      {stage2_53[24]}
   );
   gpc1_1 gpc2207 (
      {stage1_53[48]},
      {stage2_53[25]}
   );
   gpc1_1 gpc2208 (
      {stage1_53[49]},
      {stage2_53[26]}
   );
   gpc1_1 gpc2209 (
      {stage1_53[50]},
      {stage2_53[27]}
   );
   gpc1_1 gpc2210 (
      {stage1_53[51]},
      {stage2_53[28]}
   );
   gpc1_1 gpc2211 (
      {stage1_53[52]},
      {stage2_53[29]}
   );
   gpc1_1 gpc2212 (
      {stage1_53[53]},
      {stage2_53[30]}
   );
   gpc1_1 gpc2213 (
      {stage1_53[54]},
      {stage2_53[31]}
   );
   gpc1_1 gpc2214 (
      {stage1_53[55]},
      {stage2_53[32]}
   );
   gpc1_1 gpc2215 (
      {stage1_53[56]},
      {stage2_53[33]}
   );
   gpc1_1 gpc2216 (
      {stage1_53[57]},
      {stage2_53[34]}
   );
   gpc1_1 gpc2217 (
      {stage1_53[58]},
      {stage2_53[35]}
   );
   gpc1_1 gpc2218 (
      {stage1_53[59]},
      {stage2_53[36]}
   );
   gpc1_1 gpc2219 (
      {stage1_53[60]},
      {stage2_53[37]}
   );
   gpc1_1 gpc2220 (
      {stage1_53[61]},
      {stage2_53[38]}
   );
   gpc1_1 gpc2221 (
      {stage1_54[51]},
      {stage2_54[28]}
   );
   gpc1_1 gpc2222 (
      {stage1_56[52]},
      {stage2_56[22]}
   );
   gpc1_1 gpc2223 (
      {stage1_56[53]},
      {stage2_56[23]}
   );
   gpc1_1 gpc2224 (
      {stage1_56[54]},
      {stage2_56[24]}
   );
   gpc1_1 gpc2225 (
      {stage1_56[55]},
      {stage2_56[25]}
   );
   gpc1_1 gpc2226 (
      {stage1_56[56]},
      {stage2_56[26]}
   );
   gpc1_1 gpc2227 (
      {stage1_57[48]},
      {stage2_57[23]}
   );
   gpc1_1 gpc2228 (
      {stage1_57[49]},
      {stage2_57[24]}
   );
   gpc1_1 gpc2229 (
      {stage1_57[50]},
      {stage2_57[25]}
   );
   gpc1_1 gpc2230 (
      {stage1_57[51]},
      {stage2_57[26]}
   );
   gpc1_1 gpc2231 (
      {stage1_57[52]},
      {stage2_57[27]}
   );
   gpc1_1 gpc2232 (
      {stage1_57[53]},
      {stage2_57[28]}
   );
   gpc1_1 gpc2233 (
      {stage1_57[54]},
      {stage2_57[29]}
   );
   gpc1_1 gpc2234 (
      {stage1_57[55]},
      {stage2_57[30]}
   );
   gpc1_1 gpc2235 (
      {stage1_57[56]},
      {stage2_57[31]}
   );
   gpc1_1 gpc2236 (
      {stage1_57[57]},
      {stage2_57[32]}
   );
   gpc1_1 gpc2237 (
      {stage1_59[42]},
      {stage2_59[21]}
   );
   gpc1_1 gpc2238 (
      {stage1_59[43]},
      {stage2_59[22]}
   );
   gpc1_1 gpc2239 (
      {stage1_59[44]},
      {stage2_59[23]}
   );
   gpc1_1 gpc2240 (
      {stage1_59[45]},
      {stage2_59[24]}
   );
   gpc1_1 gpc2241 (
      {stage1_59[46]},
      {stage2_59[25]}
   );
   gpc1_1 gpc2242 (
      {stage1_59[47]},
      {stage2_59[26]}
   );
   gpc1_1 gpc2243 (
      {stage1_59[48]},
      {stage2_59[27]}
   );
   gpc1_1 gpc2244 (
      {stage1_59[49]},
      {stage2_59[28]}
   );
   gpc1_1 gpc2245 (
      {stage1_59[50]},
      {stage2_59[29]}
   );
   gpc1_1 gpc2246 (
      {stage1_59[51]},
      {stage2_59[30]}
   );
   gpc1_1 gpc2247 (
      {stage1_59[52]},
      {stage2_59[31]}
   );
   gpc1_1 gpc2248 (
      {stage1_59[53]},
      {stage2_59[32]}
   );
   gpc1_1 gpc2249 (
      {stage1_59[54]},
      {stage2_59[33]}
   );
   gpc1_1 gpc2250 (
      {stage1_59[55]},
      {stage2_59[34]}
   );
   gpc1_1 gpc2251 (
      {stage1_60[48]},
      {stage2_60[17]}
   );
   gpc1_1 gpc2252 (
      {stage1_60[49]},
      {stage2_60[18]}
   );
   gpc1_1 gpc2253 (
      {stage1_60[50]},
      {stage2_60[19]}
   );
   gpc1_1 gpc2254 (
      {stage1_60[51]},
      {stage2_60[20]}
   );
   gpc1_1 gpc2255 (
      {stage1_60[52]},
      {stage2_60[21]}
   );
   gpc1_1 gpc2256 (
      {stage1_61[57]},
      {stage2_61[27]}
   );
   gpc1_1 gpc2257 (
      {stage1_61[58]},
      {stage2_61[28]}
   );
   gpc1_1 gpc2258 (
      {stage1_62[87]},
      {stage2_62[27]}
   );
   gpc1_1 gpc2259 (
      {stage1_62[88]},
      {stage2_62[28]}
   );
   gpc1_1 gpc2260 (
      {stage1_62[89]},
      {stage2_62[29]}
   );
   gpc1_1 gpc2261 (
      {stage1_62[90]},
      {stage2_62[30]}
   );
   gpc1_1 gpc2262 (
      {stage1_62[91]},
      {stage2_62[31]}
   );
   gpc1_1 gpc2263 (
      {stage1_62[92]},
      {stage2_62[32]}
   );
   gpc1_1 gpc2264 (
      {stage1_62[93]},
      {stage2_62[33]}
   );
   gpc1_1 gpc2265 (
      {stage1_62[94]},
      {stage2_62[34]}
   );
   gpc1_1 gpc2266 (
      {stage1_62[95]},
      {stage2_62[35]}
   );
   gpc1_1 gpc2267 (
      {stage1_62[96]},
      {stage2_62[36]}
   );
   gpc1_1 gpc2268 (
      {stage1_62[97]},
      {stage2_62[37]}
   );
   gpc1_1 gpc2269 (
      {stage1_63[36]},
      {stage2_63[21]}
   );
   gpc1_1 gpc2270 (
      {stage1_63[37]},
      {stage2_63[22]}
   );
   gpc1_1 gpc2271 (
      {stage1_63[38]},
      {stage2_63[23]}
   );
   gpc1_1 gpc2272 (
      {stage1_63[39]},
      {stage2_63[24]}
   );
   gpc1_1 gpc2273 (
      {stage1_63[40]},
      {stage2_63[25]}
   );
   gpc1_1 gpc2274 (
      {stage1_63[41]},
      {stage2_63[26]}
   );
   gpc1_1 gpc2275 (
      {stage1_63[42]},
      {stage2_63[27]}
   );
   gpc1_1 gpc2276 (
      {stage1_63[43]},
      {stage2_63[28]}
   );
   gpc1_1 gpc2277 (
      {stage1_63[44]},
      {stage2_63[29]}
   );
   gpc1_1 gpc2278 (
      {stage1_63[45]},
      {stage2_63[30]}
   );
   gpc1_1 gpc2279 (
      {stage1_63[46]},
      {stage2_63[31]}
   );
   gpc1_1 gpc2280 (
      {stage1_63[47]},
      {stage2_63[32]}
   );
   gpc1_1 gpc2281 (
      {stage1_63[48]},
      {stage2_63[33]}
   );
   gpc1_1 gpc2282 (
      {stage1_63[49]},
      {stage2_63[34]}
   );
   gpc1_1 gpc2283 (
      {stage1_63[50]},
      {stage2_63[35]}
   );
   gpc1_1 gpc2284 (
      {stage1_63[51]},
      {stage2_63[36]}
   );
   gpc1_1 gpc2285 (
      {stage1_63[52]},
      {stage2_63[37]}
   );
   gpc1_1 gpc2286 (
      {stage1_64[22]},
      {stage2_64[18]}
   );
   gpc1_1 gpc2287 (
      {stage1_64[23]},
      {stage2_64[19]}
   );
   gpc1_1 gpc2288 (
      {stage1_64[24]},
      {stage2_64[20]}
   );
   gpc1_1 gpc2289 (
      {stage1_64[25]},
      {stage2_64[21]}
   );
   gpc1_1 gpc2290 (
      {stage1_64[26]},
      {stage2_64[22]}
   );
   gpc1_1 gpc2291 (
      {stage1_64[27]},
      {stage2_64[23]}
   );
   gpc1_1 gpc2292 (
      {stage1_64[28]},
      {stage2_64[24]}
   );
   gpc1_1 gpc2293 (
      {stage1_64[29]},
      {stage2_64[25]}
   );
   gpc606_5 gpc2294 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc2295 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc2296 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc2297 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4]},
      {stage2_2[18]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc615_5 gpc2298 (
      {stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9]},
      {stage2_2[19]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc2299 (
      {stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24], 1'b0},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[2],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc606_5 gpc2300 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[3],stage3_4[6]}
   );
   gpc606_5 gpc2301 (
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[4],stage3_4[7]}
   );
   gpc615_5 gpc2302 (
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_5[0]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[5],stage3_4[8]}
   );
   gpc606_5 gpc2303 (
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[6]}
   );
   gpc606_5 gpc2304 (
      {stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[4],stage3_7[4],stage3_6[5],stage3_5[7]}
   );
   gpc615_5 gpc2305 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[12]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[5],stage3_7[5],stage3_6[6]}
   );
   gpc606_5 gpc2306 (
      {stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[3],stage3_8[6],stage3_7[6]}
   );
   gpc606_5 gpc2307 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[4],stage3_8[7],stage3_7[7]}
   );
   gpc606_5 gpc2308 (
      {stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[5],stage3_8[8],stage3_7[8]}
   );
   gpc606_5 gpc2309 (
      {stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[6],stage3_8[9],stage3_7[9]}
   );
   gpc615_5 gpc2310 (
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10]},
      {stage2_9[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc2311 (
      {stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_9[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[8],stage3_8[11]}
   );
   gpc615_5 gpc2312 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20]},
      {stage2_9[26]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[9],stage3_8[12]}
   );
   gpc615_5 gpc2313 (
      {stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_9[27]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[10],stage3_8[13]}
   );
   gpc615_5 gpc2314 (
      {stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_9[28]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[11],stage3_8[14]}
   );
   gpc606_5 gpc2315 (
      {stage2_9[29], stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[12]}
   );
   gpc2116_5 gpc2316 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage2_14[0], stage2_14[1]},
      {stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[6],stage3_11[10]}
   );
   gpc615_5 gpc2317 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[1],stage3_14[1],stage3_13[2],stage3_12[7],stage3_11[11]}
   );
   gpc615_5 gpc2318 (
      {stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage2_12[2]},
      {stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11], stage2_13[12]},
      {stage3_15[2],stage3_14[2],stage3_13[3],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc2319 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[4],stage3_12[9]}
   );
   gpc606_5 gpc2320 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11], stage2_14[12], stage2_14[13]},
      {stage3_16[1],stage3_15[4],stage3_14[4],stage3_13[5],stage3_12[10]}
   );
   gpc606_5 gpc2321 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19]},
      {stage3_16[2],stage3_15[5],stage3_14[5],stage3_13[6],stage3_12[11]}
   );
   gpc606_5 gpc2322 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage3_16[3],stage3_15[6],stage3_14[6],stage3_13[7],stage3_12[12]}
   );
   gpc606_5 gpc2323 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30], stage2_14[31]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[4],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc2324 (
      {stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35], stage2_14[36]},
      {stage2_15[0]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[5],stage3_15[8],stage3_14[8]}
   );
   gpc615_5 gpc2325 (
      {stage2_14[37], stage2_14[38], 1'b0, 1'b0, 1'b0},
      {stage2_15[1]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[6],stage3_15[9],stage3_14[9]}
   );
   gpc2135_5 gpc2326 (
      {stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_16[18], stage2_16[19], stage2_16[20]},
      {stage2_17[0]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[3],stage3_17[3],stage3_16[7],stage3_15[10]}
   );
   gpc606_5 gpc2327 (
      {stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[1],stage3_18[4],stage3_17[4],stage3_16[8],stage3_15[11]}
   );
   gpc615_5 gpc2328 (
      {stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage2_16[21]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[2],stage3_18[5],stage3_17[5],stage3_16[9],stage3_15[12]}
   );
   gpc1163_5 gpc2329 (
      {stage2_17[13], stage2_17[14], stage2_17[15]},
      {stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6], stage2_18[7]},
      {stage2_19[0]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[3],stage3_18[6],stage3_17[6]}
   );
   gpc1163_5 gpc2330 (
      {stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13]},
      {stage2_19[1]},
      {stage2_20[1]},
      {stage3_21[1],stage3_20[1],stage3_19[4],stage3_18[7],stage3_17[7]}
   );
   gpc1163_5 gpc2331 (
      {stage2_17[19], stage2_17[20], stage2_17[21]},
      {stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[2]},
      {stage2_20[2]},
      {stage3_21[2],stage3_20[2],stage3_19[5],stage3_18[8],stage3_17[8]}
   );
   gpc606_5 gpc2332 (
      {stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27]},
      {stage2_19[3], stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage3_21[3],stage3_20[3],stage3_19[6],stage3_18[9],stage3_17[9]}
   );
   gpc615_5 gpc2333 (
      {stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31], stage2_17[32]},
      {stage2_18[20]},
      {stage2_19[9], stage2_19[10], stage2_19[11], stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage3_21[4],stage3_20[4],stage3_19[7],stage3_18[10],stage3_17[10]}
   );
   gpc2135_5 gpc2334 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[3]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[5],stage3_20[5],stage3_19[8],stage3_18[11]}
   );
   gpc2135_5 gpc2335 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[4]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[6],stage3_20[6],stage3_19[9],stage3_18[12]}
   );
   gpc1343_5 gpc2336 (
      {stage2_20[5], stage2_20[6], stage2_20[7]},
      {stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7]},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[7],stage3_20[7]}
   );
   gpc1343_5 gpc2337 (
      {stage2_20[8], stage2_20[9], stage2_20[10]},
      {stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage2_23[1]},
      {stage3_24[1],stage3_23[1],stage3_22[3],stage3_21[8],stage3_20[8]}
   );
   gpc615_5 gpc2338 (
      {stage2_20[11], stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15]},
      {stage2_21[12]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[2],stage3_23[2],stage3_22[4],stage3_21[9],stage3_20[9]}
   );
   gpc615_5 gpc2339 (
      {stage2_20[16], stage2_20[17], stage2_20[18], stage2_20[19], stage2_20[20]},
      {stage2_21[13]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[3],stage3_23[3],stage3_22[5],stage3_21[10],stage3_20[10]}
   );
   gpc615_5 gpc2340 (
      {stage2_20[21], stage2_20[22], stage2_20[23], stage2_20[24], stage2_20[25]},
      {stage2_21[14]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[4],stage3_23[4],stage3_22[6],stage3_21[11],stage3_20[11]}
   );
   gpc615_5 gpc2341 (
      {stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30]},
      {stage2_21[15]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[5],stage3_23[5],stage3_22[7],stage3_21[12],stage3_20[12]}
   );
   gpc623_5 gpc2342 (
      {stage2_20[31], stage2_20[32], stage2_20[33]},
      {stage2_21[16], stage2_21[17]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], 1'b0},
      {stage3_24[6],stage3_23[6],stage3_22[8],stage3_21[13],stage3_20[13]}
   );
   gpc2135_5 gpc2343 (
      {stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5], stage2_23[6]},
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[7],stage3_23[7]}
   );
   gpc2135_5 gpc2344 (
      {stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage2_25[1]},
      {stage2_26[2], stage2_26[3]},
      {stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[8],stage3_23[8]}
   );
   gpc615_5 gpc2345 (
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16]},
      {stage2_24[6]},
      {stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7]},
      {stage3_27[2],stage3_26[2],stage3_25[2],stage3_24[9],stage3_23[9]}
   );
   gpc615_5 gpc2346 (
      {stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_24[7]},
      {stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], stage2_25[13]},
      {stage3_27[3],stage3_26[3],stage3_25[3],stage3_24[10],stage3_23[10]}
   );
   gpc615_5 gpc2347 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage2_24[8]},
      {stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18], stage2_25[19]},
      {stage3_27[4],stage3_26[4],stage3_25[4],stage3_24[11],stage3_23[11]}
   );
   gpc606_5 gpc2348 (
      {stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13], stage2_24[14]},
      {stage2_26[4], stage2_26[5], stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9]},
      {stage3_28[0],stage3_27[5],stage3_26[5],stage3_25[5],stage3_24[12]}
   );
   gpc606_5 gpc2349 (
      {stage2_24[15], stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20]},
      {stage2_26[10], stage2_26[11], stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15]},
      {stage3_28[1],stage3_27[6],stage3_26[6],stage3_25[6],stage3_24[13]}
   );
   gpc606_5 gpc2350 (
      {stage2_24[21], stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26]},
      {stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21]},
      {stage3_28[2],stage3_27[7],stage3_26[7],stage3_25[7],stage3_24[14]}
   );
   gpc2135_5 gpc2351 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4]},
      {stage2_28[0], stage2_28[1], stage2_28[2]},
      {stage2_29[0]},
      {stage2_30[0], stage2_30[1]},
      {stage3_31[0],stage3_30[0],stage3_29[0],stage3_28[3],stage3_27[8]}
   );
   gpc2135_5 gpc2352 (
      {stage2_27[5], stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9]},
      {stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage2_29[1]},
      {stage2_30[2], stage2_30[3]},
      {stage3_31[1],stage3_30[1],stage3_29[1],stage3_28[4],stage3_27[9]}
   );
   gpc2135_5 gpc2353 (
      {stage2_27[10], stage2_27[11], stage2_27[12], stage2_27[13], stage2_27[14]},
      {stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[2]},
      {stage2_30[4], stage2_30[5]},
      {stage3_31[2],stage3_30[2],stage3_29[2],stage3_28[5],stage3_27[10]}
   );
   gpc606_5 gpc2354 (
      {stage2_27[15], stage2_27[16], stage2_27[17], stage2_27[18], stage2_27[19], stage2_27[20]},
      {stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6], stage2_29[7], stage2_29[8]},
      {stage3_31[3],stage3_30[3],stage3_29[3],stage3_28[6],stage3_27[11]}
   );
   gpc606_5 gpc2355 (
      {stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26]},
      {stage2_29[9], stage2_29[10], stage2_29[11], stage2_29[12], stage2_29[13], stage2_29[14]},
      {stage3_31[4],stage3_30[4],stage3_29[4],stage3_28[7],stage3_27[12]}
   );
   gpc606_5 gpc2356 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_29[15], stage2_29[16], stage2_29[17], stage2_29[18], stage2_29[19], stage2_29[20]},
      {stage3_31[5],stage3_30[5],stage3_29[5],stage3_28[8],stage3_27[13]}
   );
   gpc606_5 gpc2357 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[0],stage3_31[6],stage3_30[6],stage3_29[6],stage3_28[9]}
   );
   gpc606_5 gpc2358 (
      {stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19], stage2_28[20]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[1],stage3_31[7],stage3_30[7],stage3_29[7],stage3_28[10]}
   );
   gpc2135_5 gpc2359 (
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22]},
      {stage2_31[0], stage2_31[1], stage2_31[2]},
      {stage2_32[0]},
      {stage2_33[0], stage2_33[1]},
      {stage3_34[0],stage3_33[0],stage3_32[2],stage3_31[8],stage3_30[8]}
   );
   gpc2135_5 gpc2360 (
      {stage2_30[23], stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27]},
      {stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_32[1]},
      {stage2_33[2], stage2_33[3]},
      {stage3_34[1],stage3_33[1],stage3_32[3],stage3_31[9],stage3_30[9]}
   );
   gpc2135_5 gpc2361 (
      {stage2_30[28], stage2_30[29], stage2_30[30], stage2_30[31], stage2_30[32]},
      {stage2_31[6], stage2_31[7], stage2_31[8]},
      {stage2_32[2]},
      {stage2_33[4], stage2_33[5]},
      {stage3_34[2],stage3_33[2],stage3_32[4],stage3_31[10],stage3_30[10]}
   );
   gpc2135_5 gpc2362 (
      {stage2_30[33], stage2_30[34], stage2_30[35], stage2_30[36], stage2_30[37]},
      {stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage2_32[3]},
      {stage2_33[6], stage2_33[7]},
      {stage3_34[3],stage3_33[3],stage3_32[5],stage3_31[11],stage3_30[11]}
   );
   gpc2135_5 gpc2363 (
      {stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41], stage2_30[42]},
      {stage2_31[12], stage2_31[13], stage2_31[14]},
      {stage2_32[4]},
      {stage2_33[8], stage2_33[9]},
      {stage3_34[4],stage3_33[4],stage3_32[6],stage3_31[12],stage3_30[12]}
   );
   gpc615_5 gpc2364 (
      {stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage2_31[15]},
      {stage2_32[5], stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10]},
      {stage3_34[5],stage3_33[5],stage3_32[7],stage3_31[13],stage3_30[13]}
   );
   gpc615_5 gpc2365 (
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], 1'b0},
      {stage2_31[16]},
      {stage2_32[11], stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16]},
      {stage3_34[6],stage3_33[6],stage3_32[8],stage3_31[14],stage3_30[14]}
   );
   gpc117_4 gpc2366 (
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_32[17]},
      {stage2_33[10]},
      {stage3_34[7],stage3_33[7],stage3_32[9],stage3_31[15]}
   );
   gpc606_5 gpc2367 (
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[0],stage3_34[8],stage3_33[8],stage3_32[10]}
   );
   gpc606_5 gpc2368 (
      {stage2_33[11], stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[1],stage3_34[9],stage3_33[9]}
   );
   gpc606_5 gpc2369 (
      {stage2_33[17], stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[2],stage3_35[2],stage3_34[10],stage3_33[10]}
   );
   gpc606_5 gpc2370 (
      {stage2_33[23], stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28]},
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage3_37[2],stage3_36[3],stage3_35[3],stage3_34[11],stage3_33[11]}
   );
   gpc135_4 gpc2371 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10]},
      {stage2_35[18], stage2_35[19], stage2_35[20]},
      {stage2_36[0]},
      {stage3_37[3],stage3_36[4],stage3_35[4],stage3_34[12]}
   );
   gpc135_4 gpc2372 (
      {stage2_34[11], stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15]},
      {stage2_35[21], stage2_35[22], stage2_35[23]},
      {stage2_36[1]},
      {stage3_37[4],stage3_36[5],stage3_35[5],stage3_34[13]}
   );
   gpc135_4 gpc2373 (
      {stage2_34[16], stage2_34[17], stage2_34[18], stage2_34[19], stage2_34[20]},
      {stage2_35[24], stage2_35[25], stage2_35[26]},
      {stage2_36[2]},
      {stage3_37[5],stage3_36[6],stage3_35[6],stage3_34[14]}
   );
   gpc615_5 gpc2374 (
      {stage2_34[21], stage2_34[22], stage2_34[23], stage2_34[24], stage2_34[25]},
      {stage2_35[27]},
      {stage2_36[3], stage2_36[4], stage2_36[5], stage2_36[6], stage2_36[7], stage2_36[8]},
      {stage3_38[0],stage3_37[6],stage3_36[7],stage3_35[7],stage3_34[15]}
   );
   gpc615_5 gpc2375 (
      {stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29], stage2_34[30]},
      {stage2_35[28]},
      {stage2_36[9], stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14]},
      {stage3_38[1],stage3_37[7],stage3_36[8],stage3_35[8],stage3_34[16]}
   );
   gpc1163_5 gpc2376 (
      {stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage2_38[0]},
      {stage2_39[0]},
      {stage3_40[0],stage3_39[0],stage3_38[2],stage3_37[8],stage3_36[9]}
   );
   gpc1163_5 gpc2377 (
      {stage2_36[18], stage2_36[19], stage2_36[20]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_38[1]},
      {stage2_39[1]},
      {stage3_40[1],stage3_39[1],stage3_38[3],stage3_37[9],stage3_36[10]}
   );
   gpc1163_5 gpc2378 (
      {stage2_36[21], stage2_36[22], stage2_36[23]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_38[2]},
      {stage2_39[2]},
      {stage3_40[2],stage3_39[2],stage3_38[4],stage3_37[10],stage3_36[11]}
   );
   gpc1163_5 gpc2379 (
      {stage2_36[24], stage2_36[25], stage2_36[26]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage2_38[3]},
      {stage2_39[3]},
      {stage3_40[3],stage3_39[3],stage3_38[5],stage3_37[11],stage3_36[12]}
   );
   gpc1163_5 gpc2380 (
      {stage2_36[27], stage2_36[28], stage2_36[29]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage2_38[4]},
      {stage2_39[4]},
      {stage3_40[4],stage3_39[4],stage3_38[6],stage3_37[12],stage3_36[13]}
   );
   gpc1163_5 gpc2381 (
      {stage2_36[30], stage2_36[31], stage2_36[32]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage2_38[5]},
      {stage2_39[5]},
      {stage3_40[5],stage3_39[5],stage3_38[7],stage3_37[13],stage3_36[14]}
   );
   gpc606_5 gpc2382 (
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[6],stage3_39[6],stage3_38[8]}
   );
   gpc606_5 gpc2383 (
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[1],stage3_40[7],stage3_39[7],stage3_38[9]}
   );
   gpc606_5 gpc2384 (
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[2],stage3_40[8],stage3_39[8],stage3_38[10]}
   );
   gpc606_5 gpc2385 (
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[3],stage3_40[9],stage3_39[9],stage3_38[11]}
   );
   gpc606_5 gpc2386 (
      {stage2_38[30], stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[4],stage3_40[10],stage3_39[10],stage3_38[12]}
   );
   gpc606_5 gpc2387 (
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[5],stage3_41[5],stage3_40[11],stage3_39[11]}
   );
   gpc606_5 gpc2388 (
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[6],stage3_41[6],stage3_40[12],stage3_39[12]}
   );
   gpc615_5 gpc2389 (
      {stage2_39[18], stage2_39[19], stage2_39[20], stage2_39[21], 1'b0},
      {stage2_40[30]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[7],stage3_41[7],stage3_40[13],stage3_39[13]}
   );
   gpc606_5 gpc2390 (
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[0],stage3_43[3],stage3_42[8],stage3_41[8]}
   );
   gpc606_5 gpc2391 (
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11]},
      {stage3_45[1],stage3_44[1],stage3_43[4],stage3_42[9],stage3_41[9]}
   );
   gpc615_5 gpc2392 (
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4]},
      {stage2_43[12]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[2],stage3_44[2],stage3_43[5],stage3_42[10]}
   );
   gpc615_5 gpc2393 (
      {stage2_42[5], stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9]},
      {stage2_43[13]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[3],stage3_44[3],stage3_43[6],stage3_42[11]}
   );
   gpc615_5 gpc2394 (
      {stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17], stage2_43[18]},
      {stage2_44[12]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[2],stage3_45[4],stage3_44[4],stage3_43[7]}
   );
   gpc606_5 gpc2395 (
      {stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17], stage2_44[18]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[1],stage3_46[3],stage3_45[5],stage3_44[5]}
   );
   gpc606_5 gpc2396 (
      {stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23], stage2_44[24]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[2],stage3_46[4],stage3_45[6],stage3_44[6]}
   );
   gpc615_5 gpc2397 (
      {stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage2_45[6]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[3],stage3_46[5],stage3_45[7],stage3_44[7]}
   );
   gpc606_5 gpc2398 (
      {stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11], stage2_45[12]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[3],stage3_47[4],stage3_46[6],stage3_45[8]}
   );
   gpc615_5 gpc2399 (
      {stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage2_46[18]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[4],stage3_47[5],stage3_46[7],stage3_45[9]}
   );
   gpc615_5 gpc2400 (
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22]},
      {stage2_46[19]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[5],stage3_47[6],stage3_46[8],stage3_45[10]}
   );
   gpc615_5 gpc2401 (
      {stage2_45[23], stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27]},
      {stage2_46[20]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[6],stage3_47[7],stage3_46[9],stage3_45[11]}
   );
   gpc615_5 gpc2402 (
      {stage2_45[28], stage2_45[29], stage2_45[30], stage2_45[31], stage2_45[32]},
      {stage2_46[21]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[7],stage3_47[8],stage3_46[10],stage3_45[12]}
   );
   gpc615_5 gpc2403 (
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34]},
      {stage2_48[0]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[0],stage3_49[5],stage3_48[8],stage3_47[9]}
   );
   gpc615_5 gpc2404 (
      {stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage2_49[6]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[1],stage3_50[1],stage3_49[6],stage3_48[9]}
   );
   gpc615_5 gpc2405 (
      {stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_49[7]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[2],stage3_50[2],stage3_49[7],stage3_48[10]}
   );
   gpc615_5 gpc2406 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15]},
      {stage2_49[8]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[3],stage3_50[3],stage3_49[8],stage3_48[11]}
   );
   gpc615_5 gpc2407 (
      {stage2_48[16], stage2_48[17], stage2_48[18], stage2_48[19], stage2_48[20]},
      {stage2_49[9]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[4],stage3_50[4],stage3_49[9],stage3_48[12]}
   );
   gpc615_5 gpc2408 (
      {stage2_48[21], stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25]},
      {stage2_49[10]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[5],stage3_50[5],stage3_49[10],stage3_48[13]}
   );
   gpc135_4 gpc2409 (
      {stage2_49[11], stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15]},
      {stage2_50[30], stage2_50[31], stage2_50[32]},
      {stage2_51[0]},
      {stage3_52[5],stage3_51[6],stage3_50[6],stage3_49[11]}
   );
   gpc615_5 gpc2410 (
      {stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[0],stage3_52[6],stage3_51[7]}
   );
   gpc615_5 gpc2411 (
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10]},
      {stage2_52[1]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[1],stage3_53[1],stage3_52[7],stage3_51[8]}
   );
   gpc615_5 gpc2412 (
      {stage2_51[11], stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15]},
      {stage2_52[2]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[2],stage3_53[2],stage3_52[8],stage3_51[9]}
   );
   gpc615_5 gpc2413 (
      {stage2_51[16], stage2_51[17], stage2_51[18], stage2_51[19], stage2_51[20]},
      {stage2_52[3]},
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage3_55[3],stage3_54[3],stage3_53[3],stage3_52[9],stage3_51[10]}
   );
   gpc615_5 gpc2414 (
      {stage2_51[21], stage2_51[22], stage2_51[23], stage2_51[24], stage2_51[25]},
      {stage2_52[4]},
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage3_55[4],stage3_54[4],stage3_53[4],stage3_52[10],stage3_51[11]}
   );
   gpc615_5 gpc2415 (
      {stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29], stage2_51[30]},
      {stage2_52[5]},
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage3_55[5],stage3_54[5],stage3_53[5],stage3_52[11],stage3_51[12]}
   );
   gpc615_5 gpc2416 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10]},
      {stage2_53[36]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[6],stage3_54[6],stage3_53[6],stage3_52[12]}
   );
   gpc1163_5 gpc2417 (
      {stage2_54[6], stage2_54[7], stage2_54[8]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage2_56[0]},
      {stage2_57[0]},
      {stage3_58[0],stage3_57[0],stage3_56[1],stage3_55[7],stage3_54[7]}
   );
   gpc1163_5 gpc2418 (
      {stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage2_56[1]},
      {stage2_57[1]},
      {stage3_58[1],stage3_57[1],stage3_56[2],stage3_55[8],stage3_54[8]}
   );
   gpc1163_5 gpc2419 (
      {stage2_54[12], stage2_54[13], stage2_54[14]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage2_56[2]},
      {stage2_57[2]},
      {stage3_58[2],stage3_57[2],stage3_56[3],stage3_55[9],stage3_54[9]}
   );
   gpc606_5 gpc2420 (
      {stage2_56[3], stage2_56[4], stage2_56[5], stage2_56[6], stage2_56[7], stage2_56[8]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[3],stage3_57[3],stage3_56[4]}
   );
   gpc606_5 gpc2421 (
      {stage2_56[9], stage2_56[10], stage2_56[11], stage2_56[12], stage2_56[13], stage2_56[14]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[4],stage3_57[4],stage3_56[5]}
   );
   gpc606_5 gpc2422 (
      {stage2_56[15], stage2_56[16], stage2_56[17], stage2_56[18], stage2_56[19], stage2_56[20]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[2],stage3_58[5],stage3_57[5],stage3_56[6]}
   );
   gpc606_5 gpc2423 (
      {stage2_56[21], stage2_56[22], stage2_56[23], stage2_56[24], stage2_56[25], stage2_56[26]},
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage3_60[3],stage3_59[3],stage3_58[6],stage3_57[6],stage3_56[7]}
   );
   gpc606_5 gpc2424 (
      {stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[4],stage3_59[4],stage3_58[7],stage3_57[7]}
   );
   gpc606_5 gpc2425 (
      {stage2_57[9], stage2_57[10], stage2_57[11], stage2_57[12], stage2_57[13], stage2_57[14]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[5],stage3_59[5],stage3_58[8],stage3_57[8]}
   );
   gpc606_5 gpc2426 (
      {stage2_57[15], stage2_57[16], stage2_57[17], stage2_57[18], stage2_57[19], stage2_57[20]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[6],stage3_59[6],stage3_58[9],stage3_57[9]}
   );
   gpc606_5 gpc2427 (
      {stage2_57[21], stage2_57[22], stage2_57[23], stage2_57[24], stage2_57[25], stage2_57[26]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[7],stage3_59[7],stage3_58[10],stage3_57[10]}
   );
   gpc606_5 gpc2428 (
      {stage2_57[27], stage2_57[28], stage2_57[29], stage2_57[30], stage2_57[31], stage2_57[32]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[8],stage3_59[8],stage3_58[11],stage3_57[11]}
   );
   gpc606_5 gpc2429 (
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[0],stage3_62[0],stage3_61[5],stage3_60[9]}
   );
   gpc606_5 gpc2430 (
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[1],stage3_62[1],stage3_61[6],stage3_60[10]}
   );
   gpc606_5 gpc2431 (
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[2],stage3_62[2],stage3_61[7],stage3_60[11]}
   );
   gpc623_5 gpc2432 (
      {stage2_60[18], stage2_60[19], stage2_60[20]},
      {stage2_61[0], stage2_61[1]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[3],stage3_62[3],stage3_61[8],stage3_60[12]}
   );
   gpc606_5 gpc2433 (
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6], stage2_61[7]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[4],stage3_63[4],stage3_62[4],stage3_61[9]}
   );
   gpc606_5 gpc2434 (
      {stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12], stage2_61[13]},
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage3_65[1],stage3_64[5],stage3_63[5],stage3_62[5],stage3_61[10]}
   );
   gpc606_5 gpc2435 (
      {stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17], stage2_61[18], stage2_61[19]},
      {stage2_63[12], stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17]},
      {stage3_65[2],stage3_64[6],stage3_63[6],stage3_62[6],stage3_61[11]}
   );
   gpc606_5 gpc2436 (
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[3],stage3_64[7],stage3_63[7],stage3_62[7]}
   );
   gpc1343_5 gpc2437 (
      {stage2_63[18], stage2_63[19], stage2_63[20]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9]},
      {stage2_65[0], stage2_65[1], stage2_65[2]},
      {stage2_66[0]},
      {stage3_67[0],stage3_66[1],stage3_65[4],stage3_64[8],stage3_63[8]}
   );
   gpc1343_5 gpc2438 (
      {stage2_63[21], stage2_63[22], stage2_63[23]},
      {stage2_64[10], stage2_64[11], stage2_64[12], stage2_64[13]},
      {stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage2_66[1]},
      {stage3_67[1],stage3_66[2],stage3_65[5],stage3_64[9],stage3_63[9]}
   );
   gpc1343_5 gpc2439 (
      {stage2_63[24], stage2_63[25], stage2_63[26]},
      {stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage2_66[2]},
      {stage3_67[2],stage3_66[3],stage3_65[6],stage3_64[10],stage3_63[10]}
   );
   gpc1343_5 gpc2440 (
      {stage2_63[27], stage2_63[28], stage2_63[29]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21]},
      {stage2_65[9], stage2_65[10], stage2_65[11]},
      {stage2_66[3]},
      {stage3_67[3],stage3_66[4],stage3_65[7],stage3_64[11],stage3_63[11]}
   );
   gpc1343_5 gpc2441 (
      {stage2_63[30], stage2_63[31], stage2_63[32]},
      {stage2_64[22], stage2_64[23], stage2_64[24], stage2_64[25]},
      {stage2_65[12], stage2_65[13], stage2_65[14]},
      {stage2_66[4]},
      {stage3_67[4],stage3_66[5],stage3_65[8],stage3_64[12],stage3_63[12]}
   );
   gpc1_1 gpc2442 (
      {stage2_0[18]},
      {stage3_0[3]}
   );
   gpc1_1 gpc2443 (
      {stage2_0[19]},
      {stage3_0[4]}
   );
   gpc1_1 gpc2444 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc2445 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc2446 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc2447 (
      {stage2_3[12]},
      {stage3_3[6]}
   );
   gpc1_1 gpc2448 (
      {stage2_3[13]},
      {stage3_3[7]}
   );
   gpc1_1 gpc2449 (
      {stage2_3[14]},
      {stage3_3[8]}
   );
   gpc1_1 gpc2450 (
      {stage2_3[15]},
      {stage3_3[9]}
   );
   gpc1_1 gpc2451 (
      {stage2_3[16]},
      {stage3_3[10]}
   );
   gpc1_1 gpc2452 (
      {stage2_3[17]},
      {stage3_3[11]}
   );
   gpc1_1 gpc2453 (
      {stage2_3[18]},
      {stage3_3[12]}
   );
   gpc1_1 gpc2454 (
      {stage2_3[19]},
      {stage3_3[13]}
   );
   gpc1_1 gpc2455 (
      {stage2_3[20]},
      {stage3_3[14]}
   );
   gpc1_1 gpc2456 (
      {stage2_3[21]},
      {stage3_3[15]}
   );
   gpc1_1 gpc2457 (
      {stage2_3[22]},
      {stage3_3[16]}
   );
   gpc1_1 gpc2458 (
      {stage2_3[23]},
      {stage3_3[17]}
   );
   gpc1_1 gpc2459 (
      {stage2_3[24]},
      {stage3_3[18]}
   );
   gpc1_1 gpc2460 (
      {stage2_3[25]},
      {stage3_3[19]}
   );
   gpc1_1 gpc2461 (
      {stage2_3[26]},
      {stage3_3[20]}
   );
   gpc1_1 gpc2462 (
      {stage2_3[27]},
      {stage3_3[21]}
   );
   gpc1_1 gpc2463 (
      {stage2_4[23]},
      {stage3_4[9]}
   );
   gpc1_1 gpc2464 (
      {stage2_4[24]},
      {stage3_4[10]}
   );
   gpc1_1 gpc2465 (
      {stage2_4[25]},
      {stage3_4[11]}
   );
   gpc1_1 gpc2466 (
      {stage2_5[13]},
      {stage3_5[8]}
   );
   gpc1_1 gpc2467 (
      {stage2_5[14]},
      {stage3_5[9]}
   );
   gpc1_1 gpc2468 (
      {stage2_5[15]},
      {stage3_5[10]}
   );
   gpc1_1 gpc2469 (
      {stage2_5[16]},
      {stage3_5[11]}
   );
   gpc1_1 gpc2470 (
      {stage2_5[17]},
      {stage3_5[12]}
   );
   gpc1_1 gpc2471 (
      {stage2_5[18]},
      {stage3_5[13]}
   );
   gpc1_1 gpc2472 (
      {stage2_5[19]},
      {stage3_5[14]}
   );
   gpc1_1 gpc2473 (
      {stage2_5[20]},
      {stage3_5[15]}
   );
   gpc1_1 gpc2474 (
      {stage2_5[21]},
      {stage3_5[16]}
   );
   gpc1_1 gpc2475 (
      {stage2_5[22]},
      {stage3_5[17]}
   );
   gpc1_1 gpc2476 (
      {stage2_5[23]},
      {stage3_5[18]}
   );
   gpc1_1 gpc2477 (
      {stage2_5[24]},
      {stage3_5[19]}
   );
   gpc1_1 gpc2478 (
      {stage2_5[25]},
      {stage3_5[20]}
   );
   gpc1_1 gpc2479 (
      {stage2_5[26]},
      {stage3_5[21]}
   );
   gpc1_1 gpc2480 (
      {stage2_5[27]},
      {stage3_5[22]}
   );
   gpc1_1 gpc2481 (
      {stage2_5[28]},
      {stage3_5[23]}
   );
   gpc1_1 gpc2482 (
      {stage2_6[23]},
      {stage3_6[7]}
   );
   gpc1_1 gpc2483 (
      {stage2_6[24]},
      {stage3_6[8]}
   );
   gpc1_1 gpc2484 (
      {stage2_6[25]},
      {stage3_6[9]}
   );
   gpc1_1 gpc2485 (
      {stage2_7[37]},
      {stage3_7[10]}
   );
   gpc1_1 gpc2486 (
      {stage2_7[38]},
      {stage3_7[11]}
   );
   gpc1_1 gpc2487 (
      {stage2_8[31]},
      {stage3_8[15]}
   );
   gpc1_1 gpc2488 (
      {stage2_9[35]},
      {stage3_9[13]}
   );
   gpc1_1 gpc2489 (
      {stage2_9[36]},
      {stage3_9[14]}
   );
   gpc1_1 gpc2490 (
      {stage2_9[37]},
      {stage3_9[15]}
   );
   gpc1_1 gpc2491 (
      {stage2_9[38]},
      {stage3_9[16]}
   );
   gpc1_1 gpc2492 (
      {stage2_9[39]},
      {stage3_9[17]}
   );
   gpc1_1 gpc2493 (
      {stage2_9[40]},
      {stage3_9[18]}
   );
   gpc1_1 gpc2494 (
      {stage2_9[41]},
      {stage3_9[19]}
   );
   gpc1_1 gpc2495 (
      {stage2_10[30]},
      {stage3_10[11]}
   );
   gpc1_1 gpc2496 (
      {stage2_12[27]},
      {stage3_12[13]}
   );
   gpc1_1 gpc2497 (
      {stage2_13[13]},
      {stage3_13[8]}
   );
   gpc1_1 gpc2498 (
      {stage2_13[14]},
      {stage3_13[9]}
   );
   gpc1_1 gpc2499 (
      {stage2_13[15]},
      {stage3_13[10]}
   );
   gpc1_1 gpc2500 (
      {stage2_13[16]},
      {stage3_13[11]}
   );
   gpc1_1 gpc2501 (
      {stage2_15[18]},
      {stage3_15[13]}
   );
   gpc1_1 gpc2502 (
      {stage2_15[19]},
      {stage3_15[14]}
   );
   gpc1_1 gpc2503 (
      {stage2_15[20]},
      {stage3_15[15]}
   );
   gpc1_1 gpc2504 (
      {stage2_15[21]},
      {stage3_15[16]}
   );
   gpc1_1 gpc2505 (
      {stage2_15[22]},
      {stage3_15[17]}
   );
   gpc1_1 gpc2506 (
      {stage2_15[23]},
      {stage3_15[18]}
   );
   gpc1_1 gpc2507 (
      {stage2_15[24]},
      {stage3_15[19]}
   );
   gpc1_1 gpc2508 (
      {stage2_15[25]},
      {stage3_15[20]}
   );
   gpc1_1 gpc2509 (
      {stage2_15[26]},
      {stage3_15[21]}
   );
   gpc1_1 gpc2510 (
      {stage2_15[27]},
      {stage3_15[22]}
   );
   gpc1_1 gpc2511 (
      {stage2_15[28]},
      {stage3_15[23]}
   );
   gpc1_1 gpc2512 (
      {stage2_15[29]},
      {stage3_15[24]}
   );
   gpc1_1 gpc2513 (
      {stage2_15[30]},
      {stage3_15[25]}
   );
   gpc1_1 gpc2514 (
      {stage2_16[22]},
      {stage3_16[10]}
   );
   gpc1_1 gpc2515 (
      {stage2_16[23]},
      {stage3_16[11]}
   );
   gpc1_1 gpc2516 (
      {stage2_17[33]},
      {stage3_17[11]}
   );
   gpc1_1 gpc2517 (
      {stage2_19[21]},
      {stage3_19[10]}
   );
   gpc1_1 gpc2518 (
      {stage2_19[22]},
      {stage3_19[11]}
   );
   gpc1_1 gpc2519 (
      {stage2_19[23]},
      {stage3_19[12]}
   );
   gpc1_1 gpc2520 (
      {stage2_19[24]},
      {stage3_19[13]}
   );
   gpc1_1 gpc2521 (
      {stage2_19[25]},
      {stage3_19[14]}
   );
   gpc1_1 gpc2522 (
      {stage2_19[26]},
      {stage3_19[15]}
   );
   gpc1_1 gpc2523 (
      {stage2_21[18]},
      {stage3_21[14]}
   );
   gpc1_1 gpc2524 (
      {stage2_21[19]},
      {stage3_21[15]}
   );
   gpc1_1 gpc2525 (
      {stage2_21[20]},
      {stage3_21[16]}
   );
   gpc1_1 gpc2526 (
      {stage2_21[21]},
      {stage3_21[17]}
   );
   gpc1_1 gpc2527 (
      {stage2_23[27]},
      {stage3_23[12]}
   );
   gpc1_1 gpc2528 (
      {stage2_24[27]},
      {stage3_24[15]}
   );
   gpc1_1 gpc2529 (
      {stage2_25[20]},
      {stage3_25[8]}
   );
   gpc1_1 gpc2530 (
      {stage2_25[21]},
      {stage3_25[9]}
   );
   gpc1_1 gpc2531 (
      {stage2_25[22]},
      {stage3_25[10]}
   );
   gpc1_1 gpc2532 (
      {stage2_25[23]},
      {stage3_25[11]}
   );
   gpc1_1 gpc2533 (
      {stage2_25[24]},
      {stage3_25[12]}
   );
   gpc1_1 gpc2534 (
      {stage2_25[25]},
      {stage3_25[13]}
   );
   gpc1_1 gpc2535 (
      {stage2_25[26]},
      {stage3_25[14]}
   );
   gpc1_1 gpc2536 (
      {stage2_25[27]},
      {stage3_25[15]}
   );
   gpc1_1 gpc2537 (
      {stage2_25[28]},
      {stage3_25[16]}
   );
   gpc1_1 gpc2538 (
      {stage2_25[29]},
      {stage3_25[17]}
   );
   gpc1_1 gpc2539 (
      {stage2_25[30]},
      {stage3_25[18]}
   );
   gpc1_1 gpc2540 (
      {stage2_25[31]},
      {stage3_25[19]}
   );
   gpc1_1 gpc2541 (
      {stage2_26[22]},
      {stage3_26[8]}
   );
   gpc1_1 gpc2542 (
      {stage2_26[23]},
      {stage3_26[9]}
   );
   gpc1_1 gpc2543 (
      {stage2_26[24]},
      {stage3_26[10]}
   );
   gpc1_1 gpc2544 (
      {stage2_26[25]},
      {stage3_26[11]}
   );
   gpc1_1 gpc2545 (
      {stage2_26[26]},
      {stage3_26[12]}
   );
   gpc1_1 gpc2546 (
      {stage2_28[21]},
      {stage3_28[11]}
   );
   gpc1_1 gpc2547 (
      {stage2_28[22]},
      {stage3_28[12]}
   );
   gpc1_1 gpc2548 (
      {stage2_28[23]},
      {stage3_28[13]}
   );
   gpc1_1 gpc2549 (
      {stage2_28[24]},
      {stage3_28[14]}
   );
   gpc1_1 gpc2550 (
      {stage2_28[25]},
      {stage3_28[15]}
   );
   gpc1_1 gpc2551 (
      {stage2_28[26]},
      {stage3_28[16]}
   );
   gpc1_1 gpc2552 (
      {stage2_31[24]},
      {stage3_31[16]}
   );
   gpc1_1 gpc2553 (
      {stage2_31[25]},
      {stage3_31[17]}
   );
   gpc1_1 gpc2554 (
      {stage2_31[26]},
      {stage3_31[18]}
   );
   gpc1_1 gpc2555 (
      {stage2_31[27]},
      {stage3_31[19]}
   );
   gpc1_1 gpc2556 (
      {stage2_32[24]},
      {stage3_32[11]}
   );
   gpc1_1 gpc2557 (
      {stage2_34[31]},
      {stage3_34[17]}
   );
   gpc1_1 gpc2558 (
      {stage2_35[29]},
      {stage3_35[9]}
   );
   gpc1_1 gpc2559 (
      {stage2_37[36]},
      {stage3_37[14]}
   );
   gpc1_1 gpc2560 (
      {stage2_40[31]},
      {stage3_40[14]}
   );
   gpc1_1 gpc2561 (
      {stage2_40[32]},
      {stage3_40[15]}
   );
   gpc1_1 gpc2562 (
      {stage2_40[33]},
      {stage3_40[16]}
   );
   gpc1_1 gpc2563 (
      {stage2_40[34]},
      {stage3_40[17]}
   );
   gpc1_1 gpc2564 (
      {stage2_41[30]},
      {stage3_41[10]}
   );
   gpc1_1 gpc2565 (
      {stage2_41[31]},
      {stage3_41[11]}
   );
   gpc1_1 gpc2566 (
      {stage2_42[10]},
      {stage3_42[12]}
   );
   gpc1_1 gpc2567 (
      {stage2_42[11]},
      {stage3_42[13]}
   );
   gpc1_1 gpc2568 (
      {stage2_42[12]},
      {stage3_42[14]}
   );
   gpc1_1 gpc2569 (
      {stage2_42[13]},
      {stage3_42[15]}
   );
   gpc1_1 gpc2570 (
      {stage2_42[14]},
      {stage3_42[16]}
   );
   gpc1_1 gpc2571 (
      {stage2_42[15]},
      {stage3_42[17]}
   );
   gpc1_1 gpc2572 (
      {stage2_42[16]},
      {stage3_42[18]}
   );
   gpc1_1 gpc2573 (
      {stage2_42[17]},
      {stage3_42[19]}
   );
   gpc1_1 gpc2574 (
      {stage2_43[19]},
      {stage3_43[8]}
   );
   gpc1_1 gpc2575 (
      {stage2_43[20]},
      {stage3_43[9]}
   );
   gpc1_1 gpc2576 (
      {stage2_45[33]},
      {stage3_45[13]}
   );
   gpc1_1 gpc2577 (
      {stage2_45[34]},
      {stage3_45[14]}
   );
   gpc1_1 gpc2578 (
      {stage2_46[22]},
      {stage3_46[11]}
   );
   gpc1_1 gpc2579 (
      {stage2_47[35]},
      {stage3_47[10]}
   );
   gpc1_1 gpc2580 (
      {stage2_48[26]},
      {stage3_48[14]}
   );
   gpc1_1 gpc2581 (
      {stage2_48[27]},
      {stage3_48[15]}
   );
   gpc1_1 gpc2582 (
      {stage2_48[28]},
      {stage3_48[16]}
   );
   gpc1_1 gpc2583 (
      {stage2_48[29]},
      {stage3_48[17]}
   );
   gpc1_1 gpc2584 (
      {stage2_48[30]},
      {stage3_48[18]}
   );
   gpc1_1 gpc2585 (
      {stage2_52[11]},
      {stage3_52[13]}
   );
   gpc1_1 gpc2586 (
      {stage2_52[12]},
      {stage3_52[14]}
   );
   gpc1_1 gpc2587 (
      {stage2_52[13]},
      {stage3_52[15]}
   );
   gpc1_1 gpc2588 (
      {stage2_52[14]},
      {stage3_52[16]}
   );
   gpc1_1 gpc2589 (
      {stage2_52[15]},
      {stage3_52[17]}
   );
   gpc1_1 gpc2590 (
      {stage2_52[16]},
      {stage3_52[18]}
   );
   gpc1_1 gpc2591 (
      {stage2_52[17]},
      {stage3_52[19]}
   );
   gpc1_1 gpc2592 (
      {stage2_53[37]},
      {stage3_53[7]}
   );
   gpc1_1 gpc2593 (
      {stage2_53[38]},
      {stage3_53[8]}
   );
   gpc1_1 gpc2594 (
      {stage2_54[15]},
      {stage3_54[10]}
   );
   gpc1_1 gpc2595 (
      {stage2_54[16]},
      {stage3_54[11]}
   );
   gpc1_1 gpc2596 (
      {stage2_54[17]},
      {stage3_54[12]}
   );
   gpc1_1 gpc2597 (
      {stage2_54[18]},
      {stage3_54[13]}
   );
   gpc1_1 gpc2598 (
      {stage2_54[19]},
      {stage3_54[14]}
   );
   gpc1_1 gpc2599 (
      {stage2_54[20]},
      {stage3_54[15]}
   );
   gpc1_1 gpc2600 (
      {stage2_54[21]},
      {stage3_54[16]}
   );
   gpc1_1 gpc2601 (
      {stage2_54[22]},
      {stage3_54[17]}
   );
   gpc1_1 gpc2602 (
      {stage2_54[23]},
      {stage3_54[18]}
   );
   gpc1_1 gpc2603 (
      {stage2_54[24]},
      {stage3_54[19]}
   );
   gpc1_1 gpc2604 (
      {stage2_54[25]},
      {stage3_54[20]}
   );
   gpc1_1 gpc2605 (
      {stage2_54[26]},
      {stage3_54[21]}
   );
   gpc1_1 gpc2606 (
      {stage2_54[27]},
      {stage3_54[22]}
   );
   gpc1_1 gpc2607 (
      {stage2_54[28]},
      {stage3_54[23]}
   );
   gpc1_1 gpc2608 (
      {stage2_55[18]},
      {stage3_55[10]}
   );
   gpc1_1 gpc2609 (
      {stage2_55[19]},
      {stage3_55[11]}
   );
   gpc1_1 gpc2610 (
      {stage2_59[30]},
      {stage3_59[9]}
   );
   gpc1_1 gpc2611 (
      {stage2_59[31]},
      {stage3_59[10]}
   );
   gpc1_1 gpc2612 (
      {stage2_59[32]},
      {stage3_59[11]}
   );
   gpc1_1 gpc2613 (
      {stage2_59[33]},
      {stage3_59[12]}
   );
   gpc1_1 gpc2614 (
      {stage2_59[34]},
      {stage3_59[13]}
   );
   gpc1_1 gpc2615 (
      {stage2_60[21]},
      {stage3_60[13]}
   );
   gpc1_1 gpc2616 (
      {stage2_61[20]},
      {stage3_61[12]}
   );
   gpc1_1 gpc2617 (
      {stage2_61[21]},
      {stage3_61[13]}
   );
   gpc1_1 gpc2618 (
      {stage2_61[22]},
      {stage3_61[14]}
   );
   gpc1_1 gpc2619 (
      {stage2_61[23]},
      {stage3_61[15]}
   );
   gpc1_1 gpc2620 (
      {stage2_61[24]},
      {stage3_61[16]}
   );
   gpc1_1 gpc2621 (
      {stage2_61[25]},
      {stage3_61[17]}
   );
   gpc1_1 gpc2622 (
      {stage2_61[26]},
      {stage3_61[18]}
   );
   gpc1_1 gpc2623 (
      {stage2_61[27]},
      {stage3_61[19]}
   );
   gpc1_1 gpc2624 (
      {stage2_61[28]},
      {stage3_61[20]}
   );
   gpc1_1 gpc2625 (
      {stage2_62[30]},
      {stage3_62[8]}
   );
   gpc1_1 gpc2626 (
      {stage2_62[31]},
      {stage3_62[9]}
   );
   gpc1_1 gpc2627 (
      {stage2_62[32]},
      {stage3_62[10]}
   );
   gpc1_1 gpc2628 (
      {stage2_62[33]},
      {stage3_62[11]}
   );
   gpc1_1 gpc2629 (
      {stage2_62[34]},
      {stage3_62[12]}
   );
   gpc1_1 gpc2630 (
      {stage2_62[35]},
      {stage3_62[13]}
   );
   gpc1_1 gpc2631 (
      {stage2_62[36]},
      {stage3_62[14]}
   );
   gpc1_1 gpc2632 (
      {stage2_62[37]},
      {stage3_62[15]}
   );
   gpc1_1 gpc2633 (
      {stage2_63[33]},
      {stage3_63[13]}
   );
   gpc1_1 gpc2634 (
      {stage2_63[34]},
      {stage3_63[14]}
   );
   gpc1_1 gpc2635 (
      {stage2_63[35]},
      {stage3_63[15]}
   );
   gpc1_1 gpc2636 (
      {stage2_63[36]},
      {stage3_63[16]}
   );
   gpc1_1 gpc2637 (
      {stage2_63[37]},
      {stage3_63[17]}
   );
   gpc1_1 gpc2638 (
      {stage2_65[15]},
      {stage3_65[9]}
   );
   gpc1_1 gpc2639 (
      {stage2_65[16]},
      {stage3_65[10]}
   );
   gpc1_1 gpc2640 (
      {stage2_65[17]},
      {stage3_65[11]}
   );
   gpc1_1 gpc2641 (
      {stage2_66[5]},
      {stage3_66[6]}
   );
   gpc1_1 gpc2642 (
      {stage2_67[0]},
      {stage3_67[5]}
   );
   gpc1_1 gpc2643 (
      {stage2_67[1]},
      {stage3_67[6]}
   );
   gpc615_5 gpc2644 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc207_4 gpc2645 (
      {stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7]},
      {stage3_3[0], stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc2646 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc2647 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[1]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[1],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc2648 (
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16]},
      {stage3_4[2]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[2],stage4_5[2],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc2649 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[3],stage4_6[3]}
   );
   gpc615_5 gpc2650 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[4]}
   );
   gpc615_5 gpc2651 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[5]}
   );
   gpc606_5 gpc2652 (
      {stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[2],stage4_10[3],stage4_9[3],stage4_8[3]}
   );
   gpc606_5 gpc2653 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[3],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc2654 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[2],stage4_11[4]}
   );
   gpc207_4 gpc2655 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[3]}
   );
   gpc606_5 gpc2656 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage4_16[0],stage4_15[2],stage4_14[2],stage4_13[3],stage4_12[4]}
   );
   gpc606_5 gpc2657 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[3],stage4_14[3],stage4_13[4]}
   );
   gpc207_4 gpc2658 (
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage3_17[0], stage3_17[1]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[4]}
   );
   gpc207_4 gpc2659 (
      {stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_17[2], stage3_17[3]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[5]}
   );
   gpc615_5 gpc2660 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[0]},
      {stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9]},
      {stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4],stage4_15[6]}
   );
   gpc606_5 gpc2661 (
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[1],stage4_18[3],stage4_17[4],stage4_16[5]}
   );
   gpc606_5 gpc2662 (
      {stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11], 1'b0},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[2],stage4_18[4],stage4_17[5],stage4_16[6]}
   );
   gpc615_5 gpc2663 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[3]}
   );
   gpc615_5 gpc2664 (
      {stage3_19[5], stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9]},
      {stage3_20[1]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[4]}
   );
   gpc615_5 gpc2665 (
      {stage3_19[10], stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14]},
      {stage3_20[2]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[5]}
   );
   gpc606_5 gpc2666 (
      {stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[3],stage4_22[3],stage4_21[3],stage4_20[5]}
   );
   gpc1163_5 gpc2667 (
      {stage3_22[6], stage3_22[7], stage3_22[8]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage3_24[0]},
      {stage3_25[0]},
      {stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[4],stage4_22[4]}
   );
   gpc117_4 gpc2668 (
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12]},
      {stage3_24[1]},
      {stage3_25[1]},
      {stage4_26[1],stage4_25[1],stage4_24[2],stage4_23[5]}
   );
   gpc207_4 gpc2669 (
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7], stage3_24[8]},
      {stage3_26[0], stage3_26[1]},
      {stage4_27[0],stage4_26[2],stage4_25[2],stage4_24[3]}
   );
   gpc135_4 gpc2670 (
      {stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage3_26[2], stage3_26[3], stage3_26[4]},
      {stage3_27[0]},
      {stage4_28[0],stage4_27[1],stage4_26[3],stage4_25[3]}
   );
   gpc135_4 gpc2671 (
      {stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage3_26[5], stage3_26[6], stage3_26[7]},
      {stage3_27[1]},
      {stage4_28[1],stage4_27[2],stage4_26[4],stage4_25[4]}
   );
   gpc606_5 gpc2672 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5], stage3_27[6], stage3_27[7]},
      {stage4_29[0],stage4_28[2],stage4_27[3],stage4_26[5],stage4_25[5]}
   );
   gpc1163_5 gpc2673 (
      {stage3_27[8], stage3_27[9], stage3_27[10]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage3_29[0]},
      {stage3_30[0]},
      {stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[3],stage4_27[4]}
   );
   gpc1163_5 gpc2674 (
      {stage3_27[11], stage3_27[12], stage3_27[13]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage3_29[1]},
      {stage3_30[1]},
      {stage4_31[1],stage4_30[1],stage4_29[2],stage4_28[4],stage4_27[5]}
   );
   gpc606_5 gpc2675 (
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], 1'b0},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7]},
      {stage4_32[0],stage4_31[2],stage4_30[2],stage4_29[3],stage4_28[5]}
   );
   gpc207_4 gpc2676 (
      {stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13], stage3_30[14]},
      {stage3_32[0], stage3_32[1]},
      {stage4_33[0],stage4_32[1],stage4_31[3],stage4_30[3]}
   );
   gpc207_4 gpc2677 (
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage3_33[0], stage3_33[1]},
      {stage4_34[0],stage4_33[1],stage4_32[2],stage4_31[4]}
   );
   gpc207_4 gpc2678 (
      {stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13]},
      {stage3_33[2], stage3_33[3]},
      {stage4_34[1],stage4_33[2],stage4_32[3],stage4_31[5]}
   );
   gpc606_5 gpc2679 (
      {stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19]},
      {stage3_33[4], stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage4_35[0],stage4_34[2],stage4_33[3],stage4_32[4],stage4_31[6]}
   );
   gpc615_5 gpc2680 (
      {stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5], stage3_32[6]},
      {stage3_33[10]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[1],stage4_34[3],stage4_33[4],stage4_32[5]}
   );
   gpc615_5 gpc2681 (
      {stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_33[11]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[2],stage4_34[4],stage4_33[5],stage4_32[6]}
   );
   gpc606_5 gpc2682 (
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage4_38[0],stage4_37[0],stage4_36[2],stage4_35[3],stage4_34[5]}
   );
   gpc117_4 gpc2683 (
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5], stage3_35[6]},
      {stage3_36[6]},
      {stage3_37[0]},
      {stage4_38[1],stage4_37[1],stage4_36[3],stage4_35[4]}
   );
   gpc1163_5 gpc2684 (
      {stage3_35[7], stage3_35[8], stage3_35[9]},
      {stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11], stage3_36[12]},
      {stage3_37[1]},
      {stage3_38[0]},
      {stage4_39[0],stage4_38[2],stage4_37[2],stage4_36[4],stage4_35[5]}
   );
   gpc1163_5 gpc2685 (
      {stage3_37[2], stage3_37[3], stage3_37[4]},
      {stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5], stage3_38[6]},
      {stage3_39[0]},
      {stage3_40[0]},
      {stage4_41[0],stage4_40[0],stage4_39[1],stage4_38[3],stage4_37[3]}
   );
   gpc1163_5 gpc2686 (
      {stage3_37[5], stage3_37[6], stage3_37[7]},
      {stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11], stage3_38[12]},
      {stage3_39[1]},
      {stage3_40[1]},
      {stage4_41[1],stage4_40[1],stage4_39[2],stage4_38[4],stage4_37[4]}
   );
   gpc606_5 gpc2687 (
      {stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11], stage3_37[12], stage3_37[13]},
      {stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5], stage3_39[6], stage3_39[7]},
      {stage4_41[2],stage4_40[2],stage4_39[3],stage4_38[5],stage4_37[5]}
   );
   gpc223_4 gpc2688 (
      {stage3_39[8], stage3_39[9], stage3_39[10]},
      {stage3_40[2], stage3_40[3]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[0],stage4_41[3],stage4_40[3],stage4_39[4]}
   );
   gpc623_5 gpc2689 (
      {stage3_40[4], stage3_40[5], stage3_40[6]},
      {stage3_41[2], stage3_41[3]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage4_44[0],stage4_43[0],stage4_42[1],stage4_41[4],stage4_40[4]}
   );
   gpc623_5 gpc2690 (
      {stage3_40[7], stage3_40[8], stage3_40[9]},
      {stage3_41[4], stage3_41[5]},
      {stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11]},
      {stage4_44[1],stage4_43[1],stage4_42[2],stage4_41[5],stage4_40[5]}
   );
   gpc623_5 gpc2691 (
      {stage3_40[10], stage3_40[11], stage3_40[12]},
      {stage3_41[6], stage3_41[7]},
      {stage3_42[12], stage3_42[13], stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17]},
      {stage4_44[2],stage4_43[2],stage4_42[3],stage4_41[6],stage4_40[6]}
   );
   gpc615_5 gpc2692 (
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4]},
      {stage3_44[0]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[0],stage4_45[0],stage4_44[3],stage4_43[3]}
   );
   gpc615_5 gpc2693 (
      {stage3_43[5], stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9]},
      {stage3_44[1]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[1],stage4_45[1],stage4_44[4],stage4_43[4]}
   );
   gpc207_4 gpc2694 (
      {stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5], stage3_44[6], stage3_44[7], 1'b0},
      {stage3_46[0], stage3_46[1]},
      {stage4_47[2],stage4_46[2],stage4_45[2],stage4_44[5]}
   );
   gpc606_5 gpc2695 (
      {stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6], stage3_46[7]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[0],stage4_47[3],stage4_46[3]}
   );
   gpc623_5 gpc2696 (
      {stage3_46[8], stage3_46[9], stage3_46[10]},
      {stage3_47[0], stage3_47[1]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[1],stage4_48[1],stage4_47[4],stage4_46[4]}
   );
   gpc135_4 gpc2697 (
      {stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6]},
      {stage3_48[12], stage3_48[13], stage3_48[14]},
      {stage3_49[0]},
      {stage4_50[2],stage4_49[2],stage4_48[2],stage4_47[5]}
   );
   gpc135_4 gpc2698 (
      {stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], 1'b0},
      {stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage3_49[1]},
      {stage4_50[3],stage4_49[3],stage4_48[3],stage4_47[6]}
   );
   gpc615_5 gpc2699 (
      {stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5], stage3_49[6]},
      {stage3_50[0]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[0],stage4_50[4],stage4_49[4]}
   );
   gpc615_5 gpc2700 (
      {stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage3_50[1]},
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage4_53[1],stage4_52[1],stage4_51[1],stage4_50[5],stage4_49[5]}
   );
   gpc615_5 gpc2701 (
      {stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[12]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[2],stage4_52[2],stage4_51[2],stage4_50[6]}
   );
   gpc1343_5 gpc2702 (
      {stage3_53[0], stage3_53[1], stage3_53[2]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3]},
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[0],stage4_55[0],stage4_54[1],stage4_53[3]}
   );
   gpc1343_5 gpc2703 (
      {stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage3_54[4], stage3_54[5], stage3_54[6], stage3_54[7]},
      {stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_56[1]},
      {stage4_57[1],stage4_56[1],stage4_55[1],stage4_54[2],stage4_53[4]}
   );
   gpc1343_5 gpc2704 (
      {stage3_53[6], stage3_53[7], stage3_53[8]},
      {stage3_54[8], stage3_54[9], stage3_54[10], stage3_54[11]},
      {stage3_55[6], stage3_55[7], stage3_55[8]},
      {stage3_56[2]},
      {stage4_57[2],stage4_56[2],stage4_55[2],stage4_54[3],stage4_53[5]}
   );
   gpc135_4 gpc2705 (
      {stage3_54[12], stage3_54[13], stage3_54[14], stage3_54[15], stage3_54[16]},
      {stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage3_56[3]},
      {stage4_57[3],stage4_56[3],stage4_55[3],stage4_54[4]}
   );
   gpc606_5 gpc2706 (
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[0],stage4_58[0],stage4_57[4]}
   );
   gpc606_5 gpc2707 (
      {stage3_57[6], stage3_57[7], stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11]},
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage4_61[1],stage4_60[1],stage4_59[1],stage4_58[1],stage4_57[5]}
   );
   gpc207_4 gpc2708 (
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5], stage3_58[6]},
      {stage3_60[0], stage3_60[1]},
      {stage4_61[2],stage4_60[2],stage4_59[2],stage4_58[2]}
   );
   gpc207_4 gpc2709 (
      {stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11], 1'b0, 1'b0},
      {stage3_60[2], stage3_60[3]},
      {stage4_61[3],stage4_60[3],stage4_59[3],stage4_58[3]}
   );
   gpc606_5 gpc2710 (
      {stage3_60[4], stage3_60[5], stage3_60[6], stage3_60[7], stage3_60[8], stage3_60[9]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[0],stage4_62[0],stage4_61[4],stage4_60[4]}
   );
   gpc606_5 gpc2711 (
      {stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], 1'b0, 1'b0},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[1],stage4_62[1],stage4_61[5],stage4_60[5]}
   );
   gpc117_4 gpc2712 (
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5], stage3_61[6]},
      {stage3_62[12]},
      {stage3_63[0]},
      {stage4_64[2],stage4_63[2],stage4_62[2],stage4_61[6]}
   );
   gpc207_4 gpc2713 (
      {stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11], stage3_61[12], stage3_61[13]},
      {stage3_63[1], stage3_63[2]},
      {stage4_64[3],stage4_63[3],stage4_62[3],stage4_61[7]}
   );
   gpc606_5 gpc2714 (
      {stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17], stage3_61[18], stage3_61[19]},
      {stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6], stage3_63[7], stage3_63[8]},
      {stage4_65[0],stage4_64[4],stage4_63[4],stage4_62[4],stage4_61[8]}
   );
   gpc615_5 gpc2715 (
      {stage3_62[13], stage3_62[14], stage3_62[15], 1'b0, 1'b0},
      {stage3_63[9]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[1],stage4_64[5],stage4_63[5],stage4_62[5]}
   );
   gpc606_5 gpc2716 (
      {stage3_63[10], stage3_63[11], stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[1],stage4_65[2],stage4_64[6],stage4_63[6]}
   );
   gpc606_5 gpc2717 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[2],stage4_65[3],stage4_64[7]}
   );
   gpc606_5 gpc2718 (
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage3_67[0], stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5]},
      {stage4_69[0],stage4_68[1],stage4_67[2],stage4_66[3],stage4_65[4]}
   );
   gpc1_1 gpc2719 (
      {stage3_3[17]},
      {stage4_3[5]}
   );
   gpc1_1 gpc2720 (
      {stage3_3[18]},
      {stage4_3[6]}
   );
   gpc1_1 gpc2721 (
      {stage3_3[19]},
      {stage4_3[7]}
   );
   gpc1_1 gpc2722 (
      {stage3_3[20]},
      {stage4_3[8]}
   );
   gpc1_1 gpc2723 (
      {stage3_3[21]},
      {stage4_3[9]}
   );
   gpc1_1 gpc2724 (
      {stage3_4[3]},
      {stage4_4[5]}
   );
   gpc1_1 gpc2725 (
      {stage3_4[4]},
      {stage4_4[6]}
   );
   gpc1_1 gpc2726 (
      {stage3_4[5]},
      {stage4_4[7]}
   );
   gpc1_1 gpc2727 (
      {stage3_4[6]},
      {stage4_4[8]}
   );
   gpc1_1 gpc2728 (
      {stage3_4[7]},
      {stage4_4[9]}
   );
   gpc1_1 gpc2729 (
      {stage3_4[8]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2730 (
      {stage3_4[9]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2731 (
      {stage3_4[10]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2732 (
      {stage3_4[11]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2733 (
      {stage3_5[18]},
      {stage4_5[3]}
   );
   gpc1_1 gpc2734 (
      {stage3_5[19]},
      {stage4_5[4]}
   );
   gpc1_1 gpc2735 (
      {stage3_5[20]},
      {stage4_5[5]}
   );
   gpc1_1 gpc2736 (
      {stage3_5[21]},
      {stage4_5[6]}
   );
   gpc1_1 gpc2737 (
      {stage3_5[22]},
      {stage4_5[7]}
   );
   gpc1_1 gpc2738 (
      {stage3_5[23]},
      {stage4_5[8]}
   );
   gpc1_1 gpc2739 (
      {stage3_6[5]},
      {stage4_6[4]}
   );
   gpc1_1 gpc2740 (
      {stage3_6[6]},
      {stage4_6[5]}
   );
   gpc1_1 gpc2741 (
      {stage3_6[7]},
      {stage4_6[6]}
   );
   gpc1_1 gpc2742 (
      {stage3_6[8]},
      {stage4_6[7]}
   );
   gpc1_1 gpc2743 (
      {stage3_6[9]},
      {stage4_6[8]}
   );
   gpc1_1 gpc2744 (
      {stage3_7[11]},
      {stage4_7[6]}
   );
   gpc1_1 gpc2745 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc2746 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc2747 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc2748 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc2749 (
      {stage3_10[6]},
      {stage4_10[5]}
   );
   gpc1_1 gpc2750 (
      {stage3_10[7]},
      {stage4_10[6]}
   );
   gpc1_1 gpc2751 (
      {stage3_10[8]},
      {stage4_10[7]}
   );
   gpc1_1 gpc2752 (
      {stage3_10[9]},
      {stage4_10[8]}
   );
   gpc1_1 gpc2753 (
      {stage3_10[10]},
      {stage4_10[9]}
   );
   gpc1_1 gpc2754 (
      {stage3_10[11]},
      {stage4_10[10]}
   );
   gpc1_1 gpc2755 (
      {stage3_11[12]},
      {stage4_11[5]}
   );
   gpc1_1 gpc2756 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc2757 (
      {stage3_14[8]},
      {stage4_14[4]}
   );
   gpc1_1 gpc2758 (
      {stage3_14[9]},
      {stage4_14[5]}
   );
   gpc1_1 gpc2759 (
      {stage3_15[25]},
      {stage4_15[7]}
   );
   gpc1_1 gpc2760 (
      {stage3_17[10]},
      {stage4_17[6]}
   );
   gpc1_1 gpc2761 (
      {stage3_17[11]},
      {stage4_17[7]}
   );
   gpc1_1 gpc2762 (
      {stage3_18[12]},
      {stage4_18[5]}
   );
   gpc1_1 gpc2763 (
      {stage3_19[15]},
      {stage4_19[6]}
   );
   gpc1_1 gpc2764 (
      {stage3_20[9]},
      {stage4_20[6]}
   );
   gpc1_1 gpc2765 (
      {stage3_20[10]},
      {stage4_20[7]}
   );
   gpc1_1 gpc2766 (
      {stage3_20[11]},
      {stage4_20[8]}
   );
   gpc1_1 gpc2767 (
      {stage3_20[12]},
      {stage4_20[9]}
   );
   gpc1_1 gpc2768 (
      {stage3_20[13]},
      {stage4_20[10]}
   );
   gpc1_1 gpc2769 (
      {stage3_24[9]},
      {stage4_24[4]}
   );
   gpc1_1 gpc2770 (
      {stage3_24[10]},
      {stage4_24[5]}
   );
   gpc1_1 gpc2771 (
      {stage3_24[11]},
      {stage4_24[6]}
   );
   gpc1_1 gpc2772 (
      {stage3_24[12]},
      {stage4_24[7]}
   );
   gpc1_1 gpc2773 (
      {stage3_24[13]},
      {stage4_24[8]}
   );
   gpc1_1 gpc2774 (
      {stage3_24[14]},
      {stage4_24[9]}
   );
   gpc1_1 gpc2775 (
      {stage3_24[15]},
      {stage4_24[10]}
   );
   gpc1_1 gpc2776 (
      {stage3_25[18]},
      {stage4_25[6]}
   );
   gpc1_1 gpc2777 (
      {stage3_25[19]},
      {stage4_25[7]}
   );
   gpc1_1 gpc2778 (
      {stage3_26[8]},
      {stage4_26[6]}
   );
   gpc1_1 gpc2779 (
      {stage3_26[9]},
      {stage4_26[7]}
   );
   gpc1_1 gpc2780 (
      {stage3_26[10]},
      {stage4_26[8]}
   );
   gpc1_1 gpc2781 (
      {stage3_26[11]},
      {stage4_26[9]}
   );
   gpc1_1 gpc2782 (
      {stage3_26[12]},
      {stage4_26[10]}
   );
   gpc1_1 gpc2783 (
      {stage3_29[2]},
      {stage4_29[4]}
   );
   gpc1_1 gpc2784 (
      {stage3_29[3]},
      {stage4_29[5]}
   );
   gpc1_1 gpc2785 (
      {stage3_29[4]},
      {stage4_29[6]}
   );
   gpc1_1 gpc2786 (
      {stage3_29[5]},
      {stage4_29[7]}
   );
   gpc1_1 gpc2787 (
      {stage3_29[6]},
      {stage4_29[8]}
   );
   gpc1_1 gpc2788 (
      {stage3_29[7]},
      {stage4_29[9]}
   );
   gpc1_1 gpc2789 (
      {stage3_36[13]},
      {stage4_36[5]}
   );
   gpc1_1 gpc2790 (
      {stage3_36[14]},
      {stage4_36[6]}
   );
   gpc1_1 gpc2791 (
      {stage3_37[14]},
      {stage4_37[6]}
   );
   gpc1_1 gpc2792 (
      {stage3_39[11]},
      {stage4_39[5]}
   );
   gpc1_1 gpc2793 (
      {stage3_39[12]},
      {stage4_39[6]}
   );
   gpc1_1 gpc2794 (
      {stage3_39[13]},
      {stage4_39[7]}
   );
   gpc1_1 gpc2795 (
      {stage3_40[13]},
      {stage4_40[7]}
   );
   gpc1_1 gpc2796 (
      {stage3_40[14]},
      {stage4_40[8]}
   );
   gpc1_1 gpc2797 (
      {stage3_40[15]},
      {stage4_40[9]}
   );
   gpc1_1 gpc2798 (
      {stage3_40[16]},
      {stage4_40[10]}
   );
   gpc1_1 gpc2799 (
      {stage3_40[17]},
      {stage4_40[11]}
   );
   gpc1_1 gpc2800 (
      {stage3_41[8]},
      {stage4_41[7]}
   );
   gpc1_1 gpc2801 (
      {stage3_41[9]},
      {stage4_41[8]}
   );
   gpc1_1 gpc2802 (
      {stage3_41[10]},
      {stage4_41[9]}
   );
   gpc1_1 gpc2803 (
      {stage3_41[11]},
      {stage4_41[10]}
   );
   gpc1_1 gpc2804 (
      {stage3_42[18]},
      {stage4_42[4]}
   );
   gpc1_1 gpc2805 (
      {stage3_42[19]},
      {stage4_42[5]}
   );
   gpc1_1 gpc2806 (
      {stage3_45[12]},
      {stage4_45[3]}
   );
   gpc1_1 gpc2807 (
      {stage3_45[13]},
      {stage4_45[4]}
   );
   gpc1_1 gpc2808 (
      {stage3_45[14]},
      {stage4_45[5]}
   );
   gpc1_1 gpc2809 (
      {stage3_46[11]},
      {stage4_46[5]}
   );
   gpc1_1 gpc2810 (
      {stage3_48[18]},
      {stage4_48[4]}
   );
   gpc1_1 gpc2811 (
      {stage3_52[6]},
      {stage4_52[3]}
   );
   gpc1_1 gpc2812 (
      {stage3_52[7]},
      {stage4_52[4]}
   );
   gpc1_1 gpc2813 (
      {stage3_52[8]},
      {stage4_52[5]}
   );
   gpc1_1 gpc2814 (
      {stage3_52[9]},
      {stage4_52[6]}
   );
   gpc1_1 gpc2815 (
      {stage3_52[10]},
      {stage4_52[7]}
   );
   gpc1_1 gpc2816 (
      {stage3_52[11]},
      {stage4_52[8]}
   );
   gpc1_1 gpc2817 (
      {stage3_52[12]},
      {stage4_52[9]}
   );
   gpc1_1 gpc2818 (
      {stage3_52[13]},
      {stage4_52[10]}
   );
   gpc1_1 gpc2819 (
      {stage3_52[14]},
      {stage4_52[11]}
   );
   gpc1_1 gpc2820 (
      {stage3_52[15]},
      {stage4_52[12]}
   );
   gpc1_1 gpc2821 (
      {stage3_52[16]},
      {stage4_52[13]}
   );
   gpc1_1 gpc2822 (
      {stage3_52[17]},
      {stage4_52[14]}
   );
   gpc1_1 gpc2823 (
      {stage3_52[18]},
      {stage4_52[15]}
   );
   gpc1_1 gpc2824 (
      {stage3_52[19]},
      {stage4_52[16]}
   );
   gpc1_1 gpc2825 (
      {stage3_54[17]},
      {stage4_54[5]}
   );
   gpc1_1 gpc2826 (
      {stage3_54[18]},
      {stage4_54[6]}
   );
   gpc1_1 gpc2827 (
      {stage3_54[19]},
      {stage4_54[7]}
   );
   gpc1_1 gpc2828 (
      {stage3_54[20]},
      {stage4_54[8]}
   );
   gpc1_1 gpc2829 (
      {stage3_54[21]},
      {stage4_54[9]}
   );
   gpc1_1 gpc2830 (
      {stage3_54[22]},
      {stage4_54[10]}
   );
   gpc1_1 gpc2831 (
      {stage3_54[23]},
      {stage4_54[11]}
   );
   gpc1_1 gpc2832 (
      {stage3_56[4]},
      {stage4_56[4]}
   );
   gpc1_1 gpc2833 (
      {stage3_56[5]},
      {stage4_56[5]}
   );
   gpc1_1 gpc2834 (
      {stage3_56[6]},
      {stage4_56[6]}
   );
   gpc1_1 gpc2835 (
      {stage3_56[7]},
      {stage4_56[7]}
   );
   gpc1_1 gpc2836 (
      {stage3_59[12]},
      {stage4_59[4]}
   );
   gpc1_1 gpc2837 (
      {stage3_59[13]},
      {stage4_59[5]}
   );
   gpc1_1 gpc2838 (
      {stage3_61[20]},
      {stage4_61[9]}
   );
   gpc1_1 gpc2839 (
      {stage3_63[16]},
      {stage4_63[7]}
   );
   gpc1_1 gpc2840 (
      {stage3_63[17]},
      {stage4_63[8]}
   );
   gpc1_1 gpc2841 (
      {stage3_64[12]},
      {stage4_64[8]}
   );
   gpc1_1 gpc2842 (
      {stage3_66[6]},
      {stage4_66[4]}
   );
   gpc1_1 gpc2843 (
      {stage3_67[6]},
      {stage4_67[3]}
   );
   gpc117_4 gpc2844 (
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_4[0]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0]}
   );
   gpc606_5 gpc2845 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1]}
   );
   gpc1325_5 gpc2846 (
      {stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_5[1], stage4_5[2]},
      {stage4_6[6], stage4_6[7], stage4_6[8]},
      {stage4_7[0]},
      {stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc606_5 gpc2847 (
      {stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7], stage4_5[8]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc606_5 gpc2848 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[3]}
   );
   gpc606_5 gpc2849 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1],stage5_9[2]}
   );
   gpc623_5 gpc2850 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[2]}
   );
   gpc615_5 gpc2851 (
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4]},
      {stage4_17[0]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[1]}
   );
   gpc606_5 gpc2852 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[1],stage5_17[1]}
   );
   gpc15_3 gpc2853 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[1],stage5_20[2]}
   );
   gpc1163_5 gpc2854 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[1]}
   );
   gpc606_5 gpc2855 (
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[0],stage5_26[1],stage5_25[1],stage5_24[1]}
   );
   gpc7_3 gpc2856 (
      {stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6], stage4_25[7]},
      {stage5_27[1],stage5_26[2],stage5_25[2]}
   );
   gpc615_5 gpc2857 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[3]}
   );
   gpc606_5 gpc2858 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[1]}
   );
   gpc623_5 gpc2859 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[6], 1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[2]}
   );
   gpc606_5 gpc2860 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[1],stage5_33[2]}
   );
   gpc7_3 gpc2861 (
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6]},
      {stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc7_3 gpc2862 (
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5], stage4_37[6]},
      {stage5_39[0],stage5_38[1],stage5_37[2]}
   );
   gpc615_5 gpc2863 (
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4]},
      {stage4_39[0]},
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage5_42[0],stage5_41[0],stage5_40[0],stage5_39[1],stage5_38[2]}
   );
   gpc615_5 gpc2864 (
      {stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5]},
      {stage4_40[6]},
      {stage4_41[0], stage4_41[1], stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5]},
      {stage5_43[0],stage5_42[1],stage5_41[1],stage5_40[1],stage5_39[2]}
   );
   gpc606_5 gpc2865 (
      {stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11], 1'b0},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[2],stage5_41[2],stage5_40[2]}
   );
   gpc15_3 gpc2866 (
      {stage4_41[6], stage4_41[7], stage4_41[8], stage4_41[9], stage4_41[10]},
      {1'b0},
      {stage5_43[2],stage5_42[3],stage5_41[3]}
   );
   gpc606_5 gpc2867 (
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], 1'b0},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[0],stage5_44[1],stage5_43[3]}
   );
   gpc615_5 gpc2868 (
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4]},
      {1'b0},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[1],stage5_46[1],stage5_45[1],stage5_44[2]}
   );
   gpc615_5 gpc2869 (
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[0],stage5_49[0],stage5_48[1],stage5_47[2]}
   );
   gpc117_4 gpc2870 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage4_51[0]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[1],stage5_50[1]}
   );
   gpc615_5 gpc2871 (
      {stage4_51[1], stage4_51[2], 1'b0, 1'b0, 1'b0},
      {stage4_52[1]},
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage5_55[0],stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[2]}
   );
   gpc606_5 gpc2872 (
      {stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5], stage4_52[6], stage4_52[7]},
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5]},
      {stage5_56[0],stage5_55[1],stage5_54[1],stage5_53[2],stage5_52[2]}
   );
   gpc606_5 gpc2873 (
      {stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11], stage4_52[12], stage4_52[13]},
      {stage4_54[6], stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11]},
      {stage5_56[1],stage5_55[2],stage5_54[2],stage5_53[3],stage5_52[3]}
   );
   gpc1415_5 gpc2874 (
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], 1'b0},
      {stage4_56[0]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3]},
      {stage4_58[0]},
      {stage5_59[0],stage5_58[0],stage5_57[0],stage5_56[2],stage5_55[3]}
   );
   gpc135_4 gpc2875 (
      {stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage4_57[4], stage4_57[5], 1'b0},
      {stage4_58[1]},
      {stage5_59[1],stage5_58[1],stage5_57[1],stage5_56[3]}
   );
   gpc606_5 gpc2876 (
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[0],stage5_59[2]}
   );
   gpc606_5 gpc2877 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[1]}
   );
   gpc1325_5 gpc2878 (
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], 1'b0},
      {1'b0, 1'b0},
      {stage4_63[0], stage4_63[1], stage4_63[2]},
      {stage4_64[0]},
      {stage5_65[0],stage5_64[1],stage5_63[2],stage5_62[2],stage5_61[2]}
   );
   gpc606_5 gpc2879 (
      {stage4_63[3], stage4_63[4], stage4_63[5], stage4_63[6], stage4_63[7], stage4_63[8]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], 1'b0},
      {stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[2],stage5_63[3]}
   );
   gpc606_5 gpc2880 (
      {stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], 1'b0},
      {stage5_68[0],stage5_67[1],stage5_66[1],stage5_65[2],stage5_64[3]}
   );
   gpc2135_5 gpc2881 (
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], 1'b0},
      {stage4_68[0], stage4_68[1], 1'b0},
      {stage4_69[0]},
      {1'b0, 1'b0},
      {stage5_70[0],stage5_69[0],stage5_68[1],stage5_67[2]}
   );
   gpc1_1 gpc2882 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc2883 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2884 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2885 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc2886 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2887 (
      {stage4_3[7]},
      {stage5_3[1]}
   );
   gpc1_1 gpc2888 (
      {stage4_3[8]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2889 (
      {stage4_3[9]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2890 (
      {stage4_4[12]},
      {stage5_4[3]}
   );
   gpc1_1 gpc2891 (
      {stage4_4[13]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2892 (
      {stage4_9[6]},
      {stage5_9[3]}
   );
   gpc1_1 gpc2893 (
      {stage4_10[6]},
      {stage5_10[2]}
   );
   gpc1_1 gpc2894 (
      {stage4_10[7]},
      {stage5_10[3]}
   );
   gpc1_1 gpc2895 (
      {stage4_10[8]},
      {stage5_10[4]}
   );
   gpc1_1 gpc2896 (
      {stage4_10[9]},
      {stage5_10[5]}
   );
   gpc1_1 gpc2897 (
      {stage4_10[10]},
      {stage5_10[6]}
   );
   gpc1_1 gpc2898 (
      {stage4_12[3]},
      {stage5_12[3]}
   );
   gpc1_1 gpc2899 (
      {stage4_12[4]},
      {stage5_12[4]}
   );
   gpc1_1 gpc2900 (
      {stage4_12[5]},
      {stage5_12[5]}
   );
   gpc1_1 gpc2901 (
      {stage4_13[2]},
      {stage5_13[2]}
   );
   gpc1_1 gpc2902 (
      {stage4_13[3]},
      {stage5_13[3]}
   );
   gpc1_1 gpc2903 (
      {stage4_13[4]},
      {stage5_13[4]}
   );
   gpc1_1 gpc2904 (
      {stage4_15[0]},
      {stage5_15[1]}
   );
   gpc1_1 gpc2905 (
      {stage4_15[1]},
      {stage5_15[2]}
   );
   gpc1_1 gpc2906 (
      {stage4_15[2]},
      {stage5_15[3]}
   );
   gpc1_1 gpc2907 (
      {stage4_15[3]},
      {stage5_15[4]}
   );
   gpc1_1 gpc2908 (
      {stage4_15[4]},
      {stage5_15[5]}
   );
   gpc1_1 gpc2909 (
      {stage4_15[5]},
      {stage5_15[6]}
   );
   gpc1_1 gpc2910 (
      {stage4_15[6]},
      {stage5_15[7]}
   );
   gpc1_1 gpc2911 (
      {stage4_15[7]},
      {stage5_15[8]}
   );
   gpc1_1 gpc2912 (
      {stage4_16[5]},
      {stage5_16[2]}
   );
   gpc1_1 gpc2913 (
      {stage4_16[6]},
      {stage5_16[3]}
   );
   gpc1_1 gpc2914 (
      {stage4_17[7]},
      {stage5_17[2]}
   );
   gpc1_1 gpc2915 (
      {stage4_19[6]},
      {stage5_19[2]}
   );
   gpc1_1 gpc2916 (
      {stage4_20[5]},
      {stage5_20[3]}
   );
   gpc1_1 gpc2917 (
      {stage4_20[6]},
      {stage5_20[4]}
   );
   gpc1_1 gpc2918 (
      {stage4_20[7]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2919 (
      {stage4_20[8]},
      {stage5_20[6]}
   );
   gpc1_1 gpc2920 (
      {stage4_20[9]},
      {stage5_20[7]}
   );
   gpc1_1 gpc2921 (
      {stage4_20[10]},
      {stage5_20[8]}
   );
   gpc1_1 gpc2922 (
      {stage4_21[1]},
      {stage5_21[2]}
   );
   gpc1_1 gpc2923 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc1_1 gpc2924 (
      {stage4_21[3]},
      {stage5_21[4]}
   );
   gpc1_1 gpc2925 (
      {stage4_22[3]},
      {stage5_22[2]}
   );
   gpc1_1 gpc2926 (
      {stage4_22[4]},
      {stage5_22[3]}
   );
   gpc1_1 gpc2927 (
      {stage4_24[7]},
      {stage5_24[2]}
   );
   gpc1_1 gpc2928 (
      {stage4_24[8]},
      {stage5_24[3]}
   );
   gpc1_1 gpc2929 (
      {stage4_24[9]},
      {stage5_24[4]}
   );
   gpc1_1 gpc2930 (
      {stage4_24[10]},
      {stage5_24[5]}
   );
   gpc1_1 gpc2931 (
      {stage4_27[1]},
      {stage5_27[3]}
   );
   gpc1_1 gpc2932 (
      {stage4_27[2]},
      {stage5_27[4]}
   );
   gpc1_1 gpc2933 (
      {stage4_27[3]},
      {stage5_27[5]}
   );
   gpc1_1 gpc2934 (
      {stage4_27[4]},
      {stage5_27[6]}
   );
   gpc1_1 gpc2935 (
      {stage4_27[5]},
      {stage5_27[7]}
   );
   gpc1_1 gpc2936 (
      {stage4_29[6]},
      {stage5_29[2]}
   );
   gpc1_1 gpc2937 (
      {stage4_29[7]},
      {stage5_29[3]}
   );
   gpc1_1 gpc2938 (
      {stage4_29[8]},
      {stage5_29[4]}
   );
   gpc1_1 gpc2939 (
      {stage4_29[9]},
      {stage5_29[5]}
   );
   gpc1_1 gpc2940 (
      {stage4_30[3]},
      {stage5_30[3]}
   );
   gpc1_1 gpc2941 (
      {stage4_32[6]},
      {stage5_32[2]}
   );
   gpc1_1 gpc2942 (
      {stage4_34[0]},
      {stage5_34[2]}
   );
   gpc1_1 gpc2943 (
      {stage4_34[1]},
      {stage5_34[3]}
   );
   gpc1_1 gpc2944 (
      {stage4_34[2]},
      {stage5_34[4]}
   );
   gpc1_1 gpc2945 (
      {stage4_34[3]},
      {stage5_34[5]}
   );
   gpc1_1 gpc2946 (
      {stage4_34[4]},
      {stage5_34[6]}
   );
   gpc1_1 gpc2947 (
      {stage4_34[5]},
      {stage5_34[7]}
   );
   gpc1_1 gpc2948 (
      {stage4_38[5]},
      {stage5_38[3]}
   );
   gpc1_1 gpc2949 (
      {stage4_39[6]},
      {stage5_39[3]}
   );
   gpc1_1 gpc2950 (
      {stage4_39[7]},
      {stage5_39[4]}
   );
   gpc1_1 gpc2951 (
      {stage4_44[5]},
      {stage5_44[3]}
   );
   gpc1_1 gpc2952 (
      {stage4_47[5]},
      {stage5_47[3]}
   );
   gpc1_1 gpc2953 (
      {stage4_47[6]},
      {stage5_47[4]}
   );
   gpc1_1 gpc2954 (
      {stage4_48[1]},
      {stage5_48[2]}
   );
   gpc1_1 gpc2955 (
      {stage4_48[2]},
      {stage5_48[3]}
   );
   gpc1_1 gpc2956 (
      {stage4_48[3]},
      {stage5_48[4]}
   );
   gpc1_1 gpc2957 (
      {stage4_48[4]},
      {stage5_48[5]}
   );
   gpc1_1 gpc2958 (
      {stage4_52[14]},
      {stage5_52[4]}
   );
   gpc1_1 gpc2959 (
      {stage4_52[15]},
      {stage5_52[5]}
   );
   gpc1_1 gpc2960 (
      {stage4_52[16]},
      {stage5_52[6]}
   );
   gpc1_1 gpc2961 (
      {stage4_56[6]},
      {stage5_56[4]}
   );
   gpc1_1 gpc2962 (
      {stage4_56[7]},
      {stage5_56[5]}
   );
   gpc1_1 gpc2963 (
      {stage4_58[2]},
      {stage5_58[2]}
   );
   gpc1_1 gpc2964 (
      {stage4_58[3]},
      {stage5_58[3]}
   );
   gpc1_1 gpc2965 (
      {stage4_64[7]},
      {stage5_64[4]}
   );
   gpc1_1 gpc2966 (
      {stage4_64[8]},
      {stage5_64[5]}
   );
   gpc1343_5 gpc2967 (
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3]},
      {stage5_5[0], stage5_5[1], stage5_5[2]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc135_4 gpc2968 (
      {stage5_6[1], stage5_6[2], stage5_6[3], 1'b0, 1'b0},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1343_5 gpc2969 (
      {stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc615_5 gpc2970 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], 1'b0},
      {stage5_11[1]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1],stage6_10[1]}
   );
   gpc615_5 gpc2971 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc2972 (
      {stage5_15[6], stage5_15[7], stage5_15[8]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc1163_5 gpc2973 (
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage5_21[0]},
      {stage5_22[0]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1]}
   );
   gpc1343_5 gpc2974 (
      {stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4]},
      {stage5_22[1], stage5_22[2], stage5_22[3]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[1],stage6_20[1]}
   );
   gpc7_3 gpc2975 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], 1'b0},
      {stage6_26[0],stage6_25[0],stage6_24[1]}
   );
   gpc1343_5 gpc2976 (
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1],stage6_25[1]}
   );
   gpc615_5 gpc2977 (
      {stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc135_4 gpc2978 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], 1'b0},
      {stage5_31[0], stage5_31[1], 1'b0},
      {stage5_32[0]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1]}
   );
   gpc135_4 gpc2979 (
      {stage5_32[1], stage5_32[2], 1'b0, 1'b0, 1'b0},
      {stage5_33[0], stage5_33[1], stage5_33[2]},
      {stage5_34[0]},
      {stage6_35[0],stage6_34[0],stage6_33[1],stage6_32[1]}
   );
   gpc117_4 gpc2980 (
      {stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5], stage5_34[6], stage5_34[7]},
      {stage5_35[0]},
      {stage5_36[0]},
      {stage6_37[0],stage6_36[0],stage6_35[1],stage6_34[1]}
   );
   gpc1343_5 gpc2981 (
      {stage5_37[0], stage5_37[1], stage5_37[2]},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3]},
      {stage5_39[0], stage5_39[1], stage5_39[2]},
      {stage5_40[0]},
      {stage6_41[0],stage6_40[0],stage6_39[0],stage6_38[0],stage6_37[1]}
   );
   gpc1423_5 gpc2982 (
      {stage5_39[3], stage5_39[4], 1'b0},
      {stage5_40[1], stage5_40[2]},
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3]},
      {stage5_42[0]},
      {stage6_43[0],stage6_42[0],stage6_41[1],stage6_40[1],stage6_39[1]}
   );
   gpc1343_5 gpc2983 (
      {stage5_42[1], stage5_42[2], stage5_42[3]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3]},
      {stage5_44[0], stage5_44[1], stage5_44[2]},
      {stage5_45[0]},
      {stage6_46[0],stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[1]}
   );
   gpc1343_5 gpc2984 (
      {stage5_46[0], stage5_46[1], 1'b0},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3]},
      {stage5_48[0], stage5_48[1], stage5_48[2]},
      {stage5_49[0]},
      {stage6_50[0],stage6_49[0],stage6_48[0],stage6_47[0],stage6_46[1]}
   );
   gpc223_4 gpc2985 (
      {stage5_48[3], stage5_48[4], stage5_48[5]},
      {1'b0, 1'b0},
      {stage5_50[0], stage5_50[1]},
      {stage6_51[0],stage6_50[1],stage6_49[1],stage6_48[1]}
   );
   gpc223_4 gpc2986 (
      {stage5_51[0], stage5_51[1], stage5_51[2]},
      {stage5_52[0], stage5_52[1]},
      {stage5_53[0], stage5_53[1]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[1]}
   );
   gpc1325_5 gpc2987 (
      {stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5], stage5_52[6]},
      {stage5_53[2], stage5_53[3]},
      {stage5_54[0], stage5_54[1], stage5_54[2]},
      {stage5_55[0]},
      {stage6_56[0],stage6_55[0],stage6_54[1],stage6_53[1],stage6_52[1]}
   );
   gpc1163_5 gpc2988 (
      {stage5_55[1], stage5_55[2], stage5_55[3]},
      {stage5_56[0], stage5_56[1], stage5_56[2], stage5_56[3], stage5_56[4], stage5_56[5]},
      {stage5_57[0]},
      {stage5_58[0]},
      {stage6_59[0],stage6_58[0],stage6_57[0],stage6_56[1],stage6_55[1]}
   );
   gpc1343_5 gpc2989 (
      {stage5_57[1], 1'b0, 1'b0},
      {stage5_58[1], stage5_58[2], stage5_58[3], 1'b0},
      {stage5_59[0], stage5_59[1], stage5_59[2]},
      {stage5_60[0]},
      {stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1],stage6_57[1]}
   );
   gpc1423_5 gpc2990 (
      {stage5_61[0], stage5_61[1], stage5_61[2]},
      {stage5_62[0], stage5_62[1]},
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3]},
      {stage5_64[0]},
      {stage6_65[0],stage6_64[0],stage6_63[0],stage6_62[0],stage6_61[1]}
   );
   gpc135_4 gpc2991 (
      {stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_65[0], stage5_65[1], stage5_65[2]},
      {stage5_66[0]},
      {stage6_67[0],stage6_66[0],stage6_65[1],stage6_64[1]}
   );
   gpc1163_5 gpc2992 (
      {stage5_66[1], 1'b0, 1'b0},
      {stage5_67[0], stage5_67[1], stage5_67[2], 1'b0, 1'b0, 1'b0},
      {stage5_68[0]},
      {stage5_69[0]},
      {stage6_70[0],stage6_69[0],stage6_68[0],stage6_67[1],stage6_66[1]}
   );
   gpc1_1 gpc2993 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc2994 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc2995 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2996 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc2997 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc2998 (
      {stage5_3[3]},
      {stage6_3[1]}
   );
   gpc1_1 gpc2999 (
      {stage5_4[4]},
      {stage6_4[1]}
   );
   gpc1_1 gpc3000 (
      {stage5_5[3]},
      {stage6_5[1]}
   );
   gpc1_1 gpc3001 (
      {stage5_18[1]},
      {stage6_18[1]}
   );
   gpc1_1 gpc3002 (
      {stage5_36[1]},
      {stage6_36[1]}
   );
   gpc1_1 gpc3003 (
      {stage5_44[3]},
      {stage6_44[1]}
   );
   gpc1_1 gpc3004 (
      {stage5_45[1]},
      {stage6_45[1]}
   );
   gpc1_1 gpc3005 (
      {stage5_47[4]},
      {stage6_47[1]}
   );
   gpc1_1 gpc3006 (
      {stage5_60[1]},
      {stage6_60[1]}
   );
   gpc1_1 gpc3007 (
      {stage5_62[2]},
      {stage6_62[1]}
   );
   gpc1_1 gpc3008 (
      {stage5_68[1]},
      {stage6_68[1]}
   );
   gpc1_1 gpc3009 (
      {stage5_70[0]},
      {stage6_70[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    reg [127:0] src32;
    reg [127:0] src33;
    reg [127:0] src34;
    reg [127:0] src35;
    reg [127:0] src36;
    reg [127:0] src37;
    reg [127:0] src38;
    reg [127:0] src39;
    reg [127:0] src40;
    reg [127:0] src41;
    reg [127:0] src42;
    reg [127:0] src43;
    reg [127:0] src44;
    reg [127:0] src45;
    reg [127:0] src46;
    reg [127:0] src47;
    reg [127:0] src48;
    reg [127:0] src49;
    reg [127:0] src50;
    reg [127:0] src51;
    reg [127:0] src52;
    reg [127:0] src53;
    reg [127:0] src54;
    reg [127:0] src55;
    reg [127:0] src56;
    reg [127:0] src57;
    reg [127:0] src58;
    reg [127:0] src59;
    reg [127:0] src60;
    reg [127:0] src61;
    reg [127:0] src62;
    reg [127:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [70:0] srcsum;
    wire [70:0] dstsum;
    wire test;
    compressor_CLA128_64 compressor_CLA128_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha204472099f4fb8437f4f6b4f4cdd2b280ccfcc97b1ef37e0e9f25d9d8bb7de9a8184bcfe059109f2e2d6b61decea6bc796e1f5ab39124787d1bf28f73987eeab83e8a8147f179cca89a79f327793bdc5217a9ee1b73ed1ad38a29cac4d3be11e8e3e9583e8eb76be8cc20538815c8c707f6e6f298274e5e2d9b5ad4d537c338ca5c34f735cf6ede504bda27f56ea8346691c41babbc3eadb42bf68d022f135760fc0e101cc3d660369ca7400d20fcb2fe7c67a40b5dd74f9e83d2fb8c025a579e723b6c10e1c7bd1f6ebf88c48612c44be3e860c074c0e19979f0e0243010107168b2beee79a965eadc5b4f208cffe86bebaff2f203fd1dae868bcf600dd7ecc71d515d8fbaedc8d8d643a6d970b421639737f6355cecfd0dfb82b0424019637d1c4489e024188153361f123b9f9f83084d0c46f7940a4f93e2ca45116c069ceee35638c9cfc356118d6433fa477f9d78dafe42c2082cb8e685e29df6184775f89cc9927f4d5d3360a6430586a4413bfea00461caa98639a32348b7702d189f8f537690b4fd521b13bb32682c1bdb68384d811d81fc9c640413749779151868feea2517efbb8a48530abbbe1aff9a3817b36b3abbcaeb8b06598e543564467580c776c1bd03f58b70e2605b11f6a14bf077442ebf46a03040e9bd514bc6c03e98a29ec2eda002191d4c715dbd9374d840d7a503ac1cb228289f8ab658a76f4d4f862b8874f75babbe41935cb846a8fcd697e9b0ba80c1000a40e7ea5e3990f75b21f8213945390e28d14d768896ce5e4062f7bfd01473dcc2c4c5626515278cb52299aa6a046b9f0fb9e1b1234ff4ffccdefe9f0c08b48d4e65f38f23dab12ecd2621079a096c410fcc25ff8182f1c10b9786767ab9390c1ecb09a55a5ca28f260936f6cd722f4174dcd5540335b9a8436e35d723b78d117474ca6621803d79bb77344b4f0b8e5c57b336eddb7834c71afed2430e891bdd7c89d70593ac529fa72416dc751fa079acd97782096deb8967dc3ded1fba2d5e91136edc479fae22032cf5aa7e855e8c8c141ca2f971027371476cef98a1f19e3e84fb76ce7ff78f524efc355a4b90a5fdc519ce7034b6471117c347c9e95382da211b83f89fb9f2bbbb10d4e2f6ee60bbfd9c53d8c1c168a266982ec4964033bdaedc5726425e016f74eab872118ba2cee23e67329fbfabbf2827b2f78d0ffd0477138c52f2b696fefcc561c64092f5703c59839347f55ce40888e796c127653a1c79d32d1418750b509f7ec2de2fe52d330728b9293255d169864ae128a1e95cdc4a092a31c97e307eb0db140acc172397a2fe0c77d87b34d3475a05d691a35b38e030bf19965362a42ecc6a0ba7143f84b3ed3e5a825e426c15d5036c242f8c1cbc217f0377b5d4eb237b11b9650ba579040546b7d53820690bfffc6134ce9f1e1f6ae41527d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb801f1073a9e48d7086cfdb42312dc0bd830699639a53b09628cf4a8082881b469d990c2453677a9a1d89276ee24e6d401e43b178ad53d9c61329fc8958f74fd28bc1f987b9bb0f5d57721cd5aa3610de232dc8845539efa501ad36c465af6ec99cee8195db40c39e72ede1fab770f33de88ea53b0366f91c0a6dfc655350adfec02976da073847b45c112ef33c8eea2fc93f7f20853b78f4bcb6af3e335d0ff62c1a147237327a84d36adc4be42d7e113ecc7e067cb17f4705abc8e330af5f04025b1224d1baf69a5b64f25acf4b2a86c00c6ad94a88e545175664b98fcf54b8eadec2f792718d8852bf61747012d3142fcf8defe50d13f28550d1da393fab3b9cfa19d8f8d918d63189b4fdd9122f00be697a4d0ea6201d5620c71946ac8fa847c165de5bd68af6ff3327f349fd067bbe0da7d96431ad80306557ce805fc65b61e505718fbc3a3b20c728af0e1bea6ca8c135e50241b7fd67668baf701acda3fac650f1b7f2a329b0355f2150b8656427ad1c0913692b2592f5705e94fe5300a200904e59d6fca8fbdb316fb442e29c81b35cb0b846bd8427ada91535dc1997fe2dfc6c34b56470033f41a927fc7d17d321a3f2f170a7505b0b332ff9728842fc584f4d1070671c093c2a64a4e64ccee8c45f54332dd5e898991c56e82d72bc31950131f3abf6e1a713cac6f14b40d068b56566fafb3d2a2f1fec99be4206594a9b68099965296775ca7d2965ad216d32ee2e46216002c2ef5869bc520748bb0233a989352f43e69a9f6355cb101cbadace52bc03cf77a6e26619c0ddf1563e09360a5d11b3a3111b58ad601d3667f137029226893d8021ec412d5d9643969973ee88d78f4c807dd43fb6020db30cd4cd1fedf8da34c805136d514a9422c06ed8179a1fbe9356d64466abc7af827534cba6410579243506b63624c3f8ae5a49563b0971dc0927c0414947e0555fa9e0dfe67462914ed5a987132a00029292bf20de8177467e59ae29e2ec00ae3625aa4403f5d500b34fed1de437949750543282751f8bfb2b94a049069e7dbd7b1d138a1161d30f0c9db573f8f3e066b6636ffb6eabb07c02cd5800e1c914bd2933dcf9d5737ec220667b80e2c84e74209181a04516d161f3d9ccb2fe0e6a0acf5faad94a779fe46e4d06ced8ff0aaca00f0b27f29e5f84590415b52a698d2aa0d52ef368da336097b1f2af4df66fc87d609fe41369ca3b771cdc88e9e07114ae97b12c959778ede01511bed7c0118996347c1fae11bce89c8546c6b53880adff1b80a21b187f75153f2cf1328e6cb45f252c510845e64395c5cd6f68c0140979db5457c547c2d27cfcdf9619fba14ccf04188099213b26a8f1efc4398faa8417a6d5ef735cac16e110a9c0504f6afe9887c593156c0fa44c8924349de94b4075890a43beaaad5d0b48cce289966b0dec36a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf4e571f75318b60d2f645d9a20726d78b847a77af704a5cbd23912856ee1748eaebff6cc86575850931ce1e39b4447fce829e10a64aef9c916001ac065203f1cce926cdbd7d74e5a1864a4088e55dd30a5a91f75c672374c2084116c737018e9634632268c09e0ef98b52a41e35d3fa8fa3225b5ada7bafd914a56fbedd2fe38ef4031047c271e5d977e1e878c8e233b27b0fb19a73b71b4dfffc2c4fdfacf8947b11343eb7660063e1aa0ca898bc3cf83976260154f263726d748cb74f42f57f5e22c080d5b97e4108ebac60198b54e5a57333b8d2bacdabe0358a71f6d56941260af0e077bc27e83c9052c38cc23d22efa408b4808581cbba20bcec1c001831777c32c8276051b46d57c61a092a03fd72cb4e8684540d289040ab735cdca8a4927acb59c2e8fcbf7b3c1c6f2c58e913d7a8de354398c7cce1956d565c9b80fb319adfdc049ac3e663ffa34cce762d0fe03fe83a6ec8ee98609690ca75c48650b0913c1d803089da1e544bdf35f8073147334f0f820d00e0a055f007395a521cb4e1496f37ffc62609b23d0038db5b602aa2f55f2d94c6944b6f600471f2a4d2a0e2c7d3c5b3dcdfce8eae0b8df91d90187f20d7926bde2afa4d52e82bc2933b68aebbdb9dc59276c7698695ab89ffe0f49dcc15d10e7547b759d3b96bd821573c5dca92900b267b549b4f57f9823ea404c1331d19fe24c2e5b57dc7805755a3b69374dd891c99c19864e2b2d5b9c98c636ae8bd341031081550027b3310536a2cd3402bb8240356bb2d7e05b8b120681f97aa032293e063e61ee7ad2f18513fcfe67a6f84eae0f0e80d2096ca5d7b0a0c043c2249c1f37240573c69a46711a220e06599b83c5e16707d7fa4a431d5453d4cbeecb214cd6a96a9af43294a6acdd281c840aa73de5ea2838231ffe68f8089387394c454bf2b84089d679e662a51fc52d8d5b1ffd3d762220b08ca778f76d5517a3dd5864f9852fe3db64b56acc142c267d565d9239dae8ba79150c598e460d7495e6ef1a7dbd9677f2cd802a909d6747a8021ab5217677f9b350173e36ec821a6ed5f2e8061733b5c2bd877b75ff13be7ea6fcfd6e1b94a0c21ae9de81b3e8a7d3a82de0f3737926570fdacaf095287639820e4f9dfa0c50c067640018116ead86b30dce3b2e652ec51b0e065a2e6ada52344f040c28ec00887399a0c722db00e17d40a568fb5a4e8fb9e9fc76c6d9884075b2115f69c47e39038bd752d77f76fd84dd2e986f866f80b5435c926b15807edd2b3b6de0439129284d7f4c90adca4f07a071127d3c09a05b400aa3a71abd44b5d3059031679c8d68e8c5103cdae6e0de10416cfaf5fabaf82e915bb6985c5c10903c80b05f09f0b2f38b9f088aaff7d3abb0b54dc699c8ee9e2b015b70b907d3213645f291af0fbd70d4f66d1057ba12557ad811677927ae5b605a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1f1ae1b2a4b53c9a82d711e1b88825e945d8d672611cabc545fbb7610367aabe998e995bc84f24bf3cfada7e8c33579eab2326af23677c4cad279c7360b7dfe3e574952231a11122b921a5b767e33910c5d5e49d52c5de5076aa5b9773eb5774619373b2ce48ce7d45dee9f7937fc8d14f85fd590ddcecaa0c4eccc90ed44b75bed161099eb79d05f5e496f8ee74972e9dd5547ae97bd6bf2aa39de99cceb44cfe95b5d3cf6238bc0954e2464fa4b959163a1050e64c2c1059225fa26b41ad7993dd45c23c69e48bb4a42d45516107a29bc2ec3491d571a835f4aa18617ef5bff73e25c8a45d79a479ddaf6f07ad8e0263a3771faa455179a8bc1f610704420c3afec8a2e530a35ed706f17c3799e63e5424c4aaebb23a422926e6be1321e0553979479ced24c9edec8658bd482d7a2fcbbb4a88884064c75a8e75d1eae8674bb93a314d9fe78d91caaf3e67cc40b8abb0084e057aa966c17750f6879d3cc15c287a3ebd1834c93059b613b6cf2d19d848ed910da4bb1f95d31678751715a5d42378f0712010eff5fdd3bddaca949fa397e5d496df3d402e7ce2ede097d3d0aca39ceebefa5b4b57bc4a361007578bf7d2ffb8d49e3af68a5bde89ab4ba4b218057e8934606a7c8a7282d4c1336272339bdf8cc6e656e58447d25215a2436ab600f55c623690b47648c6b1d3415133c449b23fc37b63468a30c3159754e5790715aecf99198e08dcb4828cabc487d7fa27b35c2c9f25ba0e13bdfad8ef04ca3aff96191b37a9e2410425cccffe870e62d984f9276ffe98ba35b3460678c115f943db052731690b0a44207d41b3fab1af6194970a5e4d26eaa777aace4a641a1045e67c488297e471a29ff39341a813c62a3c50469f09ec937ed0de4c3ea943b270f9c5c58195b6b6297231c77e45af92959cfcb7658c780bcec0e975e671d591d0975d91376323f8bd7ea4b02feb1bd507d7e95fdeb07edc4cd1ec11b3b02e267a3f8c80cde7c265dd585762ff072215f923b3ef1fe1fd70f7202a1dfbdda66ef69c37799c576cab544c8024798716d1bc763cc641e7925cc420124ead66546d4d4930dfce2f045266e1bf2720b36ba87a4b3a434c8958e7b79027c542235d93da28a66fe50925f9918d2f2cd171c4b7f64fee2afc1bead1c3b1a1d26c067cfbc969504684e806a783eb417bac4ce5df4747dc89587983f6c16875416311b2dd3ecbad2fab6fbd9649bbf53e1b76e1f72610178f3aaa803273fd41cc6004e21600a7b04a1d66ead6c7a5e5b9b4b6e1a2481581c0fd1e3ea8ac684ed5485c77809c49661f95d54566d172bedd7ac208278bcf67c5aca73cdfce83cf6aba58c0576572c93686e4b1dd1e3247e5592a7b58ab5379b11055cd892ab642eeca53fc8c0d36c65254e0e3b0f103de4926fdddbff2d7d1bd78a1276acd66911744b932bf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52714a8d1511e30e8d57068a031a61217fac4f7b62174dfcea8512d52570f7ab6968d055cb33109adb2f1da29e0934c543d43685880122e7d4318b365c4bf8bdec1522f51ade34c6563cae13a508bea3c0c4976162b0cc80ef0ffda59aaba0e179dfa700924fe904f330ae5814ef4c8c2a06aacac6877065282e9a40f5f28b68167c4c6f6c34a4a4f1c5dbecfd91d6fbff1fed829f5854998c58e26ee80bd5ffa3a343194658110f9d9dd5e7c4bb820357c86d3c9f05560154cb7610b3d5113a1f6ddc4209f320c9b260467583369c7d72345a23a8db32e83995943375fa4eb78f46e253daa18607190d18c8d7d2d240ba261c5f52c417cf20f1bd95fd2cd44ddf2a89eb5e6dd198d29f1c037cff11e432da9afab5e8ccf3ce7eeefeab62f437fdecdafe10e7e49bf1ea1b0ca8ba4a49f7f583e532e39c33a6789c8acde6ebf8df8c5b24837e46e3534d985d2d55791d07b84d5a046c4c21c8d8e3318fd0c3d90e908adc77cc45bc17df9a8f2a631d88dc5fe8fe848f42acf36bda77c0a160c014654796a4e825bc5b68bc2eb9cc1fcd51c0a7565b8cbe5be703e2969dac8fe27f24b8df3dcd47b00fbc5e7c876a0bbb2ac14c70554894b8523fb35e0527e6a68c023fce0f17c46c3b35c4c31d5d1df6284b2db7b895bc7ee52c677ec6bfdd5aaf7b57afc8ee276cd7049f86389b74afc529cd92438fefcb1c163d0b0afef6b141f86e37ad2764bf3b8aa1fbb17279d7d406d5d841998fe9a8d8af6f284ed4dbee11022a2be7593868035e9ea4b4e4479a7e96493667a92ecacdcde7c44f3ba480a4cd5b07c387bd9312a1cc4ec28bfc0b9c3816e58b57b4dff4dd40b376e29ddc7151e8e5d9f9a109587b8341bb98739f1dc577f18b5922f4788a75fb85309f0f9272ee6fd728e1f0518dcc8fcc5767695f7857651db7ba45732b9dd44758540cf79c11eb5b66b7074adb0f837c843043e209523b2fcf68af047c13b56652fb13435f9970ee34420c625684367a75523561ac6f38fff3d5311b323ef447280a8079c071131830ca1f0cbebade26f531b0ac5cfe1d9d76b85d8fae0785b914b3da68395be8021254fb991d340c172a10c30c064e060a7f726d6a10eb60fdbef72aa644330d3e3e36f9536ecf7f07ba9a79922a5eae71cf790dbeda0eb56bdb9b28014f7d6ada047bd977757ade82469ada42d9a40e96f4f7b1c83853e2079555c5202f0a54d32150c8d9b66de0eecc85bbc98ed98c41c6384bb79d4e029399184b04d532ae4d2f993cfc10e1d1f03b90516a0c375ddd3634f941bbb7d5cf38390663c10c676b0d63571cf74214c52ec96d94d2b8415dcb1a108511d2e167b21947e955f99ad31400b7166846cb207e6fffbe98d67db0ddce70cbf5e819af3fd7c165d21de4843cf8e666346f0b71e6103b628711062344a355c02e6ce4b5c733;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf8f36452cfd747b2f668387dcffc4df1cccd6b0090dc771b277d5d42967ec3f12cb59b1c75c2761e8d092128dc3bf9e6d83122c74f86c7828a376cc02fd481b43fed77c6d6355ed26a0bb71ac48e686cfe26aecbaf598c987025f319056de03b8251c96b5cc020869b2026a60c3948d11ac664323ba6c0c61ad29084ff373aed0119157b19864ffa6fe69ecd17c95b6af0aa16bfd362cc4b75b438c3948a39034015df90fa4e889de7c41b8578eb914c2460b50107249bb5c76795b67c6dc507a09e0253636c93c63111dc5122926cb57289056d66fcc6f9998d67d5f68fe8dcb5eed75b689c2fb22b8aa8a68263b886a81d255cc2869a829250ccb38e829595dd1c7d2b0845a815852817a3d82978cb7c81b69ff62d3a25a497b93e339d5624b2f8d6330306ed46e9208a8afd3c7e6091905a50ec8621b5b7185e0701bbaabf8522a3f7416fecc8ce1007b09bc13be1a8267ff377584dd90921c6419db7c4a36aed25db4f00d92469f1eae725d95b3a7884fc5c5eb908cf58559dc8ef498d040647961e3a4285549aaa2ad2e6d6b97b1fb859486ab0e18a4e5e753d98f2743236ce98316d423d7a084b4d461a9c976bcb7e3d2ddd8f484ac258b20d962c6c72de8ed8618e7a46c6afd53f8a7b5866543fb0e9ecb53633482b8f3155accfebde15b1c323b5b18c127f9b624d29aaa823b6c55fd52d921e8c9776bc90784d28c70c598ad0584fe9485ff6c3fb1a520bd043cf4fde77aa785e94f82568c4e5a9084e0e1a978efb1d3e895687995fa14404a347d4445a99f54460db3bb19fc656dcdab8e5c8d198bb29723beea3305398486af7a597517b3c52483fcf9a9a3e031a6b26b86372b1d9cf9d4bb0223470fdc19668f288bb5a5c7970850e9dc6f1ece3481b3807418e1f896b74b3bdba8de75194edfd0058f40df81ab70f42da60aa370530d4fd70229a4bbfe7dfbbd0c0abf1725f829b8023cef41ad930ec21a074622ef3deeceaa3c5ddd8c6766f774fa2a415b6d5f8dd3734bb4f2c99aea8813d1468d60516daff55c02593730bd49493333cc8f56f2bbac917bd9bdcae67538dc05f19e445e9cfea31a13716c1f1c0ce7179a24c0b1016f07e65654063367caa7893f49f0f955a9c612638259eaf1dbb9974bfceecff4deb68920366e0b3ac50df50ed1e85c4fe0b05acf3455136a8f2b4ede11b8ea557e0dd8ab6352eccbf4ae844371be59757049300dc77006cb450bef0c576f02990e56c8e02c0d5b2439748cbd9147cbdbc0fbe300b8f0c435763399d97498c42be5970ea2eed39a454676ef63f32d3ea3649a53fb0c59325a70659d60cf214a06657a96b919aaa7227202b8835df1f80a39bad0b7102c30b8ac276afbf85a3492e044c449711939b9168700cd0b47f54b21d91068bef6b891781d08971c7314ef637ee9998960f97d72d2a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5ba8a85c84b190ffce67f37d75ea2e09322f1735ec94e3710c8f929814f50d05788960bd54d892d411c64ce82e7e003df494c9bdea8e697f57711512a056c8d7ff94b5b13e06a45b8fb2db5d636e20c95a9d2fd09a3ce303f5c42a1ef7a75e68934aeb71902f7397327302802b45950d7821dfa13362f6eceb4c8bc1013519e15a0919b74cadc78fe80deaab9a678ac53d2da9b03a5fea7d9177e94a1ab5b9b27e239f09eede8d41493871a53593577d9e1949299847c5fa5f878e92e82059462056472d0dc2794af43ce3bbd740ea9b44dcf7e418514b981a92f0115d6044a700361f14ed2afdb52ef97b96c87e7aa61e6ad293220d758d7e71945fa61ad10157a138cdd3b0e0542864a2940adef28920c2d0ab231e5b28711c0bfd188b0d7772e66df19e77fe9e2e9759f1c679621503eabf9396d5df557196ae04bc0f8934d9aa0b50946911f00378d6bf24e281de549c80f281a0c537dd723cb6d1331bdfe9299b761778d4585a7bfaa15433bce2b151a68fd940f9a1fafc07f77f48a34bbe962737245c5326cc33a4da25b704749d51a96978e78ca9a265a6090398d7fb5f97880e73c87f8d9604f85ffbc3ee8cb3670963b8ab72166998cf0685fb2538d99f6d8ef2477bd85bf0e2d87f8e70d5b2d0bf7156295962d6b9a17183b90a3534471deb89af3e5d6da92f32cf0de9e810d3dcbccbd6f421978c8ed959087961e9b87fb951f0428bf3a1b76e4f0c6a24cd8ae192628928ad6eb274f402b6cc12ce44e05d2ca0cfc0fe1ec1ab82936ae60a3ed6b8377fea140e372f29bb495f2ee19b3305edbf1b63ee0af244067f156e76b74821cdf834881bc0d85c29082b5085d9ab169ae368f90dc587da00452c430c805cb8dadba2348403472fa82d9ed001bc6b9ae8c35d373fb8c7de15af27f149a2ac888ce8b067104e4071bab2b85853b423d5ecd995ea31002bc22f18f92a37f5ee110eb955b4da426cffd3dc4c3f58f73f4c03aab618ab8153ee30a4e50c836057538cf7f3fc39deb95d09c59d8b7de0504f115f1aba93169d7e89c864a2b93731031ec3865d43d56e3dfa424822e1033b065254422f529690ebfac363a87c54cb20bd4a0275d56bf9dd77e66ec7d11a452f1a80b3865b94a21b7a812be5a19533fc986d2bc1d2aea83e2ae0bf30327f73b36dd8b4bc65a982d8b6845ef112f6c89661e0938c03c870cf2535ebde2ad150cacc2369801213402bed3f0fb824d2fbd4225f1998bd605d5cab5d92ceeda6751f150a14a1273136961c5c81d41c2231736a2d7058ed1037d0d33484e71ae2ef22400b04a956e6125ad62863b17249992a8a91544e46d24d276f3e903c857f16603d1167c744c43b9f9b76ce54c15952427ca349573d0fed7ce4e1da346f47ed912412a1275f381063795a8abb397f6f2f8549a563643e7384acfdc67f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1c6e91e8dcb69984dce402a50cfd47b9ec9b418852d81ced81b8b6be227869444cac69e56a67bba252b345f52d10e07ac94f0a671fbc08b5b7c01a8a28a19c2763e1718c2983e73cf5be831ce90dbd24cde6428aee9804992b4d11dae8c0b62d62fb026f4139b4a3211231ed4b867714cde2b0ab8a4bad4ea3c693f8c98578b8f9f4a2a1d1f90247d54d7f3bfbb1d68b0e30a45048de1f100792751c984136e727f8d461566160f98026831b7f52e094aede64416cc0b9038e2e11b8add97aecb37131b3338e45e62f157c9435ab7da6a8f14226703f733e604a4fc821a84a62f0226eb623629f7a955aa36893e6f855253a1ef4a3a90caed96b26cf602902a8289b10f07ed8e90e4d385e797f0d90c893896b0f82947f5c8fecd448e198e39aa0c962eb1a3e20e4ec5c93222261596bd4356001ee22dc31057918ed2b16edd88e75c095d29ab7409d4fdbc3db8dc26e1912dd19d248d92b72fe5ae6f3ac3eacca81d13c9d9a8fc21a820cd3773694f3b7b4423c429f2f614e42e31a403f7d96b909b51b19474f5f1b9c382f728832db8ead258c32e65cd32d5a95586cfa6fc677211e1174ca05b8ffd1b8f72b7c4d4b716bba51d524c525731195bef031bdc6511d20eb6fd942b3d3b4dd9def346d57d2803b62eedf94237c2b7ec0a49682de684c524a3e7f746194a26147354fc545b37f640378fffa59725c0ad4ee0f47b95c3906495d16cbfb78b826c23e1cf2576728de911575778f204807fad92b465a89dd002332eaa4543d88a89209b37535edf93249bebb1985a699e6c5d5def9c8eb5fe81acee5e9b276d41fdf3545bc1f0418cbd81849cf6c6e9619396cdb6e332bc4e7a8ba1df719df09b3398e3187e3dbc40c45fa54d51da5bd814cc83249d17dd84e81d56dd50fd363e0fcb077a205268e96031a45ef569a4dcd91842cf653d7cf193e22f221e8604836960f4dc2b4b8b076bac2b9e2597289aec2d13ffd58016e7c3176020dda54c7ed119533a9f91447560c1c8fe4ec3db9e6c9b0e3063f157c8cdf6aa87e9f9b0f90aeb6d6c6c00af35862f4b258b2fce558c55fb81576bea83f3447922ed775808fd8326150e2aceec6d54c71ccbb1cbf1c2177d4c17170ece4278f15bd8f59c7f87f3363f62fac217126e3c591ae3b847d5c10c6ac19d9f8b6d29f1c4794848f1175f68d0c2899f1e6066593455fcc1cc16226c684f169452c8556b3b6b18a35fe7a57a1e2b2bca5b72a69f1b41fd1acac5fa85fa017304253525ee5576d6fda0500492b536dc6410ffdc653a9fd857862b9b4ade460df6f887fdfe168a061900abe94a471a5875770b5e6d24492803ecc9f72f2a9b7701c3001da32b5db884dc167b60fe34a23140d368ead33b2beedc8f63cb820f9380d8ff65bef5a5010339b8e8d1cb3052d976f6aabc126483291fd92fdb2d6b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heff453867008e2ec653334c018441594970d7a96dbb494327fcf8790cc222b25d6d3c2ea2ad9be4cc1333caef76dfd25b60764a4957ae1ca240a93ed864029cb5a598c65e90babdecfe88663bb1e93f41b2f73b32cbc72141b7eec09e05ed7c8dfdf814b0ce046cf9f72748655f12a9b3b6fe222b052acb6de2290bcbe2b76b90504073ace25630365e700c99550c35ae88e7ecd1145486546222fe342aa2be7b53334cdc17ddccd1e1d87abaff4db153c6685f84e6884fed0f2ee38941ca16b8392d3d3560c67d8df22bb273607d3940f6b95c3c42b04b611d1f85bf59e1e27fccb601b638718ee0ac81e58ec6bafa51894b194b35bf3e6e1d3e2f7cc6ac105ad1360af74a32932e19ebefaf9d36c780e65268b6bd351503bb33f9d60c2acdfd919fa5c0d62b9687299087fc4a74973a04b09dc7a4c8f3c19508f55a95baf09249f347fbcb1631ef79a04a92c0bc2c882502998a7395a46cb358537a9c57a4267da9f051c96c62b3854183064a38cf7e5993a6919124e0c4b23179698107e03b06126cf595b525ebfcdb5afe0a069c7a1d4399893b4726b647c4f611cd917dedff29ce3c650998ea6eb9b1f50942e8151c27ff00b93667d2fc69f72e1d4fe55522151f33a1925c79d81b26777f9737019822b38dae801f0227838a0232c40db8f8fb432c2612c1b1d7e90bc9a92ed2b4eb3cc7d36880f7be4038d1c6ae62e08b75b2fecb8a9d50d6344270b6ac8a2dd37e4cbaa37bcc9ebe12e5fa042660a0df626e4094c4ac6f274661e8c82e5f189d10afe646fb0763b775750a381267f01c25cb9daa1ee9f2b5e8401a437bfcb5101f317d318d4d00ce9cf9d92dca0f825baaef1b0df5561748f2cd5c9254762acf56a1b518543fdf37e7e57e70945beb935b24c3ee9f915ece2fe769efa9fe320e87ac8a00e315b2856027464baf078371da425d6ca282a00ec59bcca7cef25e7a4d9b4f43a4075a348929702ee6ce26a3dc40e87d887117678d402087115d98bcf951f1c0f1a50a4c08c34c13f33b12b44b9ec084049817f8d6652091218aec4786c56e90d3b667f8e24e8f5f4efce1f02583a756056b692891bd9c0003fd05771fbe77ae559fd42136af951a8bcc03498effb2da53e70129432354afa912536cc0b93b423518906be23ac77c8f4e5b8cbdf60bc92900d0463e2bdd25d307fc757c6dda98d0337cedd5d23e9895b5e66a54fd5740cf5bed26f52762032b1085500dc355e81b903096924dd426e8e2c801a1c806d82bb315e35f68f3555571c185b71a5469ee46f19d0644183337d5b21fccf601db2ae6e4c9818494a73bc8c324dbbb2b89c29f79c34da08ede6486581fa7534b73a5275f0f8cf724f1d48a35b89758820dfaee5a6c7cca0eaf2630a3f82d37cf9267ee9a1503139f7c4090a574a69fdd02d73e40e7a8d702758564252;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcb6ae6c5798439be994be5b83060012443cf4fcb04aae6aeb11abcadf53119a218f211dc8ecb5b392fd4882a3d84df5a6283f025fb3563a44f9958ef95aefc7003b09a1788b7fad950540a4b262ea6bbd48fc881de0f204f4865580f2446fc9c25bd3b475d256b40eac698ba6feb84024321353a2b773efb730732f8243610bfb7d5e59ea7db77dadd16f54afe22d6c3049602a40d261755f209c473c923c405ab61323618d5585391ee33a20b19136daffc8afdb70e6d5cdd2ce47460994e934e7cda09c429a189410c4117fa6426c66aab00013410724c4012d305d997dee4cf38056bd34a6779e9d33940a36d23d1cb8b280d9df2e17d5d37405f1dd4a498d40e1d88c0f63a4731adce73c769263f60869dc664f00ff69aef474d0c7a02006a854aed2099d6c26d1543e01e72dc246f8d435d05bce7d672d17d6f7219f92d5c7b4538b1cc97243d48c8f562c7ad949537f05c7d3133e799dafcb2448de31d823038c9fae001e0606fefc0d9dfc2b288c8d613e51e1f530ddd10bcf06ee2f0b62e3051cac7bbd001941cdd7087a363d04b24d18bcfef56f2c6e5c57414c61053d08b269b4fe39a14ceb2d376695de818b008910175b56638833d0a588e2b6c6069e5bc4793433562082958a2b6ec597e671e7b4312c6191e4715013540f69fce0842a84328331639f0d81fd080533cb2581c506d510d02307891f81c1a3848990887faf567e002c968682936aa2295d6f5bc3e48921fa65157d2224d0dd045826c3c8bed156038b09d471367fecc3dfc4c209048b0e067f26ccc3f55be0f1d93eff3db65808c53946ee2be1e288c6a9b14940be862f85589c0ca6fd376ab9d61d01b4091370a662ee47e4996d86302433ea834232980265d191cd9acc93d431f64a919f6cf03b8a5df7d50de0acc08b1c9a2235a8f7ad08c0f997aab2a90105bfea41a59f6b512cf21c163f378e70e4d8cc73df0bba850d4e03da8a598f18c682ecc6ea092893dd53dca6dcdbf813326bd006929407201dd1a5569b5e6b62bc5be34ca4b6cc33ccb90c7dabd99b3379bdd4580067d7f87de4d63c871e21c4a71e9dd699083847e5c2605276fb18f050976418751b4072481bd18716fc35f55f6770acc3e76ee99af18e96939845456cdf967ce1b0dfc635a138ca47e68aad2a5228761e6c07f5c5b1a627c687cecaccb3e8ec6195befed116ab2275cbd2107920e7e2c86fb2d09b85984b4d5f840b1c27e4acf83bf2d7710d692c531858396911034449ebac86a16213e9570e01bab06f798fbc3b737cc3251de8340e1b263e41431ade9a31b667df0a8a6ef415fa80ef9c1c6dba29c3f8f404862b27bd968a0993bed488c94cb6f278b543a353dc6abef87a9e42ba03dfdb3ec2f37a79b7a17ca179cdd8dd666c29a4b48e2681d81e99028c32e86c50e118c21c822285fb0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h69ad26db01d406bd5a52e158c7c3b7fd8abdbd42ff6e5ff43360547631ad1fa76890aa94ddb427c058602246b52a2bf4f40b71d3dc2ee58a1a55052befd94660bf451b3817ec2808c6cb4926db08e66df9a78bfa9e0a21422a552ebfacac3c231790bd0c5ad57d7a98ef7fd91c6e1f90a9cc3d44979b0dca97b38022be6db19ef37b4956671cefc08659d443e0203f236cd6513fe3fde31afb7f32a9d5445a84e59afde5d27cba5d3cf0e17f518c42478f9c1eb7cb40904a60a46a6ca9dac147432fe804128f93afeba0f4777e027c652f7867c86b24355d86b669cf74d535e3a8fd0d661cd40476f7b6e6d3f9c816cbc26932667b0fb19f348ab86ee67a0c9a95e763663882ec788bbe11d6fab957c98300eb135cc91768453d4f8fd4a6343ae8b35cc408b8fc3d1f31b53414be27ea463173457921f11c3e8556df5ce64a0a878a7b277ed6ea1d81f25f0cf256466cfcfaaabcb4d159f6519bdeef8604cea865dd28001202318fc6bb7a8c737271d6302702f55d0cad0d1c38c6cc46b933468e5955e765bd92b5c97a487249df9d582895170338fcc07db6f89c3e44c4bff942fa369574a9614d62b6f20b236fecf855e8f396ce8848ba1c0fcb1943b2c94f2352f24918a26501b7375ec4d2f8b6a95aa4eddc3c4979416b97220f7e049d9447a83f284d89b9ea291b281838a2ce2bdd731c2434e6603d95f565892658f0d5735218eefd9903405ebed8ec21b7485d4e7cae59c3ec50d0864ccc05f45dc56959272c86a3b3445297f76c9ab408d2161fde9c0b7e673da2a1723d1000ddf5c35347862251d346c29d853d60ea52758099b12e74f0dcc8617876468487606c701b564061e44516b40a995198a7354fff53ca9956bd9f18319fe1fb9f96dd662f8de87837bd7b37cedd8483fc656fb13cd48a78c149639c215a192a823b17327d099cb1d7d5b1665dbb082bb51e0badfa1b8f545f3d2fb371d75f4a3b6097c358e1416a9fa8936c480bc1eff3974e800adbf55653b14ceeb098ecfbeee0b3715b9dee24e0413760e55d922bc9bc3f9539035d81109f6ef0b3fc240a97a591b393ecd6f432f59d038d928fdf15366196a3187deff6d699f74027d46476ac18f80f7da159e69823347e30bb855321886ddb0218fb7516c36c559add8deb40f9984e78d87bca73d8cc8203a8551d5919f5f9103e18dbc4aaead4f6319b11f9d4071063aa9ef0d41539489cab407298c15cfe8f81d90fbc84769d54f2e507b3f62f3a2a91be815a72acdb5ff9f0e7a3d0a2482f6892da531f5d526908977b74ab67276d4805772c601038e175bc74ce331d506f52cbaf6777d8c24d618a4ed251f6c407ce150a0d50f1a49f813497392d2f8ea848d8efc2838b656dfe93041a9827663449b5f6f3d5a861bc3a6fef9f7ffc350ab20256c3f4941c41f70436f169399d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8507e2955d03b433141dc6b9575f7c240f9938dd39777b82c3ead3fdbb825f566971894ed3fcb81b96b8a0feedb70cd6127afa62fc3a0c0624c07d6c473ff3d78f93be3be896ee297c27ca4fee6c8c3ae4f60b634d9a3471dd6fe8408445bc09e863b5919e25ec4fdb4fc59a5ec2acc6678e470868e3507be3921e35db987f2f97fd4e9fa5f4fe2292337f91afbe3d195d4bbcec3494e132de9ebae73cf0a23f21f86c46c13ab276231a5bb7e65472c7591caa2c8b8f198d2604333299229e4f8f44a633bf7cea3637df0f1c6f35af247277523b39829abb1457a0b86590548a6366cbc2dfd7ce02ae87557bc37a8d898db1aed510ad6bbb8b5e9bfe5baf9f4337e92f9033f9fed4345013ebb2d4706bbe1dc274ff37324081e828d7ff59447797c916909857bdaf2d892f1b5c3efe07c0dca608736fc0f5d6d537127c24447ea3805d731b60fbd07ddaaab033b4a7308912af895a0f3ec2862dd4e6a6837f8e0beb7569ccce574c5dae6bccb1a86cde7c9f4ea0b0af71b85f62511c8a5a46960832e465688d631d738b08dc04ea7e34ed747febce58f111ff46fbe9e49db970e94a30b789b666d6a667d84409421cda3e17dd60b307596a2298ec0d597fcadf719b81daf5a930eb66e8c34abe5953543945c23aa50b3ea5415eb360ab9a82cabe675a222e37aa4c0723ead9383498174528018f9d152ac0067a0c9a176aa675c9f3ddb2098e015c016d9a0611d01313f43122b1a3d24b32432f0acc91b0da22715c57aa1dc9af799fff0e9aa43b97e83777854c801cbdd32f32871cfc035cba1930ce9b2656d1973ee493d1daa1b97d27b4ecb3404bd4f08d8afa6658152146dc92cf90433d946302f10a7c56645dcb61f623ef726003260c39b9c5986ac7c3b33e2e5eff87389bfc2d0333a005ad8e222e34a449d2928def40cada52c24a576af4b5669f18888f7c391150ff973ff18608c290c0476f978bbd18785a48821753a4e4d474ab3aefde0521039e07138e0837b020d88d2607358c7e465d0b9f290ca89eaaef88f6cab0098653385955a6cc45f6bf94b26134c6c7a3ea3e8957464d35fae002ed6f27ff401e310b44d79e5baaebfc78c2fa2cc65908d89e15befe6f09f1f97b3c9620a5937946a468d480712f713a6f12b43714c0b443e1fc6cc5f887c4ba2b550c943cc6821ed89ca80b9a08d32bd726e23339ac4bfe84d02cd39f7b1833c0e29395828790d790596580be492dc87c8ed4cccebe6284fc8f7c2da55b338793916b819b703ebc3fc97a7ba882584699818ab9e6b7124464e49f2a0190cc9f25ab605eeb41b3170565ec65dd6b16f67e43b6e735eb4ad4f84c714828aa6ad333950e375e6adc615be1c0c5616e2e6d287e4437236356ec0d3c7e35daffd518eced9e7f0b751bc4bdd8c6be7f630ae54ab041e60df2b202aa0ba497;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4b53e018f1444701748f8822725d71f83aa8b90affbf38c1c304e24cc1abd4ca0d41d7d57af236586a2ab49f705dbb09546ad874e3ca632211b819c0942e15724623c6450a9aa0242d47b6271a7dc0faabcc91ec0d60e9a724624b04506fddd15b1dcd3731617551a4d919630d43639f81589d1c2637c6805ea33bbf45e457bd73fa629d02f0e7a07afaa27fe58f4c4cb9ee49a7f752e1223bc7ff6967bdc04e17343a7f44320ebbd97f533ee434045f3cc1a5fe332e0acc855d03111e7f290881253b24966090831bb4f17f1dfaa9c6bafb8ca4b682efb670b8ab1d6705797f5ddfca0b005af12ba1b3c4dbafa6813b05d13734d6ded64c60c16f25d201b2c83bd5523c0d2d060256af2eeb61d2998d114e3325eae5d4b2704cabcef6a12647dc73c895d03544f5148260309f038cea74a0628695d75f2d632398f82f0c8a40684ffe05d3c52a1e45675a0d519d53b6bdeb2d228410fcb134bfaa20a2fb7dfd73156fa5ece2f06e540a4436d5830d7e898a0ff06d452b07c8116ef2293c0c15cc82c06d8a9dfed78147159af07e7e6c4aa6ba7752f8182454189a7b0affa26f231b3cc0f823010ef6ba1b2a835ebb74b1c499b003edbc20c7141df8a264e46f80b7d435d621ca88c397384239e1002286786d59e45bf8f4a48be3a66e50736b2e0943e6271263ac5a49db532f8fa56b3c500c402cd08560799c5a6050c039f3e6dda8c6933dd2caf4f759eabf8c2e11abeaabba3b9faf8246f5dafab618d84a8e328bba5edca4897ff478b190af61bbda673d788fdac746bf71f25c179be1d3fa857b28c07af6399507ef40551ed2de2306e439e535d74e0f02ef0e0608ebdd875a295b2e7f5a0ec66d71eb0e6370a362bb665a08f51d174acb3c1abfbfbd444720abde1148c5c161ffc2061eeb6c312226967adb6c19ef4031415e1aef60619b7299e84d1a820fd51a1d5c9239579577ec003f4d93ee9a30a3b53a03a2be5f959f823f6c44d21e97a17beaa4a68d92a39df85f4963830d18676b234cc693f8f5127604d47a7242637b163d7bcf1e62ef65e1acdc5b607c6ffa938a0d6bc435ae2cd2fb3b77aedd0242eda97dab398902a625a120969e43f167ee2801e24397a11976c4ad1a91bfe8360d96da81486f32082407ba8a0e7bed5fd2b9965fc757dbb46191905e5358137059f88af1ef673efebd56a0b6b9fb044a799ed882fcf37b83af828559410336df05625dddc329ed9c101a21c686e7451388b281cd9b7a89e98244c38e9ab02f29c7b8289e542e5022589c8e1347ddfb6b2bbb33ee37c6203b03adfe0589c7dad6d2ef95217e241ecb8ba3a88a353404fb81c168b42207f68ae2dd239e80c14a11eb41f4cb9d7ddd4508a961967c3b48870f9024dcf0f2dcd5caaba12dc64f2d953885f6a3fe8d3097b32e1b88d708ccac0a0a9c6e018e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h63cfeb909d9a66e900ab4a184a248c6df0e6b435a276b176a25087120b9711912ecee68d31b63ca369e9deeb68fc564f67ae9801aeeb5d2847f50a455e8079436c73e43c37d4b5838be194183b00d89a725fbeca9d5710fdbb60ff54e8583e7c99215a901cfa09de08e6852df5e8b929b1d07d7a512faaf4ce95279aac7190444e96bd4efe52209317d2ba40c2ef9377d6d58bb9c3fb826a25819a06db55391e16cf7157b9bc71ba21a7fb2f820c2a091ea8241ba2f378eca34fcfb7680014824c971945b2bcf226e8f270c64153ffa3f36da1fa19e888e53f5657222fad4535f32385e82b048742f5cab68b7003d020331507368d2822688bbcd986fd80ed7516ada26004a939c7ee54c2023e3a536fb7331ef6e1509f7dac797a22b60f172b7238f8fdff6c8712dabe6094846809dd3c34d696434ddf2c52b01b50c20b0ece0279d100666d4aceae941ccdc1949aac727eac2b001afd41b614eb9eecef2444acf065ccf8c959c7a1a5ae543b3c34e9be8bd049501032dd2d3898830334cf7c2e77eead5dceb2f3b5d41cdea5e7ebb638fe0a82e5aed89a49897eb4f6217fe46f42bcf4a2e0e41859ab36f7fcc183de924c697cadaa6f52d006155cab3274c7ac6c8931fa9dec6ab17dce001d1b43dbc67c486232414de3eb5e667aa872c1f9705b5a472bed2a18688c50781b4499735bcc66d631d79f0ce30f7010899107c2f50e74ba1b628efc655937ac811100e26c39f4d31b1c9f2ac9cec02babced627a31f215795781ce7bc932d916ddccaf678d464e3a85fdb6452c63104da0d2e5d1d9f76e5b662f3b4d6c29b3dc9f2f11f4c636bc4a282733b34a14faa55429d7e5e83999e9cf19063cf14e00f32a0af53e957df43aa3b065b653752daa0ca25a139d30dc2500b7cf0c6bd5cb04d83bc07a3e8b4c09f889817cc67d72c7001cea97ee3e6fdbb8d8d5a6b9a5edb7d84b05560a3a1dc0b8a02f0b68769104ba7d84bf0bc90752ccf84f5a399b230d4a7e0218b1f14cd1278614b8cf4515347a8fe6735dc6882018ec7ea05cbe43d546068987ede539e264c399066a531172a97e924fea07a30b41f33417fea5c229eb8c40b5eea7e067309f09e966a2d68d0aacdd10ff1186d199c07b694f2d1000f198a9a94c17bce7498d2f0e32c6ac55e8ec6b0bda8cd160211f3d85c79cc00b848318cd051dfe1c33bd52b66cef266dc6dbd34773af74db2786deb01d14561ab4bccb8a694ffecd259a830c83ffb4a2689a980e0627405cc936224d82c377596b424dbc5860a7b860970b9c2760da78787ba24f69b207c1281f08e26c01178c2aa0fa72ee4072c4a105e4a73ac73cf013d010592dcc3eddf8363d5e4354eccec4dd6f8076afe2ed30a4f7c11a5811daeda30fdfc49259d8bd1810b1ef81403782122b3f9b69c4ea8da16cc7679e1735fd16776;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8bf116664373ed1fbc5c60e0638625f8c24dd1e9fab544b47991f5effe070b4de4a5a13cc97d234fe3e52f285e11689c64f266d5baea2d8842242f3b157806e11366d4d4d0adc4718d50671357625fbcd2e0cef46c04fd455294bc7cd394291b7049ec3d06729524b977807f1b31ea8a50b78fd83e7476c088d896057d985f17501d0f4777359f1111a03568268439bf9b0e6eb20c461d576fcf1fe7f75fff652535f83b3341098a1b9b6cb84c8ba59cf264a3c8ea697f1534a49697f39deee9cc4990a6f93f742077573ad090bd635916f5632eccf4089102e6ac7052dd78b66689e7922a46fdba0dba3f80d871d69576168a606dc479f75b0c6d59fc743661a18801025fbdc09659d31e3d219755666f6b025af20a991dff28e28e6f9a9ac73536f32135182beaeb9ea189f719abd26d9004fa22a91e11554ff292c3a6c54f13e6746231a0b7345dc803b0d7d908584fde3082be9d706f81adb1ac6e1c5553f6fef5f9d6566cccd233fae167bb28a33b3feaba8533def42e068946757b0ef615f33e28c573eaaae63b1f0b0a135156c6d9dcc1aa2e067b96fdff13ed657984fd01e9a588fc6309faa5af71a8f3758fd723987135b18a639525c2e1afc3e5f4cd926fa1ee3e9345afe9390749c4a6b0dc7d960408c921b0e7f87eef686a8bdfa55890cc233ec72f0ff1ac830cc7b4697300a7e9bdc377ceb73b9a15294137002ffe5020dcd793f6e41d0ee89298d14cac536fc892ee55fcad32298a8dc1d4ce05e15333b9bde92013922f4eb8c19020647a39f677ab3a2dad6f18bd17e83751b312941c83320ab62ad2798f94a99961f1d8e150bc30fe72adfa0269ee3f55079afa28e146ef18df2c00dd8c0fe43738c45d9957dd775cfc463edbba81ca37879bfe43952d06b9b1895957e3eb9c41c4e5eeff230e152a55bf192f5d0ac4566e43fb44496f7473ccf07c0901f3d2c511a8b68eb010964476917904cb8906a874bbfa674e6c725165841b8d5a343a967662fd474266622847be1ebde3f04ac1b7c8a39aaa695bc7c78239257b9b0d028e79a15ee7c34d766cb4341ed7a47f8d3a17f0c4b84eeba50232fe11f4eec16e2cf7475984595d048febb2efda3aff47d751c395196e73acd2cc24b117c24db22d3c87f2a0764ca10f3f95e5d8fdbc1d4817101c178cf1c31c32841324ffd569aa1c5d0a57e556cd580bb861b55772c9895d890fb3121c119e4f44218fa5f7f66bae6123a59d65e9b199c7b058ee4d5fc86282f3713976fffd1a0263449fe2f2a9436b2767c9ee81df2f1d3b1bd73296d4370a79288a18b9eade905882f26ba31ee8bfda5999467aaf1409cc9ac4e611572a6b9775345853293b89987f769e126caec985ed8fb18601ed082e7173c7779488d32f331473e4661a51e517b1e6d3a88ab8704b268d85b908ae62ec79130c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5d414f355f7ea11773dfef523910b3419d13a96da8c0c8837156f5350846c8c8feb6be507d1d703d3c12aa91c8438866cee8765288c6160f0066767186b6eba5b3ba97d47d68db732cd069d82ebd55976f4fdf6e18ea5bb7267694907d817a2407ecb64de765604ae0bf01fecb843b9e5fafde994037a4e9c5686c9bc69709cb60a5d0373403bc48a07cd54afaf0c85406ac74f8fb646eec18cbd1a87cc41b591a65839c838b45ec763fdec80dc222b109b100ee78dd9e8f822e1b9f5266f698e7d73764b64834e649345f9843921684977406840f40af9a426b20d15718d3aca18fe232910e92add5514800699a9547ba3f84591fd47c03107e403fa173aa38a38ac63a0df5fee9819fad288f8797b6abd4e0de6e18f3b2258820e71c26a0ed0664e30d674f02f07823fb7c7e97a9695e12915d0cb5e607845b18b76b847fab78656bddcad1b5a87eead687dd85e2a01e202fcffeb3709235acfb455fa9279c97ad8f7be1466f8d135b289629f47e519dafd85a7994af407a5acd048e9974f84c9e6186667ed392744e19e63b5bacc0af61d4bc98d710cc259cb7507c87d2585903b5235aa5b6c59d2043493d308e1cf1a1f75c4d091e9eb3ea03b59cc94d87b5a14f924881f2de12cb5b508a66bffb1cf91d4b159f55504720ba46eb51853d1364bf3cf011ffb00ecdcbdeccb14ec97580f45fffb6189d2761f42ca64fa1d21a7a4a9a119f053abed50182b373e0e3ba129cdab4b1eb32bdea79139d1d3d3182b2c6adb74bc20fe20b1042570d1baec96626db75f8be34de8299916791873fab1d3dd5e9b074d5deb034781f454488c4b368f751fb488dab9f989195bb6c7c79409c7a43629fced53e4df5da0b99e044881fa673d3a6a3162b46fddeab266a6288df0b52b2547a44e79f782b434acc353874fc0bdc4c687138bf4adc32608b8a344313622c504364fd0694b31efbda71d39b25f0f0baa562f72e4c3b697e36e07cd725cae867fc5c760fa5904c33d75afb1a0b9484c1124d4d412406fc2688bd2c3150eefc98946b54be27791274e6d3043f95cc0ae6344492b6a46e67f7c4c976aff950761bf1948caae1f1d683fa727ce238e2af2dd8202b8f3af47dfdd6f85fe1f055049067a323a17de143f002f08f9a63b5a8bcd091e181fd4a2e4dcb15c0667d7ca801df3c3b209d228887dfcfc66622967f72e0e04b6b5af656e40f04cc4779a9ffcda11a00a564caab561fe2e7e49a33927ecc4e9abb0b5477969b010074160e44de94919bf88fc96af807369c5b9b060c031f7e454972347e8039b14ee5b773098f04749ccbffdcdcfbd6e19ea96567f4b3e667fae94de53eaf588dcb4cbe79052ed3b4589c47e0a31e5eb564558efab70aebabc01e1fecba53b503bde55dfc1af56dc0f2e61eb6c6bc8de91a378a04855f8d43284627dadf0aff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h317bb05ecf330ba7e807f637b6d3c8d2bf349622dc66fcf75fdd139d55dd1b209825016eebdac5c8b1e1a11199d5b40282efc9ca729eca27f9f319637b6f98e813ebc76bb0d81827a9d90d0b9f9c7356165ea02e86536f86d5ab283fd11543412db57f470950a160e0d46ed213065e6ccec0af68c60752e75ec5a1f63c907abc2a593d4ad28c4e419523ba15f1389c5ca31fcceb149f481ec7a8c5af9a8c8b438116b20a9e553f5971740c7fb3008c0e81446458af7a1c1a64f227045761136aa32aafd76f2cce94488516cfa3212e263d1dc02dfbf2fb9a30da1f16344d3d5933231f9badd5ebf302ff4069c0888e9bf54dd0ef1379cf6d145ab1e3e240f9fc00f7971c29c2f1482596ad3f0290c6a7047f140836c5d98bcf0263952464875e72c305d2791fca9a0b3f6088ceb6be0157c0ee845a7a8e4ea139153f56c309267bf4b31f1b34149f85cf8dc7f6a10e01850b17af231b2ced77d585b134a63342f8b1728cb8f8feb64421ba6fe041387b82dfccc87b343108dd1ff63434c3d9cfe54e5dfcf0d1a15606d0bceceb012840027a4c9772bf43bc34b20340d73325ff3ea08ff1abf847e8f8b50f6d6e5b3b58ef6fecdad5c20beb5417f364c5a463c080a677ba887764b016bd31602c10f29cfa1b1c84465d24fc71d2937b328b49c1cc080425ca5eacf58653a27ad45727dddfd7ef889a7995742b52ccfbc0a808860fd55910c545bf15e7564e4f93f44d6cb46e09cb2aea4fb98d15481955608fb0cef368007298f8db0502fff7dad6541e1e52f2c317f2af6e4c6813b435900261faa7fc4f262af6f7cc709230b03f383ee2246bfcca00bffd3a376f16124cf5999efd2aae85c64dba4136b3ef237baca16cd6c98ab5415b6014d759dd112338ae86184d20e07fdd635f72d64b00bec96a23b37c0d57b3228a7bbf3ee3e4096f757b08948a393f03e4c6efe5ad7018f68bdc147ed0c3c605e7385fb9135f07b22f7ae40c9a7ad4a0cfb3d02268979362905031ea0c2e173f4488021f9d26e5485724152f89a5701c1105ae5cb85ddbbcbaffa9a36d761ffc7391809c3ed1425d72e4ccd23a2a2fc1561dc252cf49b9b9e63254de537351cde8cc0d91415e69d82d4e2870cd0910d0546d222c8dc654482e232dcffa3319b6fb338b5927b20799917bb70685f23c1d0bf33ecfff9baf931f19464192ff91b146f145caff66e569e1f0651d3e31421e5799323153a22be8ea57e3faa086321c943c4a1ceaec6201a047591130958c4feb0a306066b5e5cb7e11005c6ec37890a3ebeaa2aa5876ca016cce40691bf137504bde1e5cb0f22f21dc5b67b54bee22e530fad6caaaa34153de9a77e2a28e2eccd786742869b7ef444d0ab3e796d3e8b762d2e75fb8d9cbca0f52a2969673d70a9ad20c5c61abced615d901108bd3c4c364d1b068027aa2a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7a19d5a3a130ce2224efeec54bf5b08c7119896f0c9ab453e30459ef7d2027841e3a819eb60c791f7e5752681b302d54bbb8e6acd931152e4dfcfeaefe74e14ab5c7605b1978e30acf5b688651f16fea4969df091bfc85ce56c4be58b4becb4d972dc319fdd289e79d29593052bdcf3123d5888eba68f8c1eea0239aa9ea5b134dc3a83e180335ad1611f835c6c8c4fb22ec2e344ddc57e5861e95cdf62802f86caaaa10b661f3d493d1e0fe15a3489271455db1decfb591506ac4e5bc45308b80cbacefd57e6df5295af16c49f35c15111c446fdf97e72cc3d851fc102161b2fd72820a27c58fe1f5671413407e5eeb2eb6336a0e0217c9bdc174d598f4ababc335bd03b73f53926db72d98c9d092015c0416e9b51d7bcaf101a23abb5ce088255c75f71c1ec0536bd48060b546b3b0c1de59d2ed4fed000302a7cf82ec0a1bb522eeb1798ddf7b1f444a338e75b6e666e38b3bb2678baaae0b05376b25e7072e8de3dc3d5c2744be421ae14f2074d2e9833ff8dadf51a8238fb34795b6ccbd03c1d4c5c91e3d1f0224d57f831e4c10a7cd82880f77faa75e8f3319861b9b8e93b49e59a919620037c277a668339da87ff6eb1ec80e8b2d2b037e169aa6e50d4d12cc14800671abf159414d2bac9d6cd435c48175e53ebe1536ce0164c2a571d4efa110e4d12cc8b62d00c262502b3c46debc80cf6ddb720dd608ca428d23aeef3fc86b818728a4072561aa9e4d97e5972720c99c8a6a761996c5c83a109fc535969271a81badf0c0364d499952e1632278fe99ce63edf6d98028732f0be33fbd7c2a0dc352a20094097b4bd6a8800b83213970b99e08598ec0339f994c39492a7b5acacb148a74b7b8091978c39f98b537976a9f1e16e63a871dfeb4c28695d3cb42e920643ec9d1d29dea0902b2f61e956fb3e90185feea91058c693168df634c01dc1369eb13f6b7d7fced06d4db8929faec7e857a833d654d58aaea75ebeebeba43ef7f21667f58fa3d8a3af346d37b9dc8987714d70a1bb396f21c039a4ef9bf802e212d0c79c2dc875056cde90b6d57f889eff67f6a23d7f9ac8525edc47c1e1ad61b71850910a7a976a5bbd9681565170f293dd08896fe9060e95815f331ce73c024a5a6cdb9e46cd287d159fcc55da16575e1e4816b6431514f3cc7ecb0a5d50f5f88403ce0223f58a8d6ab7e5c48dfd88eac89f2151b0b4753b86274ec4d810b113e960ebe5dcc4e9578531914b70175d154a7b149f790a04aac57a38ac59fa4cddec912921e961a69f56f927221644acc64035182c68ef04edcc2bfe162f003652d3c41f9f0a109d5e339ded293ca8ff6dd83779887db076e72825639319404c5faab13c5d954530eceba3dfc075129aac457acea538da1f54701af8b5c056a8179cd4c8dd3c2ec7a39d90d71ebbe5ef12a16a62d2b646c3d780;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h76afb3cc89a5538f71d5b1f34a9b5a2c482b10f76d6facdaa61946c4977c87c145bb0b0c8fc99be6a006d2e5e1106c9d0e9acb6285b1ce7f24e5a622dbaf1e3e84bce0757af24133cf3312802255b9c5c0c9bdbd1bdc8e154c174ea96ae847e428c161dde3e142b78090b0af47f24c257f8e4cbce6dd968ee690124e9e644280f9330e513d0582089800a63ce51f65adecad6c2e3a6391437af08bff5a850a7daef28fc46864db6d50f6c502a40e5970e89105f29017a066cc8104f6b822b0ac4c955a4712f422a1dc3d50568d65944b25fcc260b842e16804ad5c3d8fc518cd24950aa20ca2704c5324d3dd3f0b1da2ef1d2d3af465c0cbbcaef063cc31b11e96bae3f1967f348c5401be6765139ae771238ed901c1c14df7bf4fea2908cd54e1f42d85ff537be017394cb4475129ce81648e9ebbf91b0d32793e555348a5fb94705fbf0fe5c72ff285b3dd9ae6949fdf4dd9010a9d2e96379668ab56d2db3ddaf7aa065e7e4abe817bdd61c36a00ff0c8871ac5af6ed36ea6862ae4cc24ee842ae69d4ca305136fa75e4c9f0ae6a110b30c5bef9b1140a8a541319e72b7df5460c0f62b7627031ff53e36faa57b4543b4821b65f599d5d3db8362e220049dd29eb60f88c438987cff8686c054c3742266651651e180d0e7046b96f78b2182907c391dbfd2391d6ca20fcac7f36789dd16d239684aa48da29dbb8773f43a2b1ec8372c82084c5802670bdb1c178247e10c1c64817131446f66a7a403ba20d49b79a2883b1ef751cafc9f22c9fd6bef6edcac60f9dbf15203cc1fe24663c1e24f7758e52fc071370de55bae1a2f2ce57a44ca3a7750f9672032dc35bc9425d755b2c3461c942f0544954877a80d8991ef1096bc3fd3af661b6a6812e2b87a296dd342cfaefbc56e19e56b58a738b73eea2672c6241d1072834a09e2754738f7b533fb8ce1d62aca2b3655453cb7dd1bbe31293b034e276642c5310bbea9ad6d498a11ce929b045054021c7700662687e6af5d15156b8edae708137cbd8490110024569c8ae4dfd558639e407d0add1c9d745f14a11c27ee5ce51452d6040cbd359b71ab0939c4d0e09165fd81154bc772416d170b5f7c07236989e88b140ed122608115b234fb850ace00e6b77192678bc045f01090d46756279496b7c2a64f498c3fef9224138951d0037a22d09b491456a159bd176de30f0c0c85ead5dafb77676eef9d28c76e8d1250d387c4861f8b201f86628da81f4b4868e7bfda98cfc1c4e39f70f56d093230399c9a4f3d85fe9b6ac9ec6d8b81d2ddc2e4ffe72ab52fdff3839afea0a39fa0d918809de7e09f76417cf5868a8d7bfa896763f855badffd1239282a4034adc119740c2a3c7f4cfe8ab5c717f9cf51408c2a54d9e78ab5dc3399b4f70be2a5fd49b9e8487402c55ef35e2b2aff7e46162622f4e98513e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8beb40fd9b9566dd4dbf4fc1b44d5a10987821be8be1febf6a7c922016a6f1d349676fde9800eb1c725f592c5e6c04b2debe7bda2992d91ebdc5bd0828a63363cb0d3178f13c41f922a265cf571fe3fe35844ea4fe54daddb8dfa87e711f225b6eff6b095026b9584eda1a2dbfbdcc722337edf51374942f867fa99bdc3a57c60de7074383d69304004fe932223ae290be243e768c6146490250ec4929c61f36e170a795f74e8bed004b1f98457b6c6e2151d71ad1909e99558ebcd9cbe72ef033a2cbb305e4a534097607b4ab4f5083956f7ca7901406736c0b225de016636c6f1c1ef665eab314f2d4e5dae35a30a962cbf218c359910c13d274b3935b3056de63d005dc765aa8f1340b291a28cf0f3eaf9859ce85b34dc1704e3a1c579d3b26289ff6217983ba713e4c193b58cb41f8c4fa4c902ac919cf3cecb2ebefe1b520459849286e1c157de53102423c5df3b52d4b575b8c756bf074af3acb74d707004f3fdf89e4979fddd39388964ae8b52695074c802f262742cc9230f9747ea785acc64f6de29696c2ab53839d76cc4313a24515211ce9833ff160355e77c2061f07c5d93ab920dbf151358f38a242a093fb543fa5dfc3ba4c864d2d0707a5c2ba9106e57d4a127ff321d6fc235e8f3680b91d792970e10df24e644608b57498aedc7bdeef53a086ad93f9e605cecffa67eb582241eda779ade84ea7e10ce8c8dd8e90d08a19dc0b830013ff83f04531a4a32de52ebf270360c628f9c5e51ec559c20aa69f76eb310564add606626d3e2f96e4a2eb37b32d81c4f3c5752a16bec447d3cfec258e217422a43c054f7a3aa0c8ad467cfa6143f6104078ce3bd46f6dc5a3907f39bd1f6ed87ee44ab312bd29b43f68c90fe9fecde977fba8b8be50bd75dafea421b7dc472970bd9a9bcd424607229aa731448e6d3edd9605449c40527cd86acfeeb2dfbe720e98ca49f8fb71ae32c0fd2fd6efb14c5fd66e1a37d5a679c4f027a4a40851c7f261ca999e9ffa1c09a5aeee440e612d558ea84aa71fe7dec78c222dc79d1dce3df3374bacaa9fe78e6e15d61392abaf396072b40644a16c7031a8cb49bc05196ca3d8784d9d4c94466187cd344a592715e7340b4f28a12ca0c416210a2f2ecb88d7ce373c77ba0a059dced2c38f23dac8dbd7c8ff26553ac754e87f1ccf3a83391e20df2da31d852523122fe4e3b3e10b480665fc1984321a13e3ffeb932ad920a5684f1700a25c2b79ef78553ab3342fa98b0fcac111d0ccfc52b3d909ee3a8cdf2605ae031ad4df649d25fb40c1cd07f89596f24ee5e4793ef3c68b0620ad3866d0516cd7ae513cfe7000aeb00c75f0e17ef8a1042526616871c2e9a192ae120e6ef650fe79619aae742e0bd58bf40830394bb64e745d8b09f0f46d2d8ed435dca91167fa92f7de8161a35863327e41b9af9ccee5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8e0993a6fc0f7cc63f219e27e2e5add5b8698d7fe77f1f06afe98a9537ef48524815763fb56680362c29c5e9b553115029453083f46a24e3a209c78f896d580351849eaa1fdbbb6ea203591c576330b3c9dc1ab7569d40f4d8930763c7f762dd7969f52c3775be5dbef572329ac2dec418f2245b1381e92cbebbbd1720ad863e44d7363fa2d6343582fe22d378ae4d7eb5d4e9892305c4ad63919c4ec7edc502c14a3494e263f74db5ca15fe4c6eeb5cdbbaf2cdbd92e0e40f6f031057a17f8639aa5a886b1107f63f125666d47915ee6763cab25f8686e2ea09a57b08e3fef14937ee6d2ea9a2cf020e9be8f9dc25b3c3588a9a031684c3c1c4f1ffd6b2c4628aca60bca477b634d4326c16067fe774c0e32d7087fd447bf4aac7da34b24223ad7258a76fa763abeea8a7408681b19a6763314ac6eac8565bcd53e9c2f13c289383af10b41817d346eaf809bb2cd10cf8256701bb3c44e98e9ca1344c3a91b97a518a10177b7626599c06ad919f1d6bf4578c3bd6e8f63e14be7c983c8e7923ab01fd5f69412a85af976f2b212b82ad76b507e3c864b951936ce41e78b3f2348c18361b09933278e0747d9238b922886823710cb2688dd6a4945579d9922601aeec7393e46f19b33d0ddf5f8fbde910ce148cf4d928da290e5529dfaa5fb7d02ef5bdcc2b4eb7f9f41a24fa921793311b703ee615956fa58c3f9c59441fcaee301ec1731d3aad9f3c2872812640f73789e0179000b5983e1484bc68f70bf13da74aa227cba8c4cbc86f33397e5f1c772bfaac03b03a77a8eb969654491a99229da1ed16fea596a4a3b385e765c634a78de2955e5391766b04f2335f88fc3da8d6237b34e06eb85bfd224cf8aca91deebe600abdbdc726f0c906d18033a5cc480fce65ae7a46e815f7305f056d50639b1aec025e8a6f6320dfd2ea84c1e7a57407432a583949cb4cac3e039e3414ffca239f37e5b8067c5bd3479e8a776ad25e4bbf22fdb380391c61f2f07d19c42ec0798b0b99398b5f67e4e0ccc7025434b193105e1dbb4cb5ef2ebc04cb3d7a6f8df5a3e29ccb204e45b3ebdc06dd7d783b46169a9927ffcda3eead33926abb11becfb9dc4f2cac557d76f1c3ec8aafe9cfb37cd8ddfed6ce60bb303e25c5c2084a1267b71f1cd24bd538d6c5d132a9307bbe645fb7ba7add87636ec514ce9a999ac90afc2190a1456c2ead59a3e6647f9eb1d3dbfcd6861907c72ed557352f3da77169792df3175c7faa315f92532defc841e83b3c5b777e2e2e5f023f1559203b0a6d34a4ecb4aeec8bdee58f782c9476ebbcaf2ac56784fb95106d7c31219b77896720e9e0e2617543f784f1575302564b39e8fe367e150e69ae1933f677525027796f11708669b5b537ee78cb74c62c573d00e569434eb9c947487935bf391d3087cd3c280494b7f8af143ec91220c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1779c2bd689800285bb4f254aadca6a19c8fe8690272b13d3db876403e7f122c6ba5fcc73139ee9be396e3a8d96c653fdf4f54608a6d9b67de0a468b6767c50e2aa6410f935c2ac0486d09d0ad8ca7317a0f0a0b98285685f0be8bda7df632d21277cc361583dbe03ff65d7a2f44c1bd68941656338c1eb86c4461afdb2f736d74283015550284f6f943e5cf9399c6d075d32e8fdcc6b64b53af606c21b86ff26c4402c5287475e7eac0abd2c28aed6b4991384160cad10ac8dec9fdde8f25b0598c12285938446c94ed5a444fe021f3d79cfeca2cb9403cd1af53efc23dab0b62a0764fe4c9b66a14f1d8daa0a0bede96726bfe398a04bc13462be6397cd803d4eaaa8463aee6754307f6d49442464bbcd670665a25c031aa38d414f025a0cdd80a7414a85cf0bb87b31740b10c7577509963af6f6b99bdeb3437da8a25aeb002879ef9f14ed5a639841d76046aa4acc5857edf95cbe3401879873f73f2ce3bdb5bbe681d2921904c8d00fa3e541b5dc728eb1e3d6646655027ad7a11adeb0db8bf23e8963b8a33489f8a4c3a9c06ae81297dd2ec91573d14a081192425f0eab307581fb7454233e4c45a2aec2cbaa87a143e60f05454016deda78b8d4f61f11aea34328db784181dc77fb11d41fc7b7ec1e7f8230470d7ee9cc92be60f72d38024fe87a7861ea170e37b0a2d5bd931f00f96c612560eba9c534c2abdbe19c6371ce918911c2a5ebf089318447d8607658622456e4de599293e9f7a3976c1baba0980ab3c68279a6a21a88264b4a3a74765d444c2e813ab9a0bb5f562abc81c26838c30b2518978e2a2b5d85a9474e5792718cc60d9638eb27e166d402d59719bafe30d7b837bb51ef076cc0d790e2b948c9b25328c9660d2ae469728d58b321763161b0c4b092ac61bc5651a51e79b9f0f899dbfa58ddb5893f9d7c7af8000edb448c67e247e215e91f549056571e39c5677a51687568289fa0fa27e0c107707f39094768137e01999cbc62072de712c3b87fa8578f3f94217f5600b6abecb5cb105d69956a1673429cdac151bc36f7ca11ac705e96c53792a5f8476bcc6e77f8dd7a5c2ce79ac514aba78aa14dc7cb62ad4d13c6eced304bb3f464c7358efc4c889239cbee1e4caa63a1b23f6c5c03ec37ef93e92b27042a2bb92b7f76bf0b58a55e0686077416cade700c590344a7e49b34a771afc566fdcc8b1f3de414c6a4604973ef8a8700ba2f9caec8305dadb99968ef677c7005019db49523dc91f5f9d7b82e412926dd339b819120527c463dff9b66b50d9e5328624d7a82e5fded84aaae03f00b8175974e085e6ac0b24d2a9ef55e8f1576b00024310d100cedae0f39d488f7f35d26d3613764daf16854e0aaf7278bb6d60bc87bc6a498f2da40c6ad283bae02fa2f20e820a189371d9e758cf32ceac4ebb70cd38fd863ba7c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8aad2ae4bd33eb2316b8aa850920c44eba0df4d3cd5f98a7386d4df9d6160b5d11cc34241ae5885b83d78401e6b046148f68a6f65b29025df4dc488a849fb5fe92cb1d56ed280b031d8fa5e7ac35e516c44b68de2ad276fd850316f742a0d85e47765343805c93bcb2edd6297830280e490f26834daf7d49cafad27aacb6f5342018826f11b01533a9aad1cb34defdc1d1c74690b3342ec19291cfc08c8ec196ec396b0a695724eed4df87512f6e8b7a3e6c5a6b3950cd2b1e5f45020d2e370421d54d4c0725ad5b94bf5660d76e0e5400299e87136e45b75843435956848c4cbfdcd4c9775201b7879c8b87be97751a203f03b951a5a8f836d5abd0ed1ac7da0d56af000e45042cfca9a0ab79b896c2f9c2384d1077332cc7b4e826a1cb001cde8737866bc8689f57e85a320378ef0c3da9f95a991e68e6a4329b05cec5a90b9b8b9129d2140553fb6eaa1c8d9a25c4f7ebb2d8a8cd85fab2d8fc258d9def872ea11de6d45116051cc7707f715112b643073ab62917d13cdf4033d259d1c6e2c0be021560eede52ad0475df6c1d5f46946625a54fa4e8044569288b323fdf0e2b22a7e5597b1288d94c6a7b41635885d20a055f881dc525e7eb77a0470fc1bde36d7838381d5499207c51fbdcb7d5e933cfde4441a5890bf8abee4cf653f2b0b2ee6f6d0c3b11b39064fe533a384ff798b2d651c52643329618ff80d9202ae5275be7d6d6b9f90404d2e975613efcbfc22028a372eb1c28f6edc2fbdc716ec130e9dab8aecbb15481a1ec045fa051260205f7248efcce18609e411aa0ac05782dbd8731f9b34ce2a087156c1d647165533f8811ce39077e214b5c0f31c9361d1ba7dcfbb18e8862b9184f90c62bfa22d6400fa56b2831762ffb01083c74fd0816a397635cbc9a88304be4984912446facf39e5fe3bf5d25a23a68c66211eaeba31f7e64d1f3fa002d4f76ca64b5eaf94361407000c1d7bb853ba1ba64fa44fe919ce520f4e2e928fe11484867156778b545c650ba9f6677947a8749ef84c7811a5bb4b7cc64d783a5bd52a0c3854bbde9a9acf52bb0159cd1a43b684b77e1c409cda4de690d37bc19aaccd260f757b4958723d29f28341ebbc05b7befbfa30b5089ff53011ff768a7d33275fc61dde8fb27302f2d1db2b09fedbd7863da35cceb9aa2042f8a3e0b0acff2b4d1ba88018fbb15659e022c210020bf2f5632160c522e310a65eaf874f75e8a72609d3a225ac17d940eb9a83ec605075e0e06d7f48c60c55801d71dc4e3f47d54d9a1e1f191c3aceca709e167a26cc31cd1339a4984a1ab2ec86314b29fb269f8ee4a2ae8349d3728974fe865815672582283dfd2a6ee11b0d5fe19447b73c71413dacd8243f48b9c4b30a87af2fdcbc6bb3538eb1175e271f3dcea2de6021b2a5421e538323f6a184b72b00190e882f4df6c364a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he9c950ea6102e0231c2b30b3f6421d3a572ce798a8ef3cd5150d94be53d3caecf5cede297d16be6cb7b7f7a07d9e3cf8e6039a9fe3de2b1df9498fea0f111ca8e5dd94206f4206de13b37fdda0599c05bf71b870d02168647e20cc82ce9e2669694ba3ff45287348f79223325c36c5e5e3407ca338551b2500d757e22f7b0b8741ad4d5a1ef18587e9cb15b87742fc358908c02648d12cee339f79f52b200b742a42e378e176ccf073c991d83fbec0578587a14669093827626a4f8094e344cbcad6cf0161ab93a89f410a778c881326a50cb9c5f86b47ae930d8b10b435174d1d60692269d63e3c56f4c8409ed1c3e0888e27097499f7277114d1ccb813a5771e9cf7fe95ac82c1d71d140a81d1531244f19e86aad9251e0693ce9f8e43cf6b74c6ba79c4b7ebc19810c3377c5fed72e5803a80ed5034192916285b0a77a7fb3d540662b52defa12d1f53f12771a96618f08ba1c7a4c22481fad88d6fec8295a8333621c42a3f044e1b79707f05d620bff69b26aaec5c42d4af54269f2e9fd213b7ac12d7cd22b03fe6895bed7721c59bb7f770c3a0eded050a0f94e54024084874cec2395662bc2a110ee1fffa5e57161615385ff04a1734e470d2ad19007ed583b96b0dd664c7ac13cd71c3595654204ded18e7e869395486869d42a4c837bb5d118373ab72b72f13be7115e8a7ad5d0d7669b48160866bd57b383fb36903a3849b3ac5bcf24a4ea06989134d0f5a95c4ed8a5dcb3501a566e31a96489b9c37e66f04720def836bdbaa5760b033a8168f827ed81c7693402c6ed6d5c618cc1948b8c83bf5371994829f82aa487ded6ea3e9bb111be28ed3376bdc1fb96acc2bd034db581817802887a632954953e47f46a4882ffba0491022e09d9de422b434c2a288321f5e2dbb1b3e27d208af6ed6692e64cb869b86fbc0a4996ad7cd32ce102ae6c88917649d2f60ac6054c2b4e93e6c8d5ba106c3f2674a1f103fd29ba35dfd0bf2a8c4fffb674e53abfaadeafb6ab89e01cd3f51bd73de0e9b880877b27e34166fea113116d1eb935525050b6590820ff4646434ee531924940e474a8bc8d7e37d581c69451c5b50c61a5f6f620f43773df5ebbee52a09e697b96d46435d6a332dfa437ddf92167a6a73404f1fc22d149f57833741e8e7dfca0ed385bff3f583a5c64a0dbde907d5815062247e1050cbf498d53d7b5b4f0e2b042ced7317f873c4366ec57fedf5cccd9f2511b360ffcaecbd02caaab57cee7abff23ad0e41051937f3febd7c88698e1a961f230246ab5ae2b7d9b2ce2586198a785a3922497cf2cd169fea888ba5e521678a7551486a6d67cdd1801467c0857bb67defe62964c0d1e3ba8e3e6ecbb98356aab3744ee1d4e0f4fc881b4704a5383faa5813151bafb89b6f576897e46aa8ec1bdc81971bafcd17a1fd05bfe7ab1cd0684;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h57c865663e917eb08f509eb15a88d89db4544920951ad51f5146e9f96fe8cc694697fa8f65786a928f7d29df786d250564dddf40938a5b9eefef0b28017a4fdcadd467103e415017e2142e128ae46df0b0e2fc46e74443e22f95d6fa0ee115e7e5394b786fa5739c6e347912730cf1d1651e72774790e30e18929b9faee19652a41c82692962e38c7ef8d3327e2e43a9beb93be258bcd5512631b5e1d461ad4c38894f81779ccb88bbb4da5b084729b239e938457a9240fd0eb9bae21b581f7f37f22e3fc98b8cf3f2043c0e1eb4023224423d9a5eac03cb91221e732a4778de525cb3838ba42a6fa9b41e57b0de286e08c8d2f5c8defe8107a3a6c81f6a9aef0c417a49f517e4c61504785066b4af7102f0e8752d2ab4be96c7580b4903cd8f99cb00c7cb413273d90d770842953f84f30dc5e95dcd5d97f51829157df00b3668c8951dfdb107f7902edf19bfdb97b0a38c0e867b9519f4262b83ae21b731e25b5852b73879ff775192b9d270f8387a107fa180fe98367061a67e611d8fce43666c142da71c33b95b19a5d14fb84901dde5fab0675355f75c3e79b9db97c4b1dd9eaf68c71f40a03f2614a588ed6e7809fabe20391c77bb746b466e10f1fec8739b7af5328ec36d46b5fcd14928ee80ab1be9efbae8a43fe649ee084abf908d3d9348cff8c3d4d7a322dcc27a4545dac627f937fbe0b617b9cee795662a1b07897aa70a7726acfb0c450bb435fb109f6cb02e88ac9165df0c8c34878e00f3ee8af169e4b595d43a973ffd96305533c6db59003ce701f353b3db555f6f1bf1f7fdae19812fced23e0363fd5a59aeb86de45dcdb1945a5e6e52f742d7897d2f8c27d00d9740704abe4f01f58cade70d4f420d03a558d515b22b1ce192068aef83044d887b6b9364e9242498bc02a429dfe74b5f299d7cf2e91b8739dc3db887f98acb866b6dd4359e74f4ea04cbdd17ade5b48fac98e9e5b58adf4d92aa22ac083c9620eeceb57efa6be5f89dc55e39952f66fdd79260983ffcdcec6ce29f54aea21336c62d312c08b71678dca9258b60365a5d990260b20b84ff315be90dd040c11f9071c4dd937d5f4eae0adc586e72c6b78ac88c2af64eb9c3aa8e33a7795cc2268952559febf0b0c21be429976dad454d0826da6567c634f069ffccff604ca577bd753545b075b19ec11fcfbae983c60c992d2904d0bed811bab70f50dfc573978c30c2707c3349ce1f02d12581fecb1c5551ebb741af5d5e8a58953fabf910f7e380c22b2470f07be8bda77e6b6d903eb2ff0fb7286cec9554c602d4cb946120b4258e191722e37b0aa0dd6217ae8a867ecd3250433d10f3246971ab439d83749db6f6d2bd892c79f2f2dd9a487f36997385bd307a7e88e85822fdef3dcb84a0c78d86d5695f4a92eb2fa049d6656b184ad7fb7f9fe6f593412b7b11c77a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc1f3224657a430f88b011f6caae660ac8e6d8cda7444813f1442c0930408cf5aa79723c4ac37c19887610f62d9789200b863fa99f8938e2a269dd91ecb6dd137006aab416eb0e8715d74803d99dd608aebee9d44b360a424aec0c940dfbaeb444c438e24b28af43d5d4544dbc4b3a5a873db30b78c43b6a37270eef929505a7a314160f1329323623568de30a536b5569ca328c25722f62b5ec2fcb0f21f2543c667a7d21b2b3daa1c0385fbe8b1a8eee81f0529390053b43562c44bc694190557a444c3fae9df977d342036c1378ed26be7b2a22ecafe30c4a1a2e50174c29331d5918e2022ec8fa862c25a0718cb9988fb625230a1820a2ae53abe0964d695d848b924f8cfc1922fb7671518cb46b1445c5e9cb8c9934ae92ccd4a8a314de1d82f0f488f47ec1a2ed10bd75cd282dfc8964ef255a68dda709b8ff62d5433ec4c84e2847fedf37fe8c2c86e7c97d71811ec1bd63e443dcdb9d50a40efa912883e3849b23a92a167d22cae68fbd7d0c53dc5f5c9524054d704dcee9d1b993d6705fa57496438f4634c46038b2aa6a29110c6fdf99e765ec34c0fafad7dcee5a22bcde15cf83d20918af1e131b0ca86de43c5a7c14c39d68dc60b77b73c98970a37e8ec6676ccc9254b04d0f66cafdd05da4570ba827f087e59a6e787a81b784daec684b66c6de9aa7ca7e279b019a6db0ec073d18c97f0b526268619311309093e6510aca802f9c92c887c44d886809a38d1b82920a121cabcacec178b46383a415f22f1771c12b166f88a2fa96c5ffd36f7b59c9e6b6dd63f4be3173d376148d77eebce9e67ee7a48575aa437793363e91b2907eb2485344edcbd569448c83862f3a9d720dcc357ac924e522602828e151dd700e714c25b66a82af4db36f1ea48902fe0960e23100bb8f8949b6ab2a909128235acc9a12d602593a74f99e831e8f97c27f9c4992b07f0da9b91cbb30aafd963367594bbf016bf8dda281dbaccf25a5ba6852723da5fef0807fa07333214d7fc60627d8d414fe6d8c55d3f57950678e8ebbb9265c9dc85c65d6d6524a19230d66fe9106c3fe0cfa376f0bc28cbe7d485be6fd05edbf201059102587a84763addb7a86d424aa25af1fb16d5490b9d618e277074474cfdd5186ba41e4638d73febce2013a906d6e8764cf65b02e65e38ba26cc1280d0cac3e4dab3a126c50d0f28b00e98b614023307621aef47049913e3d78bc37d76053cafc1d9b2b3b2e0c1a859bc5538c0e56d124e5c54302d1740432616f298ce12d0c0202dadb4f4296193ca53338884289a6d87f907d3f7ee77fb6907c9b147896a64dd3e88faf3c6fa4174f84690140767939c74c71d6459e5d737dad2eefebea7e6f3b5f6cda96cd8825c825b16d83de60fce70a05cbbfc974ab8fb787527f37e2f51016d5eb1b5c40b00442b3a001f59c49fea2dcee6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb2985f6f3f4979f2001c98f19ab75eaf0c66a4cf87a7675ab25da3830ba980310f9ecd09d86fa741f27aabff48f87afb0258e73731b6320b45b024333b81e797f8065ec8547758cec929bf0a8731b6950a46826b35ae6cdcc8bfd62612fcf7f9b0781e546b78386447d329648b2a73708948e2a67cdf590f24db0f20bf8d7faf641975a178041ef92126693fbf6d0441529c6f683870fdf452eda90408ddf1bf6ad4dfc1232dc109e98cb31c665ae9c1405c8ce60ca0b864aeea7fe889a7da31e489e9ab12a973aefaeba0a7ffe06e2fdfe96cb07224b520f5863fb49213316419cabe725cf64898fd1ba40f639159a26023a3f5a4c3890ae6d209e593b6108a3e9edb21e0155a7fdaf66b775bd5a763dd0e4884269240415ea1938986144098ccdee21323a394813b69be40291f65e95d730703d07654ef07dbb362a2acf9cbab921b8ec45d7bdc4fedbfe6c346fe0f642ddeb2158ae9b0d932249a7a79f5ca3b7c372d51cd4e6a946cb9f84cd180a6c5eb617e200bc7a0cfa9f0c6a852da1265c3eec7e819b611a4536da7ef9617928f4b324c08d56cdc11fa54a4e74e9eb7f56810fffdd5e522e90f060160422c709cf148537c4baa77e3c92c6ebeb9b2c0b840e0679c17722a9b1b6af3804e1e94851f0fd049f5d67a8d9039c2fb9449e381ab559ee7e208faa9b03f40d726aff6e52f1b34b925c71374865429e1ed0e7e378afbbbc0b12ea6c08bf0528b624932127c7a59fa72e9dd0d5469a7752d5913b47130f0ee6337de2755f586d16fe7d10155fc2c3e8b0b8300f55829c76f9e380ea71ed6b75573e7f4d904c621b7a6bf8c44cfda956762270f4becb3f649450d1eae3dfbaf95832aaa6a49ce9840bc20e6cc65675462d622e01f3817da24ec9052109c8861b44c98833ab2270f93a0f313a0c30b268292d3e077862734d2adfb4385ae194ae9bd0eaeadfa2bed27e4dbcf49b4e8c050a8e699cb344eb1eb611bb18b2e7fff17a68d8e8ba748b0410cb000f9c1ecb3578d53bb821dd7abdc5bb990f44302504c8bf5c0461cf5bbaab9d2b2df6df65fcf9d3f8f0ed419de8347c2163a29d8d9e0d92755d355da6ddbdd3178a9f3c284642366dd1a5e57a7903824a6c876d4cb58df59e7f5b714c97997e32d1eddc4a4e983eff70bcc4f07edde21b70ab972d27cce80f3296a6970b5c74de5336af836cee310aaf1b5ae62bfd9ca3641e7af40502be460a46eb36b86a5187a26dddffb8e93a6bc2b36ff5ac11ab8a0cb8a5e43e64f3246d701f4bce6fb9aeb2fafae2d955f31de06322491678715e1be780a3b6facef43104d78aab12fd91e4b644418030d9a07ce539b89ff9e2d49f1820bee80169d0c5fa1d540c999dc211cbc599c412fec7adac74013e343968a110a252c6cbbe9f2a12fea8c62fbe6f3942bfa9a0b291c5fba6d860625a140;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h88cc2ec6ed1a0765c1cc998bb1f40d3d9a87d41f4543a63d011de1138e3d233f2a24588b83f7e6a2472ba8834b13f17f17281f9a5f1876136f7a51dbd34628c26d901da6d23ebc0c54492e2de9d1bf2e3a34a3762daae1ba21fb2b228a63a5615ecb040c9dc798dfd5d04b4f0465271b3ed3dcc16f97d1169d4f07c9c21767bcc1b21cbc9281bb80ce7e020b9421fdbac7b402c8fb34140e9c057bf1feed8248ca7872082b9c2d12a00ef1b7313f925c39ec0694d915b009b17b9dd9790f5e3ad3eca1f4d320efbeaeab744a62dd16e25654f61539c149c225314dff1dd28cff3b5f03c14863eff57744a047c9a7f31d14c2d1422f819a96afcf05a10a5d434640e127443a85dc4156daa6dc11565d6cc39a08d0f40ae93d1da6dd4db376b9bc32e73aa9a016f0cc18b0db799624427645a009ec11d85990cf9ad5dadbe1204defb067454dab2b160611bcf5ac23390d652f50c90605eca9d3b8b5678ad0e40413bcca872680885940b9f545e493e5284879aeee2d8e3c42d756bb0c1f20aaf2661fd44c4accff5e13adb89435947a54b6a2502ad41a72e7971558b72d5d8b4efeee6c31ed687bca5c6e3f12be2be971cb469b4fbf61887fc209e3cea90d90fc827d8761b778c683489c5f4bc24fc2ba2dad0b84e51c9559a8725ca89eb400b48dc8b4fc302ce40911afcf348ebd31773ed7cccac48936eeb63c0199da8cb251ba54c92d7794c9f0aebd8f5b36c90735726930e57974dc5dfc1e57c8b1d3e216077c627381cbccc0a6d56253eeb571462043653067f7ecd4d903ba8b53e96eaded53772d24c2a6539cbf1f87bcc0bf0c311a424c84140f52348cf1992f2731f0134d19d1f5ca5f8eee08ea1accecf6fd1586249ea2ac2669621c7ddccf110b3674524b0c8675e4c10bff334755f7de83ef78e623590935085fe6d5f7d85565481b6e1fa751cc86b0cd28b22792b83e462297634386eb3768e6d2dbd1e595ee9d80e4db658ac72a2fbc31067f02e38b00efd63e92064b2c690a9f9212b246f4122f1ed9bcedf78d692b38e17220e365155e0e0021f92e36b53dc4394351eb76b0cb3f489e038cd192eb1228918f89fdc054d97db5c42f53c1a31d40fe20f91ec23ab5e82f648b606a01ff6b4a7e60a4ae13572da9f908bb4e7712fadd91db6a391a6f8a092db2ca7f124f7ac0673f9975b1f7f6312983000da532e2372634d2b5ff68a9a1caf77e173041279af31c88cec6ce3637129c75c25f60e2c96ef947f06e818749a99179b0f19f910e0c80add4260d6eb3a33c1168d705014f72a4a1dc8f3b0d31a7b3222fa55fa2322fb1d5de71720e3d7471e8f99a1c263682951aa4ef6225ec51e65b1b502e086874c8437173bbb7a51fce1a63be639d5181adb43449bf9a8c5374601c8f365a7a79e1e1b731ac9f5b99994de82b339c1d158d5964;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6900af21ee96b937180d2b75b28f101278ea4c92880ed4207e9cca2f11320401a020aa1fdce40bae9b828011ac8312da9981bb814c3e438f4ec28259f4bf9368b316c8b3a206d516740b96a52308e077ebcd649ab7a323bfc16adde577e4a5f1d0168a5896fb4862a5bbcd704074ff94f689aeb92dad194d5388ad3ae52c313eab68ee87d4bae6149b1edd6df098d5ea9810a0eea3ba4d5e8340ef30d86829020509c58dda437a9473441acea101df91c37acd26100eb460afbe4f4c68622b4a42c849df949c96902a49c4514ee4e7e387ac0616759bc243c0d77eae1025a201ecdebabf397e7008e12599ef4ca5b28fcf8a3abaa533eee573e0ff6dc23174b5d47bf7789c0f2b633ab00ed48abd3f00142ac0672fc94371c0a2de821bb9c49fd3b85d0c7894668b9895104f698d3727235f444efe7b61e06576d0a97a32a9c6e168e51281279806a101bdc3e767667c4b15a1c8fdc452cd034e7d491eae46b5c58c2254d7cb8421f4fac449245b052eebafa49fec31f3eb1bc082cf8bfa62a513f13fe6264990d34e0a4531ed919eabc6ca187466daf48a8fa872892bf4c9daec9633d2135dc5b9172aa3a247c8dc4d2793c0eb6f02305a7f61ce1a39d7b8c6a915fdcfce10bc1c6e1e37b5f1073d608121f61e8d48febfba7cc58c72be728bd2cfcd3298d2afffaf55117a9d48e641216b7599fd51ef8e3f904a74236bd915f1033ca91fa66cdf4e38f96caca41fc3ce391a566c78e4b592bc4cc3e91d73d4640ff2bd5a2e5a96862759a29bc2f339137771e898b68e2857c621450cf41053bae23579744b326d573464a23ccca1335efc07ab2d1a8a5d933f0f75112ffa1d2b1ac5b278604a9b42d215b4041f3a4e2bc9b37d994846b06ad77477353bbb2063104136481873e6f15880dc8005c88270f507ada746c4e751cf13a4542d7d671e0efd9eeefea85a1103b4f8ec8da5d797f7da596ab0772aa1aeea49db79a59e201e95b6f41e3366dde742db23323572f59337e687eef5cffb72ea11e9a34b23081b8f5fcd149318675c0b8e44f9294b2dc568ae4b0ec051853a838cb4a1b3c3491b881d762f8e92d17443568c6cfcb219254b18dcca4a75d22d8b3cfc97719b2081d55db26f56ba29e3110379caff5a64dec00bb45ddaed5e60e1fd6b2b2885f00a678dde68e4c7d0e35afab50007a0380769f582f18530f6a59868c11a61fa67beb6fa657542860820a3af9c098f8e58de69498f813c60b844e03a9b3c609c9bdc93e55da6048a09145c146266e2a2f2ab069e2b5b227655ec87b5f9e6b9766bcc462f551b119a9b85bf1b615e1c8656703f51405314608b363170217234757d0edfac6937e381073133f414f4c6e48bc819a7bc860f36022ef7e2fbbdfa85c97706399d654e656618df3857031fd415989854b2a037077beba9a557358946;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf7357027734b94659f053915bc6d7a03c910ffc2d01d0bf4ffdbf73353d328fa0ab6ce0ab0e1b8dbf2e9ed9f74236be6444c6c20bf299203f6915072abb31ccb811fd480bd42f72af70a70f77b9705a1d35e41ce7d0e9db90da5a776676bcc82345cb0bb1026fc7ad3665885fd3280a5fcd951a6188c88c56682caae73a634e96535885b4b504972e766147d6e7d44da95498e9e4b075592d3f6d753155ba989d0751f738d00ae3e317440cb3459ae77954b1938b56cacd53309fdbec9e0abdbc58798ee2796aa0d217ff4733c0ba90820106b5980c629308fb1d7a482f8d6c7fda1c70eda163c61d742d148633b23671e9ae22e5dcd4a7d5f77a7bfc11ff27bddbe2e272c94b1739deb73c531c4aa171479cd7250df8d1884559e8663220f452b76c428f1b499f8159193a6ce9b87902bf9064bc44c44817d1fb6de7a2c394bd262a2a14a67e883e9834cdadcb35a8c563c46bdd9e6aea0ee30f8faa360d01a17f57a04981b6cd946959a29bb45b80e01e3b3e4b258a305abf8a4e826b0f69c478f8ea0f623e8fd0b557d73500f6f16685a5c676ee99556df8f2e615b786162cbde62d65a965cd808c549411a4ba3ffd40c47e72e36faf6ee2c5bc4b9ba89497ed679c52285804a761ad6cba73518ebb32343c7780baae3d714891d738cf11f585ae1e9ef464d6f5d10ad977cbcef8e8cf1f327b88fb0638efa47e3c1ff330670839d3ebaa6fd6d1bfd9e8ac1f648933096680824fef8fa57c3dc3bc36f9f230bf7cd80ddcb94ad7844756104f51f508ea39c1d59a8545925f931b066578391217b42424da5e3a3788c93ea9aaff4d8f8bf039dfb6f11902ffb975556f8bfb9cdfac7cfc11e68f77db557b38e1908de71b6e6ec08b34ef6e655b9898ebee599758a1f81b46c0f5399fd2b1b8b310d521f4a2e85f0806a60f19b319053f6bea643e2af5f8a7464ec9ab1986c5e6d53ebeed825cfd22598540f375e53a00a046d3142717b3c719b3fba1d2f4aade61cbaa24bf6cb86b16994af5d50eb84c6b452f0665160053fe04d756687877d80a409b7b29b4e3921ef0196c5e8aa3635f3acd4579b2747a768a04f44dbbdcab386cc61762e5f8c6d876450ad5b461af00e91984d0b020a631fda4bfa710845239db8ab236204e9453155ea0f7ac45a04737ebe527ec76ed757975ee8195a1d51138994d7896724bc1e14465adc75581ecec183e2ced30aece3ca2ca50706023deb212261abbd0d4042e1799dd475a295ee1c5523f25f0586003a8ccdc2e6d4cdcffa4c6fdb2d65ef3fa935c841b3bef04bc6f2d4bdcc3ca465315741392ec4f01e61b0945644b889407a720219b9eedd5c75cadc297c19dee20d88f2e96176374e55d45cd6a4c0609513a112e032c41fc43c6def8397c797bce66bd4228e966622f70a250948b7c0f27c497c284562c99145;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfa865c927ca7b9633173d9a3c6a7582276a9954e0639c3dbb4e112f1bcdf05f69a39b00cd10960ee6ed630b4c24f4054df0a740fb8564d772bb2ca7d96541b438e00ab327d259c3d762d1870301d28e9619efb5bcbcc472e3017d863b2f6e866908e69d16220c201c7430786cffd89fcc2d4de35e8a94e986b4ef7df70dfa61498d6e089b37011e2e83eef928b32f7e54bd2a913b5fe3c336c90d670a8732f045fcd2cf1ea2847c179e9966e3eb649ff754fe09888dcbe46f1665b76d4e74b170b5d3ec1ae3c9bcb8c6d955315c0734aca3ccb1c3c1ab2d4e271943aa9923c98218a87f6987d171671006a8842c498f59054ca8201e52cbc85439f54c66af24920289852734dc985f3b94fd9b6e89f41067659ab9155ffe6d8c96e4557deb96653da992e7afc3a314bbc405d0780b337adabd750bb08a20660c320e1a9a6230f0fd2bb2247235f26fdd124d64017959adea1cae13df9fac90f7816a3e4587398f20a6b6a74cd3e69731b0948037b74496fd9328ae2dc0b869a2da5aeb5b7d286d38d5f9384744128b7809cf69ddf223b6305792d0b45e8e969e9cb8f81105069dafb75dcf60fa5be72b9ab526da45c42e46e0ffbedb9745d3e25d7bcc6c86b041112d1fd68363b8570ab31d943dcf8b9fe02a75b34a53d53eb6a98a8e39353e18a0d8a3c629378060f9c6f87c102068fdda152d2072757b510ce59c2e67aca33ce3fd7906e2f842121f1b89c814f2e704d0f4ff49b78c931be4e32a3caafe19c557c2c596f05022a91019d279d3242eb1ed6af434aea6ef231100851b16a002ad0a3d2244afe6d58ecd3da5888fce600b5e800eb2256326089cddb7c108c6738b6be408faaca13fbeac20559125b60c4d2aef9feed947b24d1d2fadba221899513ff4e95b43c63f72a6c6db506aee7b955e243d41550d4551e71f6c45608aa7b85b6d3c322d3d8bf3b948308b018f787dacc6a2ffce7cf1028be0e1eb59b5479c71d166c1057e2762e2e6b47ed2d6a090802978ebbd670fc3d695392d5e70297e5519a17f432c48ecd9d048a970ab1a7078790923be67185db024eb6cde31bb2b2c475a75821cdda2d24b2137c8acd270f031fe0c31bfeead1ce0888c91b4ce6911992225a37e511f7eeb0421c5644aef0073eb6e0575e39159d9da0a82f6453c28df67f4706cf34e397806e06bcc143563eda68fc32af2808fcb3cdb52836f80fb7fa33bde99dd7e6d3e1ef3a90ec3bea794f90e02dbb130a9f4dba27fbef20c9a8939aa5492f326fbf0cad21eebb7ce3674a3d7bc82417c6cfa249063e8097839ff654ca32dc56dd85cbe7f0b4689feb9d0427b4170dfae528bafbf24c69817907e1c31af4b63cd148c649607a9ac53bd58aefe846c2166fb1ba0d6dd335e3609a49c8fb903a3ccaa3386c09f7b364711372e8bffd671c5d3ee2fb3763b23e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h96a61fb32978ec464f2c25d09099d15c1ca2ff38e4e38064dbd8a147e8a8110f4887b79b9818e7f1a4668ff7e8b17552ea94427aff3157a3bb4d1e83dcfae9d0312b4ab09b0b26201081c074b02294151285394a732739b5069d38d6bcbae088a9bbbe7b7ac125ffc1e5efa6bdf097316d9a39f9c68cf36b07cad7b7a096854da10b6fce8cae2258f9c4c6017d43ed01da3aa651291b6ce0a44fb174c6bb60184e6c31e72c883bfd09b02e03486e1a8f7363102ec190ca6fdfca37187ce492a360d63ad6b46ad35c548f5d914d7b672cdf191e892ef413e5d689588bf43fed632661d4bc3d501918ac8b4597b9e8fd49b4043f5b7aad2a1d11595637e670d1df2455df20f9fa50c8072745d5b4284c64b47e6db304ce3e1ccef784ac8a8cfd25581477ca7243a03f74c44111428823070497ed0c1f6ed4c16d139f3cd852ba9f10a9c9d6864c8471f28e3ce8b629e5b555360ac4d7798172cc9563058b17967b0e4c300351d99e06c87dc5ff3c279d7e8e99cdc698293928990bec504fb3ebd8ff24b90bfe67c731049dd185edc22b9df826992c46bd16fbf32d97e99e2da4a847b24515bfb7d469569ee0b48f364454a270f98a76288b63c4a20ef87c3608a1b1fbda18fe5072d9f5d1697761e5d96b8d24356ab6dcf6bdc489b308de3cc6cb80f453614a13938cfa872fb56d956df60e0578464684872eda89dee419c488e4c97ecc154522faa50b3a6978b2caa2ebd9b403a58b43635f69d2efeacb9e60d8dda91c6787fbbfc36a7ee95188f4e2d7af02395806730e9a2e6b04fb67144cb048b2876f2610bc4faa3cbc439979b4c4a51c847d5026f415cd1c52c4b32a4769b0044501170e90e2a2c7b9a34ae4f5a21cd9954eae04c5954c4c05ab54b4c3511f2273ae2ba4c641f95dd604d6dd7dfc20aeead179dfb625d9b6deb947555404d9b537581027d27c3b887bbfda27eb08d1ed92992ec073da92250100a3fc71a20e0a6f8ffe7618c9f1d8bbf1b3decaa415eb48fd5f0bc0d3970a9b7cdca41c6441e38dee05c46a4ab8d22eef502a4dda728af77d0f0f2738a2b9afe87f2b05bd2abd5b6bac7f642956143218f34c6b497e21bcf04736f0f677c8ca72287f1b1b8c715bc79dde4330163e94d8c8243ef2d83e6c51d0b8b3c406ca28c5649640414c90e9d6b56aa074e2e0e39521f18d413c58838f653bf8dfd55beff5bbc536cd867e76d5e61899c90111e7f43bd9e8b0b87e074cdac06bf872eaf357a66e763d9c1f29d46d4dd2c372be01899e1a95837d041b7cfe261818f7428808c60c8fa2310ee0f29e1b6d5d14dcf844931d0bf00ff40eaf3293b1da3652848453673ce51e7e6182cf12db38a783da2e69183b97a06971d48dc7cfd65477cf098d95e3b631e208a18e8840dcc2f3b0a7d4723b00f96003c9d33b958ad54fb070fd338a12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h748593c8d2b758aa0dc514d2eb6ab48e1cff339ffc7bd4fe4295acc698a9e7088915207f92972133f87b3bc378a0bf0a2b9df57e7e1bb2a44a6020292f91aa8224b682d46d1099663f151849a4ce7566326ece1845457b41d350b83ba7a56317371b2f289cccb1acd840441d85791e01962051099af1721f296277c219949a8a0a28b2e3d46dbaec2a6d3b5896594e76838d8fb1c66decbc02ce266b50caad8551431452b413b7d65e14f994fddd538031c276485d114c38e2232dd105227eb6c30ef4ddacdb688d975d5dbae598fb75ac3c71111940ee46b588ecb4f1839c0347b6dff4aa7a926a6b28c81993335bb2fb60e5758a8981c776c121e203480d07ea3b9151254d3701cd3100cdb2063043366f025fee60471b8ead509820a053a027ed3733915c9c90991ab38946a44a3a467ab059f9999cd40972a0dd52547bd21db2047903712e55340d92cb119b2b89fbe5bb16adb90e4168c171a475165547a49ee76dfce2e0cd8dc9341b981ea05127f70e8b374be1fb04f296448fc78941dedb80b6280c775ae010bfec2bf7abdd6659673123939d3a888f447e85616f9d6636253b4449a8a1e86926c42d66de0c720f23acaafeb387655e54536099a0f9d7cda53004334ccef223878cd4238aa7775fdd9f407cbb8192220567c64d5ec356e6e0635a708ff9663d86b9e7ddefbfa752695235ed28519cb2b3fa59d0d19784599985a5d4540044bacdc95f03b02e7bc0c618498e3e6014b3d40578bfbf190c1332f501396b00df1d38e7e3d53185600c8f8b80690484f06214a84647826b7a0abdb1912ffbc092ec9e9128a557806f5323d3f3b9bd7df02d5e1a8da5084e65f4d280b4e3c8bb4460af078a0d19d2cfc055980988e5c84dade39bfbf7a3d5f3968bd65e47a874882cbdb4085fce41ec7b1ff13b8de0ad3548534ce9db1c4e277ed07247c60ecaf6b6e2e5fdce00c3e56f71cfbd306caddc2b1b99e817bc4bca94f0e7d78b14ccf7ee7d148c90538a58e1af2dfa9afdd41661852adac412198f0956c925b3eeb0dd6ea6e52e118bc8ce42e41b5f6f11732aacd4764a0c14219ef48be3203718d5b86d631f4e0abebc8b8f2d72af0c15697a1833b3173aa34ee939fc0bcf7333111f165d2022327529f40fa244c9bd1766912a78115e3fc3aeee5e6ffd78e4f0af715c6643d45f12a09f5d3708223bbf8e6e214b7a8b7a6549a9cd093de2cee4e4d1b49ff424b82a6e0ea82fea9b35997634f6e2c6e9bd5e7e35674c8edbdfda119d786e3a1c52f5a97f84f6266a6fb6ac767703ace543521d52f7afdd6122b91c1af45b312df2cdd15be29c725515cd04a1e580a899f7301a154dab813150746486bc02126c79d873e303d09a2b7461940c78fd5ac9dcd5760be18fc130108c83fadf06a4f4149c5faa590491ee406be9b5a8c4484da9839c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h92014efdcd094540d63a929d43e3d6c09243affb28cfc7ad6cdfa5af2f24a3d4c535cdb02ea1465f45f893965717b40d415d9b192b4dba94962938159debe98478923d6392164b96c5d224b02d02bb05d60cfdffef5af26227bffed736c08bcdcbb7b5e94a953827687c7f8aa2aabf1d66ec4441f5b7e11d6ab7ccb12a159e873b37df6dfb529a392aefbca8084d06db26ddbff1ef3955c3c6fdde48d1e0febacad542667556cc76a56d7e9aa49c25cc5cc8d21af181c4462fa0975c84c7a3660cbfb3e002d47bbc4209a43f1e0d4e208180e2db21fa572029a0692ab0c822193049beb6ab2d54fe30295b6aada9475a00437eb90dc205383f36c46d39c36a76b9573b23a36b91be43eb330fdbe3fc99f0ef8900b4f043c1c94075bb4d156e9439aabafaaa873489ba83307e62a03dd63318958b2830b41600bd9cd98bd69428423ee65f5aad469b5a76fc78dfa0d35541683b9724acffc6487c934b704629598ac83975dcdf43896441de76dccf3cfbfbe70148193de3b8a9d04e5fec12e8b0a6aaf417f82b9efa82288fb5cb6e0fa164f365188b64a8ce4628809c4b7ee814031b2181bfd391f6489732fca8e926e4839836c9444f34c53cb03bd3150f9eea737ffdb3187d074620a61edc05c762bed0f60a28941dff5fddbd542e7cea3ad8497652bc062ba9300acb7294dfc57489bd9edcfb9b585b56790a531955b03a1c2121d9d60770a074d66dd22220298b9a2b8925c1cff62016229670bb1289b53f3459ee5b03e23da73b99c56003345a901547246a161c59956f738911d5a522233d1f35e1cf7c2621e82b756d76586490962707f56b3b2493b7e8011a690feb334f8eee05d626ac5a233039cd9693372b03a2c934a689743b5e709ddfc9c9c43dbb1fcb2e4c2d40ea8bf2854d3ba09808c7dc3391beff41674c5a412a6af9dde4f12b4bb6c2ff1f2777eeee2e27a191ad8f40ba24b23f31c7179bbdecb042f60a11051a95f6dd48c447681ff09f7f24420a84efef3a650319650b5403038fdbbaa010995302d035844de4dc59318d8bb202f4f26a40ef0b182f51a1607ced90cefe071fdf310f831663c5ac9faa1a09cc352bac930b867b1e66d6dbf8287a8c27b306bbae91e82953ca86c644bc6abb8d23cca9d0d575b06db7e74d0f29f5eae17dd4922421de90d490557cfbcb39c2e7d9437733d1116de4a821a67d1b233c5002a22b68966add10dd9ea0c6fbec16009069c973c5af3115b6225c69418d70d8ad46a28240657490b708ef82f61504cc9ee63a53a60f390f6370e91ebff72639d46f724485c6eea956794b1b3b21df304d8d97011fd7acbf0def1b5405f40ab7b383512d299fa871020df7178d994aa652be4b56cf3f64010847ddf12c913aa7012091a75cf3462112bd3d7f8170931687b1142167e1adfb626d7bea8b394823;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h43bc2f09d0b90a1f5290a40a223777a6b3683e4d450d36a0308228bf9f1e0399034a4272a5057d481d07dd4d71551c99643b40a4515221911bb1caf07de76b19cfc9415d5c679766ab22ff35b059cac79dc78d37e3bae22ed370b5b3a4770d11fb4b74755f29058aa76f48b937df8b9ce1121a2fcdc913a91fedb53ef388b46d9b7b36024cf33815dbbc08f981a905e4ff05fb15fd30c2c4cecafc92784c3b6ecc6035f9889ac3efe9d44d68e4a0b1d10e1f79501d3b6636df8afd4d4871837292c9ff6ab04f8d671e55497d87fa0a5a281f7b8db9067f6a0367747647d665891c5e516cfa5983aeb31a3b69119bfd804015700d50636af793f153cd27d5f91b5a47d932c1217340de3f536e170b1a6e04f937de88710420bf639b951a86bb01e6d4534d2bf8eacc3f92f09831dafb5c246bc6098ea584a1169e644e6cba9e6ba90e35aa3ad3e8704b692ef9bdef338a5b901c83cae5db10833c5c3de0db50c278d57e807fba08042fd1d354dde836192bb18523446c94663f6ab877319f0b6033ba0896cdb8e3e2f6c79f93f398b5e755e2d511bfa46a3206f7be7f55d343ba0336859325436d9eb8c7043e7008b77685aa333e26957bbd7662aae8a064ab40d635993cb40de28356257d45ff75e9528fcfb81d93e96c0061e3a2e879d99aa2b11ec5b3cbfd4f2613522aca04ec617cfbec5f7aa8d4630e9d5d45b52f971b99b6885efd9d9ada34f1d1f2a3ff0b8375119ea569360dabd6dc0e8eb2223b836802b0b0d8ebe65805085607fa8f167986f4f94842cc29c5236f11fe856c9579f69c8a25ab98f6acaad0e82a9d493aa4cd25bfa6ea1ffd80589a2b8cefbf13214367bbc489d913fc920ae123f5061f00d5df02118ff7e92fb1b5cb961bb1e8a2a41ccf1c6c0df20d1b1fbc71ad81dfb0228b701076bd6bf37f22241cee534c50c2bd2ef7b11a22936bf61ffc44e98a6823078ca92d2409276624ba89a7b9208399c70b6a2a2189f5499d635f46a24dcd33ba5b15f93e1b57c67552808a6c234fb3d5e859d4b468700fb1e1c51e9fa66a62d5d4664148e8e9dab99ce479963a826c452bd8494102db65e1c102e3dd4cae8f054e8f97f13795b45982e9455a014ae83a39183ca9ddaa1ed80e7123d691d9daa59036fc0b7c17aa76686c1dca4542bb552e06ccc5cb507d0c287f3436a091807004971a5a02024bf1162a1ce9956662037ac6a876ae3964983b6b11a5ea3c1ae322f35b0d0f5b21407716532e62d45f7a2c74b139ced57d4a0e6d66276d36a1448d48900a0caecb3a0e7c409c9be3d02920646058cf71f2149e041430b4ab8b5bfd0bc11e3f3e2baaea241bcaa78bb87cb47dba9ef8c5cffeaf4a0893e85909307426c0c70d0a46bd33111453bd281af4ab451035bff33eff0a9af3d55649331a4f414ef0d5c04cc77a730ded422855;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h51bdcfec26c798214099eb3fabceb069b4e49283adc11d39f0ed0cd9a3bd396b01de4df6203df4255263da8e946375b1deac803eda228fe6259a756399b8e0f21f1bb2fdc073dfc7bd496ef79bf6ea24eca4270dfd1a6adadf624baf5e95a9fa70843fe5f98ceb51749d78203fd84854961689a265504641b21214022cecadff157733b24907b6037f2c44e4579826efb496d3216c8ff9f513d2bec2a9bd2916e0d6be1d504ceb4e500c452545627a3b2fb2dc278f0c7d55761eff0f339ad5f60cff20bb8846858fc425fb11aad76df9a56564af395d238041ced999f11f87ed321038feef84c82438d50ecee6608f529bb9e2ec17d41338398cd58dad3f92e95b610967c19334463dab5afad856c8390e82d634fba390699e5315f8234332a2a434e04a9af7472747efe2453d98dac1e794ee08cb99dd0770351b01af71e2b326f726b67d21f437c66f42900c0d4b4b357ea901cca65b06a9b0df851402dc4afb18835ae59821607940eb19f8ebe329588e9ce470f821f78204b692dbf7036bf3610fd9915b4128a0ec12df632fc116d46eb8d7158e148e6ff565aad911327323837226cf5176d71446a0ebe4eed7bfbf6d69875f59ba8139613b16c52a66d2373a94082465cd07122aab23680f420c5a12ad76567008da0c5a46023acbc3d56f8b1111e180e84626eb7ff829673b7bc905e2ccf989ae33fb94a23261e03ba88c605365c2bee95c4f551787a4961a61bd56dbc014f1d1e62d859085f3dd5f44d263668b63ec442ed82f135df4c54fc799e64d91b046d701f7a770344fc15193fad9de66d47002634f7efaccbacb5da7a34ae604c410007ec0bc4aee3e7170a529588eb75c4258f9ad4a1c5d0f0d516dd93d81babbe08919d8756d9cbaad7a9759ebd759773d2330415605a43a43f8f8d44561512d3c6c355949a9e89998eb9b82e9f2ca7aac2a113122e0fd29c5a711ff29f03de21ce9d7ba304275682a011d5c811d5eea5faf2f7771d5cf0e33961e69026fcbf6abb662d72cb53dd8ae50dd1d6435839d55d3d5ed91695b64b2ec2b735c36c363f7ab82de3436f216bad868dcb642cebdf8f55a96a33551915981f1356773d4c426f554b149a00861d24e489c91e772a5d295d4f927b0860af0bf7d4c7f6f4d31d2d2578cb3873a058e24b94c079b879af8670d47d84d9d2903f4e0e17cb3da8c3f5228958977837996e127afad473f3ec4ff1915977723a9ab88255c7a5421ad7ecf4b46fff3f38b9794b9ea2c9510543b01c73e0167586c11b63cf517d72179bce8a9d258e1faf64b0cef52a3414178bc78290403e0b1bbae253854af2394ba35078acdacb45042936aedc81406c1b3091f9f746743febe00222d8446e814e9d054c36fd2574a26a418c7064e7957769629c897fbaeb5284fae1299b3ff32108479cbaf82a2282d0e450;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h78ed44152012c81114599181bfe2709e349cd633e73490e1279c47c3a5e04b604a2cd930133452ae6623b36048062809542d4711104e74c2386cab29a9e65dddc963a1cd5bcbdcfafec1f04b030f6977a031e65b490c04de4b1d17b37690b19b0a1eb64081ba03b15074008a6b3835210689da361bbf75825c5ad74f239a730817aa9846438b92e2aa70e0cea33136acd5ba82ebf52ccec0cc48a04b70c8983b050676fa25e0e800ad17b7f6a19cac8205176e6e4df272f30f3264b608c0ff63dd7806a16f7f1bafa0fede5b54f6a942ca4bd6efaf67679dbc52b8429758cd5070c8dc7921296a8a21c374faf504604deaf00f0576196fcba385aba670050ba2de6aa553c0ace31fee48bf935fe73820fb9b971068fd7b87462bfb38c46dfbd01900923b3cb7d3bd87168624b4f03e4b90c5409a48ba2e8c347154688fe4d45315a3b5702d8bced09b04a82626ea6326133ee483a2976e96ac0ff0e3985bf201700f01f93b042b7fa236dfb0328a0f5e8b46371b834484dbd4163e08daef71359f79fd7d5457febd87054d4410c466da90c9e25362e0edc98faef422f2db43e2c697c83b9d51542b78f0d8817d660a555ebd5878a225f350e485c028cf0ac1355eac9d6342a583c3dfb5cf8b441d9f5113873fb8ec6bb175894942b612f6986dff2fa3f2837190acab97ecfb771a6447996845d27abbdce722aad88001ac51233baa189626e5c73424a3413cc47ff88a2ba728747936d41f0eb25a39b3e82084947e5a8b5ece8b3eb890903269e1f9791fefdbc707f457158d03a56f09435df670f1bdf3b75634b5c599421be2c03ce5fdca3b5d997829092f864d4e04ca3265af22ec90d9a1337c3bfe51f2d335ec86a4ab5a9022ae2ce4e32266bbfda7b35b5b30e2ae7e968972183973016be20803c0dfc4a3e8f0ab4e81767e9e589943c027246feba1f197c096fde89d9d51329b5b00e49ffdc48e96c83102c248d70f59c47054b95156b4155bd248175a2bcf1c6e8fb1966358a95adc1e5480fbd2b46ee644a10b396f79374cba566a6093baf297062d9954e1f02a248787dae2c004a371d682f75888199e498b047c0b45344d4302569cd966120b002f6632f249ee81128e43f568b60ed43b7af700e88839abed9ed1fa9b13012f77c4cae699f88874ebecad6e5115d771db812468d1cdc605708bde5f7b944938a81944d8e51162355a52a1eaf80c176dd67a75430e1c4b51d53dd6594b35e54c887ddfae7bcae46fdcdd13de7ffc0f610b5782c6b3bbcbcc531806223e5faeec72694cadc8906ef0c9051e0b30e87dd0f74b3ef467219fc750c46e5316d25836320e3f7106e5b90f47207396bd5b8b8795b7f70002d00e35000d43fa638742249591d5f6239539d26ab3fe9a97c0265614b6b8152aba8d4aeda4dd67f8b296c82c4d61c6a3dfff1d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3475cc87b1db961845a1f6ac6cd38a3447d94c1ec83b4597c6a29275c646cca3a6d57ece18cf9e56db5e84438b3b2a9c55603f55c9196d12b9598ed79f785af836e258adcea5b0ed28c3e51039fcc79a98af47c3d058adddef89f7839c74ae8eb99669ace1029f81ffef5e15d06edee55c5b2a942e61c7cb7b021cb91132d4860f7a3b989d75805cf93c3b81024c94b0d17f5f49da9074fdf6590cbc7a2709dcf0567ab6d08898fc8538b86d0cf079037b664f5d2337b59834fc73f6c5e5710e69dbd93259ff7e5ecd932a1bfa2f7c9fcbea40f03c48b30b331023795e9e8a9395f8ed120223e113e895f757d2cea3c4396dcb67846e8a19fe8ba0e582b5f312bc4f7c8bfa94692b0077a100293e371effe9ed87b844ef5142eb91edc0395f93f33fc722f6c4f8938aa4c83c8990113dc75f7a40d7f420ff404e210dc4681b3338bbfb58ff57d7283b634d4bbec0409266653c9e09a152e00bb3cc431822253c7afeb81e361ad0e17a39040fd5712d1a10db6614d56f2f8e2e17b0eb2dc9bdad79b46e1d711a90ffdd071b904e28a93ff90a3c3d0b0261688e3aca807e3a0b42b689214a75aac84357bb68f6af5463511b48f3eadfcef5824647f39b9894174e685284dac5fb6eb9c7fcc608d3c7ccb767989ee9e188e873f201a8d375586372afd7b53720e05fa65214fc4d6f813b8c8363d2e57806a50b993183f1f912c4991ee73b3dc44d1f01167be4647bb1013bde9c13fd880cd569c986365b5bcab88c45d6447de572a8f5e25f064bdf8b25b47a6209b231b5ca899d4b1ff3e8cd76d3e35e92ded8549f0dc8e65212f943492f5eec112cb7b4026575a925cd6ba87dcf0ad91d6aa4fc9b8f1ac472b631f1c99a77afc4917fb911abd80d1930d2764b76b454a154f0e86b444adf066dbcca9219c8b80e65c526c0c8ea7272b66c61b5f4e698431315b6bb0c0d2ee60033d11c53215d22ebeadffc31f809a2b57049fe87c857bdd47fd74a4409aa1b2e0c689c83a98ed1a226b61267f62435135c9b343c31ee515503afc664667c45b52c9d4096b5a5bd635a72ba0a03dfaa5baa5f313567561138d2e3caff9156691f8b36f7c1888b3044c9843f74cdb31f73f5282b6dd085f40fcf8db330bcd5bbb4222d4b1bcada15854ddd9c87ee141c377a583ba527c8e715a6e156994d736eb164fb694503e7cc6fee5a50884ce32192405181ae88fec40b8339c94f9b0ec5fde130eb8e385c5cd983dfb534e23f51fad10adda284cf612d243fac1768fd34d7bb1dec3ed59dd1a3bfa93f9b96f701737eef997a1de9c25732e0b3a5e86ed27f02467b492c0cb447e34a30e4d791b36843b1aba98c8572c7c9c6fff9fa283b287a157e527a486e70b853e96ac04e8bb562f21512732b04637fb221178a0bbbbcfa3d53e9a70bc35cfc8a465863fa5d995a48dbff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd4129a4eea7548515eef00c43542d2c99d03a909d06cc665619e76e1ff0c69f46000608cf5531476c2d4741e350128f49225ed64556cfcad01a77320b9ffcd869a26091e751e950ed2d060662f0e973011709f5ce3ce3d24775f4c2c41e21e8418a491359069423d78edd49d92b86a586365d6c21ba2d3c5d04969881b350da76a7bbdc774305120205111cbd6bf94e355a486912bc0c8a79e0d2ca8ac9da1c25639507d593fee6377621f7514eefc0b4b4e860ccd7321df5d800dabd729ec6f3384a104dafd52605154c793efe76854ef5f98c5f7d814014b77bf3796791dc73ce4404c5c4dc9687c0a9a5066eddd966cc2e99757b9302fd6d9f317232df056aaa969b7c412a35bb2df8e5e3b943cb7b684d1a203a3357b018323c94cbff1e0d71385f8d586b63700dae05e6bfb811871c4ab0fbe79b3c0f3d2690cb11205dc47ce9a59f53f5b1044da3c1afb6b146ad11b7d37b9910487c4e940bc0a375c4a63471ff8ead67a679208c3cc00da74f2aa6e8283cf22ed296ade49e900bb3d63ef8ddafcce775abb2bdf6b54c835d77be69e2ebfb728dee6a3c3e97a4a53597253c9c40845d90137739f0a56874829be5c1aa5f1417945e534fa2c48f7277db4bfbc01c7f76d0b6e46c708801b3631122d4e81b73ecb173bae7cd17e19af32fab724318fb764013de14b897b885aa6ee4f3c4a74fd78c0e740ceb8e3b03e6318f1dafa4d066199599bfa740d1e223d24fcd0a61d840451d652428d932b7bdeac59ac07fc7c4169fce8920dc19d79d66247a3b7737c905524233d2e59daa2a1ff11bd43b404c44954da03ab7884c07b220f6b11a0703a99fe11c94799e2acc246b5a9e5d681e9be138410e50bb4165104915a9efb3674369fe906509cd5af19e32f287dc5ec3a9d637493ced3f8d4cc20868503174cfd0a25562ba16bc6fb7c5d43f32cec4c102d4a5557cb6b0c9a153ebcf0025de685ef53bf64eba6abed9bdacfcb78f90c92e9c778b5f01fcd990e05304f9045cc3a33a7603efdc6ee12f1f2649db2a9c691b9991216c753510d3f5743e8fef4c7f82fd726d24048ecdde540d7c82f946716f855f4fd1bd89681e73da14b3764fb86210d48be4e40a441a9da2faa6c9decf798e361c1313d61fe184af5df95ad17ac29bf5374e4271490b5a3010afcb046fdec320fdab85629394b2065b4f37dd98f19df85cf9a0067486c895de572ef5412e121080527b991859fbfc5effa28feb8a17a2bb3f33588debc703b7a66e7111579ca08468ad690a6dce3beb451a836b60910731979b42def270b13a341bfd01200b75d22b199a77a81404be281d199a6c3ec4f631ce683718dca95eb0aca4dbe334c5831b0100dcb282d2cc7ba96fac9bc199afbdafff77a5e4b2cd70933955e428ef142d87b7fc57bb7d0993bdec84993463cf17d1af9882da;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he6c154f4e2c8ec08d84dd4dabe259c3e0554e76de972194f48efc18f9de0e79bf65afc3ecb93f82390abf8362ed1964c2f04977dad845dee95917984b44fab81fda723bf7092a1d4ca4ceb5ea96180ccffccade04b3aa715778c2c80ff025bccc9c474c36e8d9af72517e77f7819a1b9feaa90b28ec077b50a159b4d1a61cd910ad8a11ed64e18d9bd76751921057a2d3365cb07156b5284cb9a4ea674b11539154ce4892904b49aec290d9124ea9e56c00d7dd89870e5f7e193749701753e7144046f76a152a36cd9ce2e0869b82c545075b728aaed5ca44409c5d18e79819533d2759a76bc338b8f4497fe5a75d898cae69df464062973a32cc2b81ba98953f41953d634fcd756a8e38771311c4daa7c045490a1f3911678c78b9cd6ff39751b5639f5417b3bab346101253ea5d4f3bffcac6f14e691b2ea7ece0ecacf86f6040d0d33fff3424f09d790d6f63e8c46223ba216b419b3ece9133c77a3f850028da48d101c2b3cf7a5f7327301e749b3c88ba4e1977ea62f245a730aeef04f5e2eaa2da5506226136b7fedf19ffb715c3f5b1ddf651bc3ec45517d30353d3ea04b40a42f25f7080f181dd1a2dd67fad2cceee10f9875a32ca2fcd24e821ac8d9968023cc5fd7becfd66ad7f1fc25039487bc6dce13699a7d5086b158543330df3479f199ac42ad07304acf1ba9fa6568af6622cdb69583ffd2ce0bdb6875dd497da94bad93c6ca6d85fdd02720ccae9c5ea79f16c6c9b41288f28f83f2956b5c3a10eeaab6febd65597842b6373a0af49e2974bbea06f8f19e9321577003403393e2f5c64c029e0c1db855bf37bdefced6915247af9c2419173c3ba0c128134d7d4d93fcf724460a742fe43e86028c62492233b8d740fd1a2d27fb6026a261c49583454030ee3472a7fe35247caf1b355ed069ee38cc2fd6ba49601b2321121498e128fb59b991580e9cefbe1fbd0f467648ac5fd9ab38bf3e0d2e898123e978b0e82eed6a8d38a2ea7c6b8d3ec52a427362bd452da05306972a076f7e48fca57821ee43f39ab70373e6a20f5d7e534c2bd4ae80f5419c77171caaf66c6b60eabd5357a90aa1ea6387245cc6df7067b6b5a9e7cfe28de964dc21c1b62c4b9cfc77efa4d48e4c01f7b4f7983c6f1fa47bb931133d007377039a57d555c0530cc1b39f14d30404bbd601ba53c83bcc1ee6de8808324f5db87e58c77147ee606df3a3f0b4bfbe9514fda9b60de6facb889716f64cdd2c4809adbca60bcc993ae0f28c1705606f45b8b03e69022fcb09ab217c2b69f7e478c82c3328b2fdeef50a91fc77d2ca2b7083d252c0fde3f5ee9724bb57d38355a7151222b9f328b19c6e1c1ed7c8d70283149c0a2c1d5432aed1b6d792d66bd6e82dba176420e175c58b609d4798bc0da6f049bb270e3257d05236e5cd909aef6711a06c63925ec80fa9d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5b2596e4a346a4c8b6b2aee2c3ec91e36c73599de6d4b4b1c4a11fe07394b5248d4f7692aa305b4c1fe5ebaddd826e099a9e769e1b1784329eb0c69c50973a9068d887ee925aca09d1ef28e19ab2dccf3764015e9afa30c51643391fb58b38307b6d78452f0e7dfe65651bca9371de46b5ab7c74a0d706973a7926480cd79d6cbd47c9f17e9aa46ba3ab59a3b0b448f433a213a723822e0270b09071c3bcb9acef9efc324774a1980dfff91e7b7c511b090e6e2666cb6bf6db9d97adec38692aa997bb53651e5ab6c55cf5ef3e269175c0a9f85ba13e366506f6435f39af1f228dceb22943e539b70f50ff92578feea4bbb56aa5009b4550ab6c75d327c8fd5015e81896348e4d2e9fade3e8eeec1bb229de6152a5a9be227c7a9bef8d5c3897778ed2e9a586100fff53803e09a838afec318b59a1535db9ff47f263f461e9969f9fae69f6572adb181572caf7aa4b432386295868b7d1e89f8f8afa64d1dfa45f2defc417c056a07c6ce96593ad3b3a5754acc258d144fc1da550e00bc3d6f34b47663575160b83df458bfd8a768572daf298743f29506ea2c77d37bee7a273db4d67ee3935f7d7af7959c81c1b66939cfca2bea003d4785478d60162f818cc4f207f73c15657eb4495d3fec330f54904f88359a8672f387ed4e21368e8d579ba27d1c25d4d87a41e9396d5c24e644a729fcc5aaaa94e495d445702fb86942737506a1b6f91b0b9e80fd53cb150dbfe3fc0a328caa0db24284f266477f05a259da2fadce1666d558466e012d5fc0564c2445e7f0bd609aef21edced2aa66682af554a27f19219875b24ff270ddd83d6c140b29379ee7cb7fcb9485864a76029f0be27c194195697c448c19713729b22716ab30ae408ff2077d21f5bf74c7f68c361403a15ff315e56412d1c88f9ce741d25c4ec068e3354a5b8adb274942a1457456fa9dc2dc17147433e9f43b16ab748a75184d941500941266fc29d0cb85db68f70d9a807fd156d0ffb62233940d8ace49e7deaf45c4c2fcef6c3748f1bdc01ec0750114894d8027ca4705ff5ac256282746aa8c9df20dbea2d9918452076bdb1ed7701b1a050f3ec90d255d7285e886b5037b19aa8fde5e7d234bd3d93d4993eea1c190d7ac5b876aa02fea430114ebd69250f96fa85a22528d1fa2b6575e28cfda93cfda532aaee21d14e2c05415a104a70fb5255f0d612b332764f861cd3bee1b911f78b34dc8d7fd9d7bb797a8fbf862a435720d39ea96ae73e12ee28cc3a0a00ad738cd3d9386bd9dbbd91f26182cd03bb55b76b35af46b97e40c63ba525ea78ae625b25801337eac310faf5d05d7de51486f49e2a169b90b0c4d53c4e413dfa2f4b46667970db5cf6aa7b714428ba993b3cec718b2cfc84c9ffa5d105bc3cc4a112e1c9b7632538d29d18b6b5f2fcde574f9bbf99998a2dce297729;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb919bf489e271d5c87cc995cc893353ce3e061080460c45ba60f27dd96a6428b55555782782204d2c9e0e47ebc48e1a7febcd1340e2d9b456263a16fe24803e572adc7ed99bd6caed0048d356d1993803067169028c81032a49f5dea4235f8bd9cf18467d31f32febd437d3258b366caa7fc8f34d6d6968a6ef3534168f2c08586d44bb5cf8d855493e75f712ffd4d479774cb1feae1675730f32a913931f4fca4e03034cd828172d3c2b55db83455716b2a7b8ed378c5a8f78557dd26b9446b14019036bf9dd0e9f4e632f40f5a8f8a3d7d5ff90453e3c13d0544a93afb233e27ed79b32182ebebf16d998b9d59beb4cd77aa923f72ea0106776947c6eb40dea63dce6464f629daad80024d913bde88841373791e7ea611698b829f603a84cf2939243ef6a7ed01d64faf06e0c778a13c5f8e719c7a15e4a6edb1315eeb591971defaa685b1dc9e317f4a31176d75a0db0f76a1523feab0824eafbfeb18d40cab5805d44f8f6a97def27200ddf7c4dd362e2978d9926f32ede05fff5bd965db1c4e6f124d64cb2763b948fa873021490ea21d258f1f290ebbc098a5f9c118ee456ac6a0c3aba8519aef20a968c3dcf2ceff17608e805034c3308aefd670f7e2adf01eb7b7b5c5de8cf484d30c901924f6ae6100c0faf838e5a8b125d6f2f431302ef2657b74d9246227b22b5f0a4b1b574e01efa7830798f480ceb762f061453a334577e732a9ca184ea319b66d8f97145353f874ef00b41f794a47fa5b71afb2c78eb661109f158b6960d35b1070cc8f2e979b155b5e0a0d14f7a9fae69019629ada174f76dc800ab00e8583da66e8ee164b7e946d1c7586e8877c531099b2979772a1222fee4c088819d3a40a3850d095a15b9113e80721a6180b55d18353b0154c4e97fcd1c3870f59f70c8e0fe359bea64323658820eefa0c4381f71e5a6902de0b9e93cb87def5480539acc2aa061682b1ff91249e1f85a63abd9fdbab517d9b0961bcc97317b8276be19c62d9ea569378774e798f8631b974f0df96d21f7a90326346838929ec5c6817a331b9952e6c2245a8bbaf253c18a80a01468807d747eca4a36ac4427e153758c2286ff7150e7913b3b131e58e1950638ce48bad7db5b95b8e35c132fc2b3532e67db58acb6303e2cfd107a34efa858a69ee6067391a0348d0f4db146595d1c3cf18ab571add104edf7c35545a398addfda5a799318ad9db9782db1ea37cceac530f24ca6e1215db45c2b7aea3961546b6ef4d369b803f755d28e710956b589b2047e5f02fd4139ce2872614002c95988c10b2bf1f608b6ececf0e62d67b1a576ed73000836167fed2cd31c1323eb6f660e34fc71628d57240d3addab527b0c56876bcfe1619608dd27098eb409551711a76b4543f42ef20338567a6d82661d3bb9338875b6907e2dbb6a86b84bd4e1e5df8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h71941eeed9f23b866ef99886ed8ef9b9faf298a60e2339da6c6fd0ede32185990d5d66baa599cb915b571cd6fb1fc968c384d2e0017ad716f9274f3ec075a224634536ab979ec1cce04af79b2f6b9fa45c6fee310c5e5634d3927e838599ec799fe1fcd99d45a20f2784e03e328384eacb44d66adffe91c509b29e574e263fb017a4c92483064f8c4e9f4c46ed073df81c17965bdda103c911d84791bfc2bbb5c95da3e62d8eda58d8021d869b911434c39780dd18d5fd415f245319b8fb1b180d7ee4fb07a077b984fb0afa482b0975688efbee07bc816e5e433a529e82b49d6a84e7e0f6159e1b46009bb012af20bee2debd99a8edb193f0c7adcb6ee5c12f3be94220a2507ff3b187e1ec9c14bba498e8311fc85da41ae02360cf8f4091ba3ad4ab3f93e3e9680e209beb72e3f278cd148eb8cc6f64e600b5573e5c665351731bbf8bb67cc8985b371d02120564d1ad4dae4eb99e03efe0bff7ce1617cfcb23151f472371b2d3945fa2a8f7d387745aa59d3b9b46d2cdfe6746e19b51a045a68349381e3815b1d49bb6044f267fe4f54f9a7b8d94282e9e57bb3432eda05f396cc15e55608f62035a0e451978c75407cfd4da8c607b77ad40b8aa52a210681be9306eae229dbde2a3c8b7dd2927f915c84bea79d9f7818d746e3fffdf3fa5cd4ef158ccc7de0cb6342686ca8588bb8ae926dead5c3752b6963273c984357d93b41d617ed1599e0710f2ae56a3b336e7ad851bf96444674cd23d9db6ee7b0858d70f31ddc9a7c45691c77b3bad6a248affc135ce259cb6c3f80f54811aee9cecf481549d931e104983470af3c7c121e52e30eb7a6825b3128f710a57e4dba84c24687b37a3e6bf70b6a5796857b4462d143a0a902b8bb63a4ae7887cf47263e1dfd96b5427f7dd444fbd882c77bc2b8869559c8b60278a4c3eb60ee8b340543e8370c0bcdbf6974683225edb2fe5e01ae20b48f922e0153d578eb09211be0032058d53f93850b0e86b472c47a180869c17290f2d48cff03d0d6bd3e89a6ff9c303245f7400ab2d77da57e6e9abc194ec24c37f89c24f4eb04a72c95db8e7ade217a3fac524025d33156c5a30d782cda09923e9b30506d632436301e372e3cc61802b84bcb96daa05521994d79edf809100d87489a1d5e2d7c8e1fce004a5c0b8ca288dfce4adcdb2e6b82c9882cd34bbfdb25afea12108c9e34520480b015d8be3f90c4f64a40b912a719f06a5f2636cb9136d6f45113fdc4cb1ab7f28e1d386d349e195358dbfc0f6855c96babce6395a61268012cf80e9038713344df62fe9ddbea36fd6ffb74fd4bbf39fa59d8342bf00fd618c2c5c3b67c2b38c2e93d67ee401c8d89ec7ec0d29db19fc6878af9345ea296ca361ad2b7c25e7a808dd34af751b4867c9aba468d15936e19015fd8df6a7cc6e01122d820a242ba6a449ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9babfa798fabc8da811d3e586f9b2e69109e745c3ee874a8fcc54720dc7fe1569a2ca27068df94a0cef9381d41619f28e72a3f9a2de7f1710c93f4f4a3d98fb226c72e286e712c2af9e1936094a2cb59d2bfd03ecb2885b2762c5b5cc70baa032bf4f809d1e48e0d59e7d36a6b61302a79b1c18de0791683aad761fbf814793fbd8b36a5dd1cb387c4cdc7bdd1f102dffc71c68773b0c33dfe6ad1056b5fb5f983948578a250be53158b11a0c49866d758ca5bd37ec22b1869f2a6a0b881c9c2812a12ed8a64d00cd14a7c4f591228f9c39a996bb922a8cac1ee4fe5501e19ce9a045431ee5889d740b45c234f979d3d1d956f8fec86c93471bcea357a0794cdec5b7bf8651157048d5e4a09655fce578892e626d18f2fd1c6a31199ffe81906d54dfcf5237019eebc526796aa46c1b65c0e36558fa493eb28ff9262ee891152f720beb9a06f1083855d70db875552e7b5385ae7e6110b2e13fedd2b61869dc794bfaa32e57163390bd32dc2f006cdf844a16b5ad8265f4c8f6d3174a32f527ab085a2820957cfd1c4fd368fae4d9de91a7f44940d2a4d8c39817bb04dc226f7ec753daa3ff3ff003f1d3aa99f1becd72795f55b28c1d6c9f0863de525181a07e4dcba838488334fd128ea47bb4fdb1deaf9ac1d3411506f663145aceda2b4d42c8c2adb0d6ebccd9bdccfeb0463d79c28abc81d54a7d0f394a2d0149e1b702e0455de7b6001b3d8ddfdaa92ed27e0870f05561c3785af4bcac4cb1d1787800b9a993cc10bf6963b836ddb2a71377b190ccf728ebd4e8f76d0ec0a6aeb2428e16c77c294222ab955b9cc23b538104304f944e06336f5bd593556409cf473d1957fd31518f934af428f5b01a566160a7cd2c97e95634e5ffc377f0f648fd3b90cda0451ca04b9f46633c42a16858b8f1bae2ff015c977017d55ca18f1f2769f1812912cf5610306fbc3ef96801f8d051748314933efc9825c9147d9807a8f4bb92e746fc4ed24d99e3b3f585949a83181264e7ce8a66cd7efe58bb5a35bd9cc4aada2c23caecf6b67575863b24a20faf84412f7042309356710b6dda6de427b43238c7bd2fcab6168f9a811cc2cef4a26f8bd573deb96d945e642c6a4f8810f96580b3cb5d45620255cb68d3e3b7ec01075a18a9d426063bb6e820889797ac2746a43ac8fdea5f036974f07a50f75298e54c5006c14ea77d80e4a4fb582551fbfc8f37a477d6e363476d9e497a573e640da08cdb0a24b799395bf70012cdf2e2d5eced21d388a8044d1910f967b03df7a7df2b3aca4774674539997dbae29742a1402833b59f062e007a7dd0cbd134e90a60af5f0f116be23996df7b804957d62cda70c96b9fd89a1109d60018bae8d65ca3b1a3322f568ca3f1f28f035dad37d2a403875c722014877c41e85e38ba999da289fbf20c5f0480b3b6e86aafa55a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8cc956598cc7713dc9d40123472570f7b0269806b6c4d3143c049e3050c91da35c72b6e0af24b8d03138815db7f661ffcb10afa9881c78cd65a00da5f8eedfb11d9e40da6dabc7dc5db1b9925f0c282d336a4a622fa6fb1e98fc9350891e7064ba11a21613ae82eaeffff7ed8839afeff92b7cc3dac05ff453b4c8304a963db7432d951a181e70ad787913e8208d5b1e1d9231ff88a94b266331ca0316cd74a3b29f1ff17fac41ff135adf13309f1f77d3e1af493c53f0b5937711a5c757f2ec2728fb70012348ee0cda4ded876d6823d7bee6847b53a33f4c6f68f3906b929dd01396ada00defc32e210c168dd08452ce7d67c49824aa45a1e92a1306d82da2a06097bfef139bafd7728d0fd824b93ac3256c380fd30939f0fe528719b6dc6526d121c3b838beb890611f1b03098516197109c30a7a19f8dba4bc65e1b3b9b6e4d5607767c9c3c7c1bae20649e34010ef1fc9010fc50ea1f036b1741d42ec37ba5e1bc8071fd4eeaf5d47f703bfd17695de329e56de90da1fbf98d6534fdb74240b93c047c82b36d20410f60e1f739e2bf9f9ec3f3dfdf5f2e1b47e4d42418d82e53016ceaae18e34d8abd4a7c8464ee1b39cbb3f23b613a7329f23fa43c486de83cf111e341ab129c3566b237e3121f45d1bfadbb474b8a5cd22fcb1bfee65f910ebb9e5443712a0c957682edcb6cbdcbc1e36613810d7ab2f341c662c7916ee52a8e76431066ed908bed91f055bd2f1c0141e993e0def8f7cd37ba6c7b6631d5358a47c1201076b4a9b870ddbb464dbd9e420aff3554f3c788cf3bfc7bd5e0c96b31060476c3380b54bb83d5279c28c890fbbebfce3d507f059183aeb43686f591e2b6c39fe10721d0777651d018753274a209a97226f19a5400c7ffbb43bc34029d70cb3bf1cbac631fb2b281427a8b55628207c9eb98633bc15438ed138dbcdf73673632705b2146d888a5500a65a7115fb4bf846ef8cac7e724025f8aded4af966a403163a8f7c51089f452f0fba06338a2fb696a087681ce01e02fe2b71897f1aaaa0cc22ea63efb581cf2a1af9deea22e78cc3a00d79762ceb7e3623e69c3cbfec1b80521ee6bcd73277a6420963c9b9e49d14ef49a30c45cf1bbde692320f368df23b88d7e18381ba8ec3b529642af4a571d0fdccb56b82ca01393b2dbbb96bdab6a8d0818d4352066a478473a857b85625c2bbbc51b9aac9bfbc8cab2f54b52333836e4d413cb7c99f76315372332146a562c916f6eacd2a68b3d780e6f269746ea33269fdd3ece1ee0437165e7095ac464a947c67b8fad9618d4482422b8c73e3a96760eb4ad753a7507e0f70a1ed1ab39b02d1ff34b2157072c4104b72993f949ed55c59984d8523a2d2c5da88a936b2f8265a43e605f7476d77a01984d7f430dfbda5f6fff913ffb5f89f0b21c7cb1ccd7aafbe115df8704e7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9def5de64bed7e89a218e496d6619234d5e39a6b47300e5ac5fa5eb9931c6c562f245f107a1e7b9ebb32fcabdd1d6beafb2098881fcf4c44e5f0091e196dbbb46f9d26d4006cf69290efb98559ffe983f50c44fb69408fe92ec690bf1ba29c4790c22364a3e01be83ae61dae988de55f6115eea2e2914efaa8ac0286672318bb3999e5c7b0cdcc3b62304f317e60d8620129e096667adcffe7f7ee3fa4dee7e267a8ad3841f15acc7d8a72533568ddf874cfbf65692de463ced66ac50043800439a5ad9b18e09a140fa925397decd61dbecf35f273c13218cc5a1ebac89dec8874d68625327f052713c3b08462d9d2f82c80885bfdeb10668590b5cfb8633b138e2da07db490587f9b1a00875079f7a4b8a67173cb5a412b15a82c054d8077d2940263426eb2b307b97f870e6eab7f3a139153c1b7d21cd293084ac3cfa3ecc10b7e0cd1d7711af84b2b9ed8998843402ad1a8a7ba6f46c6ac6ae795bcf010bc4ff1c4fb6a14e1fcd8873fd04c61cd52d0ddf4c4297d11eb8a545d1639d3e25caf9eddc89090494bd7ed6e53947b93976391c89dc3d9719fc084f82d8c3ddd8ad5251267b69be09f12ddd96fa635ba609c3aa33310c275ece98b8883d35743aaa20ca73c7dbd13096b54bf037dfe373ba54b2e3e2dbd4e0fc4dcb26d617c5b2ecfc83ccaded44328af4fa7ed71626ae39d5d194104d29d84a541faf186fb791646d8ba74ab66125fdcc897166a482b80f52a149ff075b6e06bedda0b3b14324ddb0979265a001fefab3dbc9006f082dc519763c4768fd48a2bbd4d11658239ffa9b2ac8eb81371243f69be76afcf9dea2b05daa33c0c8c90329da8a3a38b6e44a0b3027c183879a318fd81efc7689ef13a889cdb58ef47db68f96d906442d8800080f1c9f9ca21b1b32c31124c9035f7e1db1ce7d3684e7519305494b9543ee5b975726ca7e06fd83c5457fcd34bb6f66b79842da324113cbad78ee85468a0e61c1a5ea5c4d98c9499f89bbd6172498f249ca7441e30b578c3d8d9f6667e37b4ddcd2c46a325e5b771561788b18be35185b7e464e77d8ae5ebc72c5075e21e37135f7272479c482feece465953604588864f7456d65fa1986e4790540f563a742c1ea946581c2e00dd7fdacd9ee2698e44361b01bd7c49691eed59ef53d95db378f1fc2c42295984e220b371cf45b1ce46fc384b99137c9df66175a30bb454dfd62f68866382ffddab3bc55abc8abf96ad9f18d8992e11b72edb75a368b263e85fb621803f98cab971b57c0eb1a245378acf11452088ad86af2ea8fd05191da294ae026fb7f40ffebb6ea1f8e729f6c6181b65d8074e3872b8810b9c8ce43e4297dec19c9704619507bca7e1dce4db1e9422660ae346ed17ade483fabd20ae999022ebff6c6f3c3b693c8e158e58c01318c0a2fc4b4641db53f4afcf3b9870d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9aae4bfba9920a7665895503a544594492cfa88a1852875b7bc4caa277cb5f653b11dbedc56cac0c37a98ab8063efcc5a4c096167b6a505eb2327012aa027f41d0cbda2e00b094707259cfff4f8d02a8b7bcffa422cc605722cb4c1a0721129d361a47349a253f95619c7636d11e970e633011b0f7691e4a2b9c876a5b9f6c1f26cdfd1ad0e91d83ae12735331494c9be44ab92e806baccd268eb399f74ad30e3ef0d9fdc345eaaf82723a4cb3ebeba233d6b39b321eaa22d881671ea788f310660a2d4f1e6809ba4b352947e3f216f17613303fda555dd45542b886e61715f8e8a5ab69aa937f82d9435a5c63373b253a76016c6825cf6be49783e2c32bd8db4deeff8fc38f844863ba08c061ead041df36d4c387249bc2019c02daba7dde2b53352dbb493e13442adc88b72cb7121ca74228a206c6fd1f91f3feea534388465edf114dc5dc4e34561e96aef9f588fef3360883e0a5692804690a23d0459e726a3b15ce3575d97752b4e32064b521144f27a5909312b20568d575e1a86132ce73fdc7d5d2031bc1375332f7530481963626d92b0ec86cd781b60b9ba7ddcd7cc3e230b6d0df2cb9638b46794f717cc4551f855f51ca9bf6114e15349af5456a144493cdcba817827c1f0838ad3329bb56fc40ba47fe81a4a23a094cf0f199171812f96f0cddccce0ba0173cba3968be58c27ab405d95eb9892ec7144b09991d916c62a5f43e76f0f6666a6962137af6a857d7c431a226641ca2f11c2598e0421c6582bfdc5599dd293fd7df4af7737a423d6d59ef00c38656e198d57ad05309cd29caa9785d37177bc58388fc027eeade1808945a133b21857c6edbc57cf99c46690f3bf9ef57942ae22fdb4699b47d026eb3ba5a428aec5b5a34963691ee44d4fac56bacae07f20c55f67f2ede5c060076e8aafa666eacc4e03bb345a48f08277a7b9f80a13bfa7cc9288bc8d548316b80e242857af28e40bb3b9acd046af46698ee36d9ed4373c43dd1b29cb0a3cedfb67ff180b5e62fe12afe95bde24a2d858e2653a575dba4627f6b288ddb8af8892473258d29e425cfdf5a4290378d18486e7717774b7643b7047d0edb02ce2f54dbd486db081a3ebd1b7ef29d434405cea939dfab0ad34285574bf234cf6696096b125b54042a1fd437fb1171c8bcfaf941536fe98d9bfa950899da3a01a0d5b202621a17b8243bdffcaa711e0bc0fc8fb4662504f70f059e01eea9c77473c424c4e09c0d3d5985867dd842a37627564e0503c1686dbf6759fae9667416641ada430facef2249a31114c5d99f7983ad39161e7c39abcbdf93d44e6cf9f35311d363ec8ff4491fc30d70cb58ca6f04295835dbfc690cd7023e93b4de633b2069e698244db695b7ed01c3aac717064c2c0bab9736559bac7b75b82e0e017ecbe3a927969b93c1b216dc1552eaf672719;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52f222df0c0272d297bb815d42fd000371579dc526d1fc2627cb61171978c7cd5eecba968a1eee58aa223f343a2743d72ae01b25e2671c6902ab3b9e2cd5737ce228eb9bc11abdb91705a9ec87c20eadb65559fd329c9aaf89d42f2706cf8c3cc3f57dd242fabaeedf5b8feea294c19919eaf22d497a56b24f93c74cf589e094a33419fd95104778e18dbb5ef844243496d3106ada43c4dc3681e9cd281ebab1bfae9be872b6dd55523189e1327957cf35eb9b6ecc29bc355316df0b4ac8dc13ee757e727f71301306ccea2dce0989ed4dcce75056e07e9dd44e8d8348d7a27eab612a9b4bce615bc454b32ee8a7d48071c7e9e3fd32b724d3896a3ac405ccc04b3104f349a97a2211e565011eb55fe07605a3fce7ba41b0cdecccdd38fe977f759611d1b8beda7764510e3e02a4c6324584566747ba455d05a258e765739b45ca935084c93fd6f29810bae746f2a916b2dedfd6a0debd36db15c3979125eb0364226aaa4cd41a81b11f042b51d753c6d896436b88b7a10085a0c7d0701a1c5baa761d39810bf1ebe44550891b32bb94eb8f006629ee696eaf9f4113ddac70a041f09713aabc9355c2b2f05b0d84e6303555f61cb77ae023c5381dd3091d024fef2140022e721fd035113010b47d28329c1bc40ea89bf4253af5ed395b1453320578a193b76889a466fa7412b9b4a49b07866e8ba06ed28ee32bb7367f2358fc1820418c0c36a131dac94baff79b45f61339a1afc322e1e6d4b8fe5f4942cd64a98e045a036b4010956d11d236d19b979ec47038ac41bd66ada84a217abe76d8e63b4081c214b31abf5ff5f966de80f010275ab6189379e19906ee5784a766145032211cdd3926f78f7352606030062a240cd70e9ea0f73a33516c6ba9751e3da089114c2917fe932468535d81cd1719bf874e259f9663dd6a8b39c0fab114541cc14f1d1d8bed0cdea6b9acd190043fa4d5a41c337dd7919301f334b6380f31ab5f74ee51324ac03bebfd6cc91099db7a71f4a90ae3b694ffc6d23dccbd7733a63a3a175740c1a4c3c8ce49e1c768d18496d4b8c609093e7af1a90930a1e70c602320e1641f96fef6742a36ca5208ed9c5dee367eca93f79c349a24b8658cf402ecc02f59533af843a951b56372aa018c75b50d8b8f582d40350bd8d458ab1562e14f3b579a771f4b072c35868f493e05c9e0a565b2f57b71b7b759e273d92aadaa945379da27fc104dc176d763b294de623ce1d98b086c01972730453f573cefcc35480925e4a645b12550a09082c83f1eae8cfc712ceb792c281e45f1fa9ffb2bc987db4c01252fe717aff751dd680f271b291450ec594e7dfc14f90516710b583d534a8931f52797b39fff8d5d35f9af869b903dd983fd167e57a8f8dc261cd39327a8c001891d6be2026ff5bdbd5e7e9e6fcd212b573a49697165b3851a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he487603dfd39344bbfad462d9a2d00bc2dae2c443d6f93da024300e4e88249caf3bb8a4b61e97f2e355f217fa75a91ee9b54b9704f7de8918ec1f2a1d5c85ebffd10fec1d4d1650d6c4501fc251da71e56cf0f9d94d2d3b38340f34fbb2f1c107b84daf0e57542476cd1818ea833dd68047a8a85c4a774dc87a562cd401b1e330f6f06e37db73a3a80e53d04fef027289b924400cfdb854e30d673debde86a1d21116d5cea88ab806c42dbcb22840424dea344538a475673ef2906b5616863f5fcb6c2236431f643ea3b1530161ff804ca2a49fe856787b4ad7a234578010fd57c42e1690a0bdbeafb2e91ef81773b6a73ae4694ed8612a39358c0366c3e1c760d133fa7a6182f773ecd48603fde9b0e866f2317f1d745060e1df36a15f96a863b39f2da7a5ee1f9cf91899a6869c3dceef430242ba08e5d179a7c0cc5ed69bf3742bff546bc8b04d5f97c554b1f0eca62faf932757cc8921457ba58611c8f22d6583e4311ae9dc681ad32eaa9113cf6a1528e09f3d283a9fd46affa6fdfb276ba73245c00333538c4361d3d1a81a01e511369e7f7c1705d3467019f040ef56fd2c4069c6cd75b42249cfa935ecd3967c2e216cff4624a814b20e8b801e03a4147f016c919561e71a663528573bdec6cccb99c971a6e4c696ebc938590ffb1cb5c30a83ae4cc2f85bc0961e66da8874f28939e71fd295f4a6ed34fb24fa44a8bba4bec1586e13ca0efabc553994f39a00dd822e85ea25131463333a640dd0ea2ecbaf1424e7f2c122f1d3c08ff90c3f76507751d29579046d9feab2850826aca0bce7c90c8ca85b0f985be40c8689c77d9b504a7cbd62e663a71031be2d7511dc81d409fd496f73c4d6ccefe14271ff274c97c91b657f253900a410cf5fdfdad1c72e3fc46939b5d607322c9b647125c8bb20d2041a657cdc099ec01369bcf4310e3ecb575102e18e3495564a831be80b03a79b54771d5b679053c59c446f2c74996ed07862d4994b05e6437153ab2d4267b1c4b8e875e0c8041524aae72f4a3582a05ee55c1e8ae5e80735320c621dd7f238d63af1fa730ba5980a44c811377f3985f14323b1ddad959f93b2c9b48ee77ad99c95fbd78a1f46293ec683e6d499e2a1f8794fb45418d506816794e5f687647eccd7bbb252c9ef3644771c602eea36f9d0f8c2816cad5440fc4af213b91f03bcb5d601f3ce728d8035692624b2036e22706f1e512eeef7ea54bf6d6857aaae574ac7011e8898ce0f16977a14fd368e9460a7ed28629d565b41dbc8ad50bcf53d493f3680e0b288e65e2811e49c33776c46cd2fb951d128bd7e0822517eec95d890da88952ead378bdd4cbf895ad59b784cdd777db747a344a24b32b52b18737219e20858e9be3e8021d1c2c3df3b3a49511769ebba22c50df61fa261e814cddda15fc3c8b358a9b3c262cb10ac1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h522d18df394c7e5ef5934edc62161d7465835ec43ed573ffc5652675b682eca8df6814433e4e3dd0dfdd613b1b4cd2d4372c9eb59f600e6937a07db5dfc6c6e055550239451ee9c959546c44ca8268ec4759e9fcfa7c11e00ca46b1573bb5a9487e0c80fba0cec28ed33df2987ac563357c74cf85871999cab9f902a3efcba77097f686b4126a352863e0f5bb2b16d6a1504013a30de9b4a86b07f23509a04a4243a1ecd03b10c16d315b0f70fe8a63c957930d329d4b46636dc1fe893fc3a805dc6941cdf5ff15829ea472d9842c0e9a891e319decfccc237b5df80a58846d3b78e9945b9be103ae91418a2b65b307c2704731b6ffb7389d86cca8766784754b4208c12a7e272dfdfe34983e56dd9f6dee446145ed8ce9a0549a10c24089533ce05f5059673fbb6e8e8eecfaef612d3f023a30458da1e045dfd6a218ee7f378d500aba07bfda0afd7de2758db43c1401a6c4075ddc4b0f8b56a27169e90a75565671456265f2474130a43c2f9fd52f7cbd5bc0ace3034d307b8a46a8b993e56bee9e48e1d7c9e45c3a688ed08484529626cc54a62cdd5314b5e8a843670829026a7e01cc682a5b523009e0211cbb31b7d1acfa0a0eaeb0cdfcdc239af841dff8b68203f52d63b1ba53e827341f4ce2d1294515f4cc91349540372a3d24e5812eb6f2928280de792f0f837524179f0ac759debb720eb3a1098def1a91b12878094aad9b502ed11009f0817301b4615fe8be11f5ceab4da3556f07633c096902a05896d10d79a7f3ba335a4ffaaffb3ef3766ae35d07e7dc39fb536b1e260cd0d40a4c2fbe476f7e68b188b8de0dcdf4daefcc5bf8ea1111c5ad80b2ae773bfe3605ae71afa6727b6bed32f4a0b32c1d116d254d2d518478eb6d65301c3c06a4b14645d903f0e76447874346e1362d4a6a0289a59aade0889f3d0a0ca19340a4a43139899a0504b8965e4e4c9b8661099cf91bb6f92ef3ed96adb94e7207f4b87a9ece698dd6ffc6ab37a0f3145c67ebc5fa8ee019109c12ebd46884f74a0477e033ebfab3cad44f66aaf5c19f2e6bf492ceb78cf8b0b4a4a2b55fcea6dbbeaede81719e2b4afe9533a284b0f254488ab481f1bcff02d4d56a81c1356dcb5a301170232921acc0a6553bf497a613a78873f40810b2356172a896ef25974e9d9ba9b78c941ff3b3e36ce7ee49c821606287e68c82e6f16f7df79d78d90369b73b09de7fa924e5771a97b4d40adbabbec55f3a0bd98bbe919ecfe636d33f2a0dff5a93ec8e98acd221ebf826356330f3b29f9608812b31ddf7bb7ece56fd3a4bd22fbc55c58af42d72a43376041decfdbeb5e35b50c5f223e3f20664871416a19d26e21b8a6f325346f91406f3d5ffd78994e1451f51658911d5c2cdacc0defa74fc788101a926021e5e08801e11380cc00af76f08e6e25dd76d8fd7abb4d92da88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4eba68f71f1bb0aa10230d31cf4948d49e9194e7dce4cea274807a603985c84aa72060c29d482dd72e670c2a0567358f358efe827f2947952abfa774e2bd63da90b6df4a85f1c98b23481851388dcb78dc7472c9544a77155f7fec36f32ab1bef62740154805b2a25a228c08476a883fce4e06b4086d82b683e3868422de147139c105f088ed25e5e0627a83ffd0e6b69b86efd4e28572e3a9e2612ffce785ff4e3bbd74f2cff28609e4f1d5df552b051df30b02bbdce48acc3e5eb5975d1e5025a2aabfa04c02a49917708d7062017cea63d7da5faa971feb79f91761c4519845dc918b3b4c7b2ec3e91ab3744c32416109ef1814acc4d06747bce0079cfbf81e9dd24751239c9b6d4bf2f3bf4bad72637edce8bcb8fcbfa9881081d00ed67bfecf0ee61104a6b3284007aa16c000c877c16b8ff1b1b32a96c42972a50131f82bccb2743d02bc9017f1d9b445c71712bb8bf78f7443dadfea207d0b6f3e5f20b09f95bb3e8b1dcc1e6932efa1e5dc8acb678040c930d989e34c19dfd5d1b21332ae4e84a5a8f1a7349d00273dcc01ee515ac02402610dc01cd0bbcf3f3ad43608d2676b2e1255d728e92981cbe1b40b81a872ef01f7b5d88cbc9d370ff42225e33d9a122fa61c7430c7d251fc5196800b24ee9ddd2ec8549ee6000ca22514bc29d65b1b1d13c676bfd39ffb14cf428511bb7e9dd74e5a1c79156f73db6d2f020701e69008ce99887162b2229efc3b9385ff230d7a21133dfc657ae67d8647874bd89ca38f19240848adf7ad6f37cdba99858ad8efa643d22605bc5814dd63eff328d40fe8644d8362ce0687a42a497f18cb62aefc9074662fb051ee0d4bb6a1e1604c7bbb20cf0f9fa98745951214e9c3611ec4a0ca0be690ed8e4fdc952407da4dcab967dc4c4b5c33fc839785ec5f75655693593e67a6a28010c0b4e47d8f9e9e52aa24094502dbc69d76bcfac3f72e828a400b2e7879d9e5ff4c71a3cfca1d1e8a06f8c380b0dd619b982dae549035d2dbcb6ed76158e63da0bcaa85a819c23cb6564ced270ddd9d6d539fe05b29a7059145099a35aa06a8087b903f4b13d101e90a91881f26bc9477542a8c10cdba0757eb1e087c9f0972034caadb93aaa3df6cc1ca77e339db6fc81d16966cb2f5bfa994b3b46f3caea306d3913bed505632fc6e5b13d36af9ea3d0e96fa352aa1c2fd13a5e1de7408cacfc336c170b7e1a2d77746e7d6d39b7116d66ec5960aa97beb622d7f584ed18310a660e12a33f034dbb55b7d14ebed23cd7dc2a5b2a244bd2c268fac345d7c43a96d269611f81b4b329edc4c2b7ba4346c129e10d273ddb9c6fad9f207cfe3a30c4e770189e0ff5e3b3e18476733a5e8682ea59496de7f53f96cc66030b906906a39c3f9647e31259ffee60da23da17e87b0b3eed062e09b3dcb880f1c0d286fec0ed3a3e4a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf725f99588ca9978e6771a891fbb2a9284438600c85494d04b18fb94e3241c3c0f4a7ab6bbd2296c48e7a2d6ea1307160231515f390f821f3c5eafcfdc5a4590b50d6e9fc3777f78d585b0f95736a5e0789dfa0f8c32adbb533ba73914c7abce19634143223065bd87a54b32b04373e2b7d2a159c7be8a64b7f282893efd81f37ffaff75060b3efd2fa661fced54f45e8499baeeff542ed82ceaae2dd34908fe466124bbf7aa37096adadcf0dece047726e317fe5c254c447b84dcb331e19a4fda9edd751044b307878e2a99bb8fe0f7217f8d945fafbb64fd05d347a24d1437d21af033e3d3a183a48dbe395f429b1ac6126bd28c39c323797e66720a7d0529d2bea12ac46d8df7aec1fa93b09ae87deb310e9d5955b55d176baa07e673922b73be4f5a8f8678bcc2a0c5cc8f6d5a2e2b4d51993845667a6463922bf151e6342c3655c241bd523daf6f358a527340f11bfb5067b34aee68224c323118663ac4e220ffd14edcee884d7a7f31fdb8042c13694bef8b2cffd82f6173f2ff00044b7fdeee701d7f98e0dc535a95f75e8c5c72b579166a451d230110aa5a3b15333ad6f51413e3702fe54b7cd67411fa3d172daafda21fb30baa6e28445004b9250c8416fb5a5ac49386b652784324f4e9f8fe6ad3686221b06d86ac2336ac59c918a37331f9f3523af2fcf18b800e1c2a795caf662a4b6d6c0c375f60b82078fe5e8d4ab69b0725aca4e3bd1949543c4f451633586e638af0c31ec9c9b3e7ddfaff44e47d4391acd72faeddf39e68a61c1fd9686f1acada576b1f562bd19563e6e2cfa7c4197ab79df7fdc7fba3fbabba718160418e728239d342244172d1bcabe5d5249add08ffeb2cbd974249b9b761260512f0b7919a145ef4c64007c001e0784299aae33c624bac35bdd73a78660f641051461452ca119391eb662ece5cdd36e173294f5bc17fb1f8577efb4da7d4ef14a299cac9833d2dad8fdd9d7709f0fdd03033b5979737192218757587fe40592590eb7c7fbb4219b6c87bfb748ef8cea7e862e171c81b21fcddeae5e2e8e6e6ba10dfd1c5339893b2ab1e19c2714643c939c70ee5865e5f745e6a3233009a9fb2d22c2273057bb99d3bd4618323d6bd3fa12db109a4ba11d3e6b0264c4bc77167647676ebebc332faf5bb4ff783a05c4f8db6ce230b0b8bb87476a5fb1e8e869741a8eea2203b2ad19ce40a5cd50f5c7449e3f9d6bf6ce88e538bf69ea8723e1e3c19555ff49f7443ff6fc6733862bdd8b13592d12726beb7a6bfacfc7c696bfee049d8850b5376b046bdf91b5248b80e30e7bd26e3b662b589adbf24f016d593543ba022f60f92ad27a12b025086375147cd9ae0288bb8a2981b4ef11369103481684b0f1176cef0455b45e18fb054d4593fb4d77eeb6c68b576b1c26c650c90d86c23b98aa66a0573484c6028b9ca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7aa77807a6f7bc459474247d2767abe8f3268bdf41d560f0836a83bd0a50a39d6781644c719f5ac28e209d0b0972c27a4a4c7b1b31c6ed7f2a24ecef4cacb8cfddbda30a555ae86431603cb1fb5b1284938e765a2f1eba239f704eca0e8a9f513c365bd21a47a2717922e7ee94cc4d225525bb42c281c64521cccf9de7918dfb8e6a105378bdbdff1a0926fe084414bf834e96cc86c4075eb5458c066a128a52b16a3cddd406f05b9ac72412c1ffaef2059f809c8ec788a0c62523c33cc0d29be55dd825cd674b4e379f28deee6e43b9d4f0c115ac92e49533eec2bf9b7f4bc2498a180dde96b92e7ecd96c54eef26bfc873ee20bfddb5b837158b6a914df69522d77379db16a55da61fe657db691137e18eb77d82742f9887dfb2a084019835880a40724dae80f61d2a2119653f152eba20ae0831a7ef0dc450f0ee59dd5c23cc6d87cebb62652d6e68b99677c2da13ee554e78a609055e728019eb7195b46e9186ebb517e818f16dd8d8ae209c92d8a9c4d38e89963e79633adc00e67e53ce5c2fb38003152ee32dcc4b64518ebb1ae7bcc82c5a9434e1ba765062f38775cd05fe9bd4b0966f6861f9493ef27b46ba1777e0929936b1e13e12db56c82a088f1e5cd40e50d436f270d3f368d9cb3e5da6604a694ac52d7fbd95dcb08190239f014edf2e1424d83589b554366d9f981b9a4d488d21c8a1ffd68be31e6331cff0e0d1d4e560e9cf2b491db5ec23d5c03a5874915b3f6392c481eec781455dd932da549aee8212bc2a587e6a97f064b4446c71e499f1cd16660277a0ced3206a4981013e59f96e08d4c9032692781d841c230a2035623c39d04274f2a225eaab2d033ff45f425ce918cb0eba865c80226dae1cf6b9fd625e7b67bc3392f2d3d049993b75911b830d48fd64b1c2a94a993257b428b28a6ff32d9ece88b4b4a441bfb30bef48360c9e4cdbbc0d2b15e23a8e53d5b1e7d8c9a825978d3e06da8de301ae2d891cd6a9d32f3c98c0fe45be7ae0039eba808f39c824332f627e7509cae113f793eeb2756cd732224de1b250a21bb8369910300f14f92aeee54f26a590c7b2fe478f13942b5095717fd99fda68f505bd622f9fbe7862d6e0a20aa4e6933f7ca55da38e1cc2603f02f4cadc895b090a90616c3a23ce3be55a57fbfa31b0b39666ced214fc4df4bea84b6f1eba2413556b5ecea0c2c271eb86a8bb90f570ac799f7c15fc015b955fbdc9993d6354820e04ae4d111101c307719111bc5078b78ab19abce91185f8cfe0da0769423a2591183ffb71b279e042fc76a09058dd8e550492f4acc2ecd427621eb2f6f15a5fe9def701112d09928fdf47aff031f99df1de24bed7a61dd43b10d1d085e1d33ad68d3d8ab7f0c5b98eefa84176274e2d0749fb8b43057ec1292ede484e9e59abe697b7330b02ee959680ea9253479df4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h55710e36f59aef6169b16121856fc13ee7739b8e8cede1ea6b6093ea290705e527a28cec0b5bddd7466f1a3757b0a4b63a9feac5666633a874dfa5598e8cc485da252c06f11449828b1692b032d351fbef5c8c86e666272f9899a0eca3b56d0b2a57c5b132ab16ff5c277b534e2950765a0697656798bb4c4a1b1136efcfd2ab06102c6ec2f221c9bad34741c6ea27274522684c7933c8e7dfcbfc6a2fb5439c44bc6019251c12e8168ed504869623130f4481c90ce5fdb82b54373170dd446c086c5d263ef94bfee57f16ca6ec4f3a345a81507afaa85f0b90736588e71198cea0e3308b344b6d446cbd32f945009455a8b0e20fa4abda6970b208ba4ffb0d84c3b2e327ec5509e79e213c9a84c76eaccf2c4061b1e096bce373ad016498ec1b307593377d99192128b1c3f734ec17e9861acf2fcbd55ddbca32cb81d015032b1ea9585632164193f41b950d6a0e7c299474d8434ec5da188cb0e38b32ddd64ed4ad470ff0e9171b030de714ee29399403dc8949a8f07eeec9b74a674b4d4bb34c3c34953d8c6e9205a3a72e0f16c9b56a5bd06f1064c329566f3f758eb36ed73397b762b0c1c52a0c9919f1c99715ab37c853fe0e4138faa81b57767f6a28348275ef9f9e5b9ad5eecc27d104f684c14ebac71f2a37f53f19584d8bbe7f32b8b3b404859e58c93b79f3d69362d22d310d4f2525d02e0c37d5ee75b3de84403a363077057a0105cdca092a807c34f580d6b28cf75172b91a26bfdcbddd12aead39076c756df4f085381413492e6ca39b855eec8e06f894d9f29c20acafc86d50c063e544e531098e789f84b07385a03305f2a7ff365809352b602287377500e9a6d88062f9dfb3b8adb080c8f9944c27a7cefbb5305156a73d7552dc7835ae797d616a082cfc8a1806644608490f7ca07bbe61fcc77d13af2bfc5b94e2c160f2b248ce4da26760b4963771ca21735a0be6ad97e0068c020953d5d23ca1ecd5e07ed7b7496514a25e6d1a4c0ad4dd8ce644a4568396db9ff1cd1bfcc06acaf40510fd1133d32978bfd75755e447169c6054feea7a3ca2d53f7884a72666e15337471999b0c4d64fd0ef4eaa52929901c5eb93c7f856ec1bab64a538e04ce7542881fe87c3eec149e53f2918d75fc61ef36ee6ce43da92c81ff6278724c22c4b2f81cf053de36c0e1cb73afd8ce9320609e04e07a8a2913fee6fe1b13eeb9c92579f255aa5ca3ab80b3864a362fe3f8ff663d0504d763f96ce9196dd7fc1f1157c619c39db822eb9fee1e57d0b8f6723de493a95eb066d273303aae446cbb050a213dbc16569e711b2c6de8f4ba1a8234ced5f025c2e218b2120d7119924de2aaf17719ca771ff33da6a313e0e45c1fe84584c4ad15ebb8d14528659e5bd660524e150c432df0e1fd7827092cba5b6252250c4c87f06ac2c5779e5619ab4a0604;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfc33863445e3fdb8001f22b80200d4c5f7cf13dfa63f0a4391076ccfef619710e61e4734beef5a687339613cdf2b26ba403653ae3ce3891438b31fb3d522bfef4fa1b96a6fe4c7945e988a31c9e97f0ead1883abc496d0f8a9b0c24bd5cbca255fcd241c6e8a00db622f652a62ca5696793c8b3b19077f3d7f58c653e1d2dd1aa1852ff7999e98f74c01ed85c00a19e49dc4fa95b542a2eca40236ed8d2822955c80d954b24616fe98679fc57205c39a2e6836cc54c8d2cab6fef76b30b4478af7b6d1cf21cf5c8a98f46f3e6ddd8537dcc33e1626eca7074f9c209331e47660ce537007c0273940a46c1990ac894f4e2e9803eb487120cedaf53767bfde92f6dfda3eec9f86882af6b2d725cc88435e310508829276a4da06ecd7eca1f52aed28a3d8a8c3a3bbc5829e6aee98f9e414c7f3a24caef9c6df548cf5a311802c1ac5f0725bc7974682b5ab0207c958d7da442dc872405134456159336f3ad9fd22cded75cbef9a4934fa67b9e0b5fd829080ce77a1c6a06915c22e0973b00678af1bf901a24d9e87adc08bcc9b109828895371b3a3e577a2f3059a3185b8bb934800a52c48f7579d21b1e85b4daa5f0b923a2cbe0a163a8261d95d2e0d1ce36dcd9485d8076511bd7e0bc1f7d49c4b8e5ca7a12ab0d92bf876fdc66febb60ff5821fe167f6a58034810e194b356e35e514c17fa52d288d67c26daf7c771f71e4393cee9e642b198f6f8eb52f0c87f3788d6fd4a300a7f51196d9a02c08b52577f4c9bc11ef68f917f05fcb9c8781590aee93fd8e4a96570034830917272531029005d2e913d3f372c4227e75190d8b5e74c7849a8d072b27e58e654dd96eda31d539d418d34e517546213c6dd8ee67efe34705e26eac68e6302071b937cc0c754934b8556862a2c38ddd05aff4d266d046e87808cbb198bb5eb8033b67d74c33a8050d649600aba3d539ea353b004068d6d191537e41ba34839dbdb6297a9e77224f9e4ac6cabd3c0b344837bd6f90c5c1ee061ede0b6d665c9d57da03aa27193cb51a878ca629f5cb9a5a7e6b8873b4f1f1b33d4dafe8edc7993b759e8169c0ae475e3f399080905fa25b35b5093c0df7e1fca8c3c39bf676a528dfc73762020a4a7aa07d9f2553a3a350f190193b201696b8762ce07bf2b721b5c9f96259d918e1ad4cdf18d00ebd843a726e14a2f575c8018d1584e99abfbce25b08b343482b92ce77a85cb96f659b02060a74c19dac6a0564cd0e5354b73bdfb78b6db1773ba0616b76c75bf9125053c73511508f5201fc3c1676efd0d904e9019149bf778af24a075337bfc7ea0d8b6a4b1e8e31e88f2bb143eee9afbaea930092de5ea5492a85cd5d9afe87c49bfea1aa64b32dc2cccdf07a1bcba68ba2f0fbf57124eeed6527e82f0605663c95b33400c684ada08f83250a1b5db5db68fdff954dafc848;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc0cbba0358460769ed553561bf3b3708669c29356e55fe14726d423d62edf8f91932554ced2c7fdc09063184dba0d5178ebb6f4c838c8f4bd892e893e56cbf5fa38ba79ebe7276726e3f1bf2eb91170c91e60035f29c1988ab64f996837ddc8de87c3febd206ea7fb657adce5ce301d690c198adacbfc478b1e3cdd2afb21da694f33bba11d1f4b1c946b6dd41c4e8f94406aba5b7d87515ebbdf8cba29d13a31fac2400d106760d4105c9c8fb2cbfbbcf9a29bcc6cb843a8d4cd52f9092b83d91cabcf2d8d19bdd6730a8d9b7b800712ce60711e67a6993036f8ef57be93c0f1d3dc6b2e25602691e3e0cba0dec22efe0cd8f3d6abb6ea0928e8ed4469765448f3a9128e71ce8c29453d89e68f85ab2824b599c9c98181fbb0adbc70e98aaf2c72ba60a1286fba87959c374ac79a8c8fa4ab0e256e61c31f6556f6851e56131e7c30b0022468d073298d9724dbf19fa1ff90119d3a3b331f855f0bbef1e7cff485a23e82fbeb78ae7e493d4420757fccfd77104aeb1eaecf8c7fe4cf2bbf93f416dde4ea2874b19d079512c820bf0f446eeb20c3038756c4aab8183c9db62926d9c204fab81b8e13ff926349f7071be05613c3b8d96dd832e5b38029a2c492577382ca44a422b5858446cf9d85e51fca98e643928439668301785f49440884fbef69fb92e13bd77886979e93614c3dc0ce901639e7311ecac06f61116c4f79c5784dc7f4cc971c4b8b4a623b437eba8704fcf45d0b7b6d7beb8d6e36f71704463ae9ea2a9205bef2d4b989d48dcbdd5d7d7100f3c24f21450724b223d4e6beb4f2bd11dca9884264fa89a89909d444281f69df882841b44617d347529162d7d504500380b6041219d85dc970ac6c5b3ea5a449187606a53c123e1eb43d93b7094c4a7a3598c639ed45f0bbeedc8e46a0a97acfc5af013c4e9766b4cb94cdf5bb03b54bd40109e1afb3c75393bda5da25f04065e70e386c36679f1f1bacdd6352169111b224351a567a03a8b95e02d5e61dece309c327f1c865537a06149bddd5ac57a256ef097c3e5b9ed771f6f49186d7e7e1817459dd81147b3863a1d3819a9cbc7d73c42ea34a94b46e7b0eb88e0f21ea81c09bed9eae56db1156cd697415562d9ec43f48471efd0e20ccec7b40d0e7d122978d1f4d860fc472b271cf395ef8d831bfefa4204bab280d5d5aab901e6e708b51b697a71bc7cbca0233724499168c52f387989b27d196fde4a75316c3167b18674cd4c1531f5d7532a614efcbb74299dbaf9b46cc271a0b8b617bd832ba6833cf2939aaa339d767bdd70d9537d139c1e0ea3d8299a391360598f7a34032b489002a3ff2d67969ed49bc6e9eab969fc225801e6f202a8c5deed608fdd7430b26ce90947c4cf132343f16a92825d73692a398cd89df69080cc904b505a4d430dd7d565c055b99a9c01745183a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb849ee02b69bd9098497a4fe9068436706aa82e26cc804f3d790c253094760a23ac268201486cd357ddf023b61c78b5a3eae4eca165276806fab635317a92164354612c5cdaf09f82394168539186431e08c7b0dfab0a9d3fe4e588ab75828b7f2fbada7944b3b0ea2140276f0450052c30cefc05de4d579a152aaea3c502908d9754f5ec4461711eda09ef2f49d82eadcf8fd40f41fdb3887919539b49918c8f688faa2230b6eedd43dc2d12081ccc622b3d97fb2a1fd43e8317a055c45abb167befe0f163d60009f2af2ed4cda1972cdda13f6eb2d5520217ddcf00057306c498ebb07893a7426be63a13a15b5a3110d9981f2f0ca1bfde640eb7b139221fb389afdb9de88e69e8583bebeb05ff71d65b121319003ec114a6adb053c017ca6629b4ccaed26205d905b159f87b111376fe94edad333c105f09e0c9a69762a8f2e5ccd2aa0271e68bcdfb45c999598d54429525de81ef20ccf051369b4daced8149ed04d9f787abfc07f9266dd2f23e27fe7439a9a234ad817570d9599340b74ec49f838c2823b495480ee4934c3388ad46eb632b5409edaaea2eb069c94747607b677a81074a221a6051a5c7aecdd8445d12f080437e7117137a9d38ce094b11dc2e87110dad56398addcce4fea8ed24f651538f72a6755ef52c675b4a4d81c0482aef4c587569208c3d4cca2937545fa6cd5443173496fcde0dc4913c5685611069599f4b404a8b24acea36c1464b16ee418bbfe6ab34617a8c9c62128a786120bb858d4f945c5d4313cbe7e584d0eed5ded39d10c2487f013f65b127b872048d67867b2243ecdda550724dd559d6a5e37dba91da4b91fa41c059c4fad2b33aa0def666925e1bf058986fc574e108ead60109800d0c9790b76093a0fd8b5b83f5feec8c778e8245df3092553720ffc443a1d826f3ff268053a5945a6cba3af115b0fe6080a884e586c6e320bb9a0d1e76a739a269d1ce32a19eb88fa66a60b5e13895d151651d78f49b3d5af0bee59f855213d7b4f42a383c91f905e9e392d11f33d314e6f2b0efe67c2613c9911820cc37de031b6d65507ffffca55e0ebc83024798b7ca0dfcc75f83e045e46abb3f2c0c6794b88809f2294e11eaad47b8ba29eae421d2cfb0859cf43569f88711c893bfa61334c00b185a0f5e5211efa447ef709b8f1a499a6e2d81a9c85f092e59d76716565df6e949399e83fdda99e2b60535eac8bad1dcbe56d02f700833d613d09a49cb977b415f306c400cbd9eb0ee82ef3663c2af06969cf0be1ffaf399a61d4d868c443aa5eef24198b1c51805ef0e0753c7cf33ee8fe5802b51bb870c8912ef407ecaa19d86a021d84c14fc3de8d39c27e0e5a7baab6467c617d14b570b612bddca7b7aac54324d6e9d6c178c2a1dcf690e38a6a0da542943e35e40e25b7bd58b1d05f9d098fcd72e8544f7e03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h407a91b5e4cca6e6b550381d7b4a0ddfac5dfa0bd1c8f8624ab80f6f95a880d9b38b4121af9d5dab7e06795c7f07fa9c01ce7e52a036c637cd154e0cec2fcadbb8e457f9811abac93c0bd68888b34e39995a1a5605671d42321059de445311b4c0a28995ebef81ace06bd0100339229d94ae7af396a6c73fc2e20a903d8415b3e3aaa6ff1a8e03c142a98dbe8780ca8a505b4da8c3e16e7a1d1a3dedfafee929b229a03dc83b3fb046a90f57ee68eada6db0cb20fb2c9a3e6f42f20c4bd6e3ec945e5e72fd59f530548c7707f386ce57f6b53d0a96d5b7c02629b31f56b6e8dd08f7a33b617268d74d0d218d7298bb767daa0a122fa9758d909af4c69fa94ce51f1f73e03955a926634ada262726c65f8ba882a49b8eaf356f33d15f9a051a4db52527d6b0b64e9183c1b76dff73a834fda9d1d54722b66df6f36dfd8743073cfd25d3631b2357eeb43e6609065bd1ef2b7a30aa8b4da9b0142f4a8222f1105964b86e47fc604cc3e35de179b563948445aba8c720e3e8927f644298f8cb0a55957fa3bea236990d5ede930a76d335d973665252e5e621a340b43ab4da4b2149879da6fbc755d05862c1fad23daaf7598dbbb905e241414710ddda7b595bab189f7f88ee641c03a0259724497233526ea7b825e63b5cf962887c3ef68ebbba2cb4d75dcb8fceaf14a7a3f6050b46fbaccd0343c999ce3d74544955d3615e765a84d5b1975823d92384fc74125e5f84687a79cf8063f574148598d96877d96133bfe2c3668b8c685fc765b980ad516ff3df2301e02d156f31eae8aad6f19063b262b98c84af410342b20be9fa3e8a2d4f6e6aed24e33b2ed39f2c7570e7e87af200fca13bad701f6df49d7f89caa686ae501849cd74fb496dd4adeac08b1e30f40b5fc9772283ee05934525ca23aae5b7c83d21aeb0cb1479bcc8cde2b802bd25dc1253ee7df28757e02dd69836feff9d24aaed116f94d559d79884c4bf5b8271eb832135501885ef7510f5f1b2de7d528e062734a0267d6e2b27328dc438b222c41be87825999b15ac462e7fb5d3cd27d7fb927262767feab989a231235626f7cf251005e416a8b5c183c5adde693aaf55630712e977d521463d0de81c9a7378ba07f37f6b67a8b324f3ad143d630575a61893f81a4ac3fa01b8d288cf7c69f5dac481f04d3bab1e056aff5076940724b2a6442313b797a2df867f6c2158c59ed8df51fc219be6b030d16dfd6d9e71b66454a327dce1b51f9885e8f60256f99044b096c9ea63b7a404a242a2c672f6c45d54744a552d5e55a79e7adf15516de5565709b8a8f08981662e5adcf90c81bcb58716dcfcc6afca45427846800b999a9974395ec9311c69b34f686f9fc60c40593873003b40870cc43e5c556d5babad22c18465eb9285ace9165387cabaa3a780909695936ac85506c985cc6c4735da;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc778e98d47d1d8ec5384f392b548c3780864dbff13e725a8bfc4630a9b7f9413c6d88282bda87864537ddf043d85c019ed490c9789c56e783a565a14fae49f631f2f9bba6d27900e620bc0455ce80a7678eff4bcb2b02fa9b607e62652c212927aee0949de1ec5bf5a281724bb86ca3c73cda44ab817fa23bbe276bdaba06ae53a1c3c65becf7e1890ef84935f170ff95c28e99f435241f156484a96e4abeefc8d67a79532a61580c766d9ca5b8e922d5334ab4d8eb1ebe9263e5c9b0a2038fb4500f5679133e30e7c417c26dacf9be9bfba5c8f1b75b8770ee2b524499027a13f9695a3d61a2cca54a4fa8285c76626bce61242205396ff146858a0ae8263d6f4700a01f2d9c11e2acd9043dfc09e71e9c56a9065aaf92ed06561cd5c5e3a94e66369ef31ae01889cfdd29bc144d6f10bf92c60587aba46b6daf07a638f9a03a1b6c5f8679762589c1ca8f82597524fe7913458d81901b1e7048702da8854d87ce7df582e6f626fab4bbe3a92eb6c0ac850916bd5e70a664e532c3d4001df9bc923398bfefbeae34c06d7bff779286b5bd4212e0b5cb778e0674c95cc7731a9c0b0ba8b2f3e67da92eb97c1d9f4a6bd0c231cd4c3c6915b6d9039746e05bfbd45dd7f1227b2337339f0f059fdc040c6fea043a1972eac68a9795b42b0f432f69554b53d403451c419f0206594e0fffa20c376765b66f55fd1f03f4ffd1c9e00f26891a8fa126c1bd93b47368cc169284fcd6ffb0d041cf65f04efbc1ffbd4543967a0a18ff9bc632e4e48ff7a36cad4b302f4e72199bd4ec95d59f81d91396c5f691f9ce06fa4784e11dcd901c98a6bcce31f211a3bc38cc310e3602c80fda32089e64766c6c339e635b73d69e2f5f7853f8275107b78fb878c8248e740f26a0d87ad9c846d2c9a0efa7d6c90f6019031ab4caf9756d4b4b4e584b6c0cbabea0f9a0ba3844ecd413942b767d8adf6a2cfdeb1ed51356bcb4bac72388776d8da30edfefa6d89b58cd44479361d31dc7c6e1de86b8c9cd46ac615e4ec0a39c7d57cca449ecb2a17b33c8de94cc51f4efffe83c420a2758417b887bedbc61d931656fdcf5a48f559aa9fe2c50c363bd26c94377f1d2d115c0b226380b4bb3fd0540ca51d2680ae948a4d93ca2c01e3a92ddd9d8f5b13c4ada0941001ea92c54a09a11d77af56399f58fcdeb2fa5b05cba4d35eca9a327e943d341b8195b7e5004a86383d392c8696f1faf1896df3fa1bf19884277a18b261f25bc3d6c23be3d5cc9b42b1df7235e42eefca7535c72700b10284379fcbca5aa6bed6af0e529e1c9b54383e804d37c047303e6d8ed8fc66d876b45c9721fa6fe4710356c7e66d51ed4c183cf062c5988753d50d2b9d8c0218e7acd7c527b812265fdaea6b26146c5796cf65608b7aa80ff21c42e35826afcffa3e6479b4f783b1402f72503524bdae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9087f9e0a4e7e8233ce31415f58209091fa01421e245c544f67172ce5f2d530e59d642db0e6554caac6f19c0c6e4e77b077487e6ef547b34789b98257a37481dac9d35dda6cb3ed2cfa8c37c2e0233c89b8a605507297cfe8693908eed3b65aa087aef3a67c97a3767753f04f11ecd5d388d133a2c526d645bd9763121800dcc4a9e649a84cc235da848bf9dd5426dd4d0c76356fac86b985a534e2dd52dc17f3731a55de3023d3e5df9e83482f3148af10d3a2ade2ea64418160a70d94e2f539b992b0f2be6450c7f2d8541fd5dbc814116d882ca6a09307cd8955d83d079b923e6c1b205caabdd1cd9535f1b2b46f6d6b4bc66d92167429056261894676b2fdd5d845a8de6eea95d415d2ec0b276579b203cf5f704cffd5703ccebfff3f72b51a6823e2a3bd79de166030a5384ba1b09995745ccc07744f0358601eb2e98848fbcbf919cf2fcf8fb781860ed3b9209e3c2224f92d57af04cbad06a442a769b4958bcadf612ba962386ff003bbf790a7e7e2a6414283faa810644dbf67b8df2e2b26e6f82318e9ee639aa70aa1602e0b46c888270316c937e297f678f441f2a05699c7d7d81ac079699068555a9c697ae7d832760f5c3111de1820fd0d529f4c574502d0491794325d72f2c55cad7d4ef5da4445e3c383f8431932a138012b35650a084b54ac39d380c19f142b30a9839f7ad54fdf2db8cf9bab29040d040fdf15902ea338b8c47d1f4b0b7d92eb75ce237bb8ce40041fbb61dd9e915d3857af06b3251271645f1c2d05ac9c362dbf73f0392277886006f5929a157176ae288e28d975d6e3bbc954473eafc42a902b91be8eac519b0c9dcadc20e2e629dc4c7014365358fdd1231a4b842e58562e758f4925ffc5914b4d0a535451d89a0d22e23cd86c61bc9e0e9aaf4133a8130cbd2ea3d353d695ae3bbd40d6a496b8196e4220e3aeb39add8ea9581090400714eb697eec424bab352861f54861cb313b38a54b2c81c8373b8e3a2a85a67821a29fe8dcab504818ee9c28d3edb5868c515047ed52915f72528fc0c323c67ffc2cb8ea51fae5f37af557f102b2d8dffc98f05ca6ae1236d69755bc9b5d16566c2b754fe844c005f51dcee72747eb69406296320b7f62006005d049a4919234b0fde58ac6a236f7da704061cce81d58e82e94d9cd363f32c4eac128c6b7ab3250000854741ffa1e06779d2f17437f29dec04d5357cc517bd3146c4fa29ae623da99916aa948310d0ba4417cda8204daff017189ef72f78077b910525b2d1e5974841e6a243bb485c8dddca91c049f2ebfb74919e88b452f66e97ab500126037df73981de35dbe316b55c463b24bc9a1b98ce7272a1923834a8063f5a707f751644101ed569500b74a1533b280feb26eac5f0a6b688e62b6836c46ad4a5d58ed5874e2b2a0d272970f3bf4cc1130cb0ab14c55e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7a042d3cf454e0483478063c2018f91fe2fd702f8607d27a67f27db0d63be60e5bcd39982a3631cf6d1b969457c5b78c73c4dfa00c74c36fd8ece274d763546b3d25a523e71251ac64d4e5d2c4f046c7ec6e16eb5dfed76c9ddf8b2b60412bfda9ad7f2d8303ace5f6416f6fd29f7a254771a432dbbd5c542dfa7a3226df5607b7040c2f1f129e549a1d4640fa7e2eabf9570d0c2198ca66bd76a8b7b5f0cb09c89bd91960a7e7f7026a19b7214807c886d495e06ed3f2db019968dad196b78546771f3be799f18fa02f6ced39903000bc11ff561bfd43092388e22377eb072f10c057e0efbb3ac93de0f693bfe839b853733c0849e081011f6443c54dc33eb1beceabccddf952d2b90eae818fbfabc7f68ab34e3e67636f3ad45f74398107889f1ebe9cb909b2f9784e940518f659278fe81e50f36836c70e6d4f79dea3f01b3cfed2eee5c646307919f50f7c50cf5372487957d622bd8fa6581b58b6c65451a89aa6bafe10da10a375f5513769224bb10ecb702e52c70eec5b626fd4bdba3ac9f74beec235b45c8bfec2af611df2a574ace902cd6550886bf141c0406bbd0a0571fbb14492a85ffdf19c292e8f3467860bea94eafcb2bbe4b3e58d77c757d9a7a22ac3b058802e2001e0ae9a8e42d0e3662d0bf2169f0b73096b0f7094b163bbf9546903d4f3e9a1429a6b8c03520500568c11740e83d00f5c49453e1a2bbbada635be92f2c4d3db849c4189db046762b8897d5e4b3e9238c4cdb26ed6a3cb7399bd39d285ebc3b56a9702112ab7054ee2aa3decf251dd1ce8529d6a3a4824f0e5059353b29bc58d5f141deb614cb8d5e24c6a4e731e6d779bd792fd7e8044de9b1e2d1fa2b93bae24d2b195da8192ae164d768de64cfe20938a70ab2407e404771937355f3a59ae1aa01c5c48752f388992499a49a4f70ce98ccba810158bb6891e5dfebe6c1f9e07fc01b8c4520a032831ce692bcfc4a6354626f84eb1d05ecaf669674545b889abcd2d1d2814748b3cb764b50f299b6ba7b7387976c89b86af0ef172bc484558122dcefe939f1519fdb9b88dc8c9f28552616f16346f684241a07982baa14e64222740dcafdfb524405c3fe4e1a6ddf5fb6a0d2c3f8ad349606cb2982537e3a406b225da3356277afdb240d4dda426476ddef8ddda61c5d27972b05b3ed1ca9c7ab6425dd793cb5ca42bfc42c1ad98ea9ace4321bb9bb399d534dff3a01df8495e35d591d811e73e2b4da0d260bccd085307d45caa2aa766ad7fb6379836c640b0fef92e9c317b9c8ecdc410f6e513b30082c292c6731b817ca56985b60811c833111f094ad0b4cd2801309d26c09ece7badf0f4219425b2af8fde5c79d66eb3da5009daf1fb59c7b7667478a8341a24340f8b3821b2d1575b7b93a28344d5c305cbb507300bc114feb26fafb2b5f2551a310edfcca72;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h61f1a8d942b05b58f3fcf4dea810162e9edbc4fd1225c198addc34dbc6808b555f43213a957b73fcd604a8011602cba92075bf7f52c2900f88a1d3addea70b140f0d3651f4585e70864c24486e57fe3144daae44820f0795cec65b7211049b47b8066917dc3179be58daf1c36ed073c217c511ffa5a672220d2bd9ecf9bea33895084e8b4df2039416c55330b5a5a143ed920a9bb0d726c1a901aa9a3dd1d36ebba6699c520dd1be3c0359ee497eda5d5a66dc0103fc7df27e2f36a453a2869861da66830790f614e4c2ad4583b203a269a7d5afe189f01c7b5f7bd4d8056f4d045e53b07c218df23089f5d0e99a27010379467f89778aac337203945b4e7a3325b44a90db6ec39466c85d6092984a6ecfdc6a86afba43ce78a488662c5a58ca05e3c32e8fe05fe4573f43324089a427c54762d9a36ecfed27b144ebe163b47e11da276271718f1859fb707ba8bcbb730ca0342b99b9342b034e13e3f3c7e1ee279d5828b14683eb294878930917ab1ca97f7e3edd68f51a0d77709c5b3c0ea73d80c0060b5a8fddd31fb1ef5e7515afedc9a353e5690305cc4b887904443a514b76d777d8b8d880fd008e430e7b4ee0bba40544c12b9b9477f8ba7c50f43512bb143dc3726d34767dbbb44a4361f459176ddba9318b6a12410da1032ffc039720e0391a13a3a7bcc7be257f68440adb5c60397badcbe60ac11da2aa44a9ed51455b67e94ee72fc1db961f627dd6efd70be80b91a904e879f7be3739de729d24a98a5c03dd52f400cbf3be77500b72cf3679733c16e5e806bdd685ceda5a985d7292b381c0fce32f194fda4c0451b0d76b76ca48fd1138d4ebc290c655fb89726aec4c3c39fdbec5406b9ff3b3e77236bcf7e8433d97664f9096312cd11d79a02a7623ea0a9859beb6018e1597ccf962ecbcccea7197791b243737923634ad1670669527610e9da43e47a01c27f18d20784890da2de1afb9800f31fcf748252da38d255b769cc4b00854716e3989a822502c5fbb4b6f3cd4861b5d505267d37f3f40be30f9f6276f517eda2c1f758e3fdc083266bc59c7f28ac9ec15d276993fd4e8d7be561aba82371c937b4581e1c6fbbfb1edd7cd60b115ac5791481077546f2ffa99aed4c86a3cbb0c8237e6000e8ce5a4ef25a2a503c0880c4b087cdec7a415769d8a1a7fb01401fc1cc5b47bbb202de610417d9a921e9561efd0293ff05e0600638e5e55824efc581668fa453d77e49a581798f501fadeb999a4b7ceceea59366ad92822b01bea1ee7f7b7adbdaf792c5f19ae03ddc25f05a63ce4f344894e477e245560346f4bedbf07e4af60829cafe85430976ea97c898d3fd501378c83314170f35927453abd0792271b247500a9af82f29341cd4b0f4e2caa1849cc3032b1a87800c809cf036749e218405fdd61b125eccf996be1fc81a4b80622;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hce864c7441be7143b82f39f2a929ced25835ebdf00f1564db8f1f49385b20e01bd647b9de9fd47ff05357a6340fc33900fb4df5f31b23d2fe4505a93fa6ced45ce2bfa4a52513861ca3accc274d0c7688ae775b55dde79b283f68b133bad09af73baf7536e5fc21e72787540025e1dcf2c51682a934483c45dd5bb4af9e6db085a6a7e6c8c8cc66d906a4744abd17fe15f2a73d67548dc54d7d14b2d4ce7d75a8d90274b78fd1d85f89df1b47d2a6eb94effb48c03b59c1014c0f605ddfc0fa71d12d4aae1dda1c8b5f052ae1fccf0a4975ae6ad1c7a5204479c2520e93b82d6a2fc4d9062edfa3b7ab3e15efafa82e3473a4f35f06aed9177b607050cdad71fca2072a54978018966c2b8785181b9939152edede0039660a9bb5b427035b454188211a81d9ef14bdca1d74f825e2fa08e4bbb9af8c88fd5c176ef6dc4d05c3ad7290ba2b55d6d91b762a380b24f6da3493a618bfc08c7f51e292a2956d80e2c69538cd93dc8af6ed220642eeccfefb5edfb88707a022c3986a5f3d1ae602c70b8d73766fd670f687542fe540ec9b32391548d6b4f04e5d7134d4e6023b61257455726c11721f2a34b6823c5b665f9f3d7ba43a1ff1d4edd2dff42ce1362cb0df15c8a198afb24cc89d1389b15b19f102d3b6c6e1e6348b12d67354938e3e955ad863760b0206b68b420c61d2c18dae66f381bcde17e4226e5a3f7191dcaaa2aadee716443dfabb6110160e1931b4442655555f5760e6dad565e79d27b0124928805d29319c0e73a95c4447a0e88480e85105f2c250c953e939595b322f27fe254f9b9e3c4ea1199c9baf5da8b1ba07838c555bdd739f76fd643b24a98173fdea19b6a89a9979758369004566fd8f1cb0cd57d6ecc0e1d40e300fe0ad0f27d002436f73f391f60e956e38109fceb53b6ef0787f69cbb615b3c425901fb2912e48c232635cfcfcc04314472ded71fc5d6076f6ed1f16351a0457a65b7079857009cae67d7ed4358bbbd114257fff68582136fe38aea0b6153fcde6abdb5ea3492c733331485f08eda3a8b15e081eee265a4d2de094e3bc6dfc46a914b31cbfa23b3dd6f32eda5dba188ee26535068f78e921bab05ae9719055f55ea29f3ff7b47eb6096bf0b03e7fdba6d7139790cb90062c5fbcc15060739449beb74c46216c95ad373968eae793dd813f76c4229602419ec934487350783d55428c2994f9f9e51c068777bdbc436a7bb2d02da770b6d24ac4920537e86443f8281cc01652bd4f0ea9537c227e5c3be57a7eded5b88c33363959106f11e94884f1d5b18ff284cd61e857a9546a11dceb38c66f7e0c6206ed5b3c20603218d903e577d7dac1a011aea58a88d3e0940144c58ad3798eb903aac1d03f1b229c15106b1ab7fb1c26338f5be64f21fa150dd9a4aa59a5caa62298dfdf6a4e065ac6c682d4583a202ad;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ac4c4c2bdf0e3f4e4cd8ebf09044be9e17a4cfe8c740afec565236b7052726215291ef7b3a3ab3dbc2d37b0077936e2d65b2dee28147f8e9cd03b5bc9133c052ad314f07b915d381d5b52d8e4ee169c42c5c471457d41aca3da348c43da3a08cb2069c240da30d4069807e1386600ddfa969b72f7f0eb4bb50616ec391152630ff3c9de2ddb80630359df7093dd74c79a30511e99d37bb5c243e209f132445ce1f64de4e03cb5f4130855efb4a82744c7574c6469028eb5ee9c11339d0e8a8396af2d5522ac5f944d1e2fbb3821115fc74b1533ca441eee659b388f5904a90a95593bf672e7d29f8395486c88d4df0e320a734afcae2218c0b695ca96696f9a055aa4949d91b8ba7616f8514e08ea5e1c5d32c7128a1328218df47a04e1fde455ce2a2621a58ca5fa2a086d306120575f1f8bbad4587afd2b296c1c1d58745913a3323ff42c8b94d072ec5f86e8979fa207bc199b701a8a2e5799be33650c0f5d6b44f0bcaad7975bc06e209312ed890034d50251ee41009d64a54686742d49eeee53241c9c101d64fafc4d13a7aaafd2c4fb75e17cca89ec84d3a24143cd17dfd68812b2c0dbb6b1d91aecdc064be3dc9d85d8572bb9f8b5527d0c7572d1147bc0ae570bf29cfb543c36859bfb1cb76901c1d045c27984242590509b433394e25cc750c7a48bef4c2886346623b50095a9b813b5d427ac478002782a5dbda2c0fa12adaeec2b2ef560a013b636c29afd7b0cfa5530a6bbfaad6451c8bd2a20515936b53068e4f9eac081841adaea40c556db57a2900dd339debaa63a8d2e4787712f2b9ced9f142a89319ef2218bbb1d4249aefeb4d182d0d6479812a1e52a26b4adf1168d3f4dcf505baa14b455c05a72ff360b0787460c22977de688e30e2796940bed7933a7a2b11dd0c9f208f50d151c0e180a0fa4c2d6533902edd40dc223e1c644eafbb531b294de0ce10764aefdf2e631a5fe286608a36f575a696d88c7981043166375203a6ad93d5e38fb77d04dc11357c8099cf7932cd242b2f323a8dbf47722981ea0718f32dc3f694939ddddbc7a0126ccc3e700bc0f695555ee01ca871803cb6c8192a3a5f4a033c8018dc9e5d5f429b053a4683773dfd73ce3f524d47bfa2923d80270bdfa1657d5e65309c469afc60861448db3fa95f9b4778b73f4776cb57f8e9fd956b8c6f7162a95d6f26465ea4bf055e1d4f40fd303740b961e9ea85043ce214e3ca0579830d660d0012e6bd94f6963297c59973b60c5dd4c48ddbf37d7a60a32250f1619bb59b1327cd6ebb09cdf54e193805c1e4740f7ad69ff0d28865e5f8271060500a1fd9e23ba03fd92b217201cb434536edc8d2346091e43de468640da59257dc32e10ee9c9f67184ee40b41f0f1ed079728c7cddb109a617ee959c567966efe7122d3e1c63100c95a95cfb734a92d915bdf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdb692ce5b3033436aebb91c54d853e856b85c8dff24cf0e3e04c16d0f5e2fdd937c6945df56a256a892947027ef69d5434fd490d29047c58788affb596dd62074b7ab32d18fa12d66108f03d0217c9b942668a7a8d510153a445f1fc9dd57757b086937abc9eac4e0c0a7b3b20cc03bded47d355ddca24823a530a68f2d4ada754719fc92dbf703eb27e081fe5ae5cb5c90161559bbd8fb24456a5ecf3188086e28d3a4169eddd72dda9c0e37cf4c439fe071a3ae100d86d0579bf8163c5b1e38c9d399e413a59f9a28e71e8c685377f8a6a14df2d552e5d67b67c0e794d063dbb6f57dfd4607893ade13555924fd80fbf4582679e18711e610892ebb62377e5994b435e6c9193fe3b0f11a5eca74bb85ca6db66764f39a6756f60957f68e9d02d6d4350e6ef161d70f8f8bf675f8d804eaf02ff0985b86f2314fc046eccbd0d6cff323da32bb666515b6f655fed830e44de0eba1544fb918da516fb0d9cc5775b30834a99514297edd8dc4121f2f2e33792ec3d294058259ee620e19531fb117d68d592d671c168e09b788f323dfff34a495a5eac9bb146206f58ea08a34ed003bcd46461a29fa96e31bee35ea6e1b8307ad1451da16e0031b127678f0f01ac1977febbb03056ec2eafc8ce7c8e358af14183d967dd91f947e65a7978f8a66ddb64e26daa67bb4223e39f01ea1b72cb2a2a245441cfd385ec13a51ac9305ec370175bdfdd29e6b4ba9dee8100d629d101ec0013afd67c44351d7317141ed53c285d7ba5e6509635ece810cd8be4ad3a1c65b3d4348e5beb6d408dc38851f112c060cb6261f192ae8cd67408309d1dde60b7227049f35668a11a99fd3122948dc2c6bbec7d6cba0da6f89d0ce41bd507b7ecdef888dd595db18fca0af658057c872284d994b31f73120ae9334528c81873f3860c78720c81615952f2ab049248885989be2e187711887bce6ee05ab8891e9311c4e906a4f3319f5ca7c0364d1834907e85b5cea785589ad7ec510f844bb2356b0571929aa5f2fd965a563f47a7bb5d5f8ef15f4d04c569d476867f7a4ba54b92c1c78eccb2aeb490e5bd3ccf3d74b341a685f83053dc7dee3fa7790ca34386a6e57345eab4a13b9ac78a891ccda5b70c4dbcd135cf1d38869b8147682d589d028f85209a4d4604d4f2990f257653a4ee078b22736d004604c2475bdd4b481b45aeaf1d1676edc34358eb54ff1f14b418e216b1dfd558f37e902fbe81af580e5baa63ca0d3e48ad83e79c85e4993c01940f8c6894ada6ffb2af8185358edaa1c73b9cb0eb6382bb8990c71058705cbd7f5303bc5601e0647170be1f6a18ce4e934f409e7b84fb8b9228a7dbe40e2e7d7a99d7092211303ff9435ebea7703091a049c91b6ce350191dfaaaa26008f304f5ea85b1ebca89d982866c53a0740cae11bfa907ffbfb6977ad3a421adbd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h124752437e6c26477168b42a4232ea0a766d7a47d03d796bed6c1dfd8f73c771758b248ce7888b548a8305f3b50c73c6536115d2daed90f19dee483e61c2fdf1c0f88b31150b3b0ebf410991790e60832b7164b2888866726635185f1a2d7780c97f7afab1da6c9cb86527752ccb31a133848d0314e8bdb4c6933e51a4c52d961c5d6cdcc688978f89a5cd077398dfb24a8c8c157fc364741218953ab13d0ba288c1c591b6ccd2ee8f52dba7e9f6e3463284d987fcf33dfb07e76e944505bd54f09ca706dce8aea0e31eb401bff2d3fb14c30c4b59cd61efedaee2b589e617d4c07db9b5f37ccfde16d93494b850e359c59f65f1f1babcab3550fc628ef660a6ddd7988c1f6d6e6499e4d1a46953f7f5ba8986e762b75990bf361dcdcb5f47914f7f8c448b4aea82fd1dfc2774b68eb88954125008e97ea2991b9b8d4345a19aae6f35686c4e819ad0cc0416f7ff74a5071147d80cc75ad7790e488f7f2778d228e8a3ca399a5984d9705098e5bf29995ff2d39061c217e033034d8ad155f59b4e40d38255812d5d06506ed01d5049b0f8771ea37b2bff69b6b602e22688938327e48ab80cb712070375d55adfe773e746cbbfe5dc02e099c6cc29e8fa795756a67cc4a07ab6e48f36a6e3d26ce6c612476e6d84aab4497bbbaeab419ff209e7da5d21fdaf9342f01df2e0a3c884529bec52ef545671430c3a2718fba68b1140773c7e041787df9222ed08044f589fa93127432cbb135b007146f040f99e8cdfc6287880ce083271e5eca63de4b4bf99deae5277c05ae1303d731b77c0de00e9d4c672c198181097e76e11b9df26a8ca47e815830895297bc5135f36c9c7ef7e4df696d4ce4337ece543475ef831d741ec37b0c4aa64d0bcc5f023729907f468c93e6255bea47c48a948c884c6c5d1607bf7fe8fbc64fe85d7118f313cc4fe839282d5374eb1fd9f954683212903a13e44153fda28ccf1c4f3e220284be67b008658718027afabc0f90885c00430c2cba519756cace7c67f8eb6fbea4b09c6c57d1b21f4934036717dc6d437974db3f8075f4c7b839fd77903383140f83bcdaf8b173decaf2ca5a31c82ad9a40672464b5f9de25b48806bd7b69960c5f57912991e19771eab84487ddfee9ab66fea8680296227cfbbead6942f70251e45574f7e135b6630f86f1b065a755d2bdbc0cae9680ad2424a8e16d1944a5abb45455a82c7300d8c05dd5cf6ea37a776b66f9af8c5327ff0f60c5855f4f49ea33046f42be4505cf312756012ce0ee9e94a08b0ab8071223aeda4b56bcf383b4619c70ce6238a25e5db054bb5b46e3acd3ef3a15db5932f03552aa3615f522b27e005bc3c8a2e8f543688a3ad4dc06509c8ffcb1034b4975015e8280402503bfe11ef1d4330da7c4c845f4ba9c89cb4312175b63038d971cd50319b2ef911f26a68198e6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h84c0428b895086abca9714fb8ea47cd10d07ab450996d7d0bda0983495708b069175febf03578d427f80cc4f17f5e537fd6537341426d16f281bd1dbe6753b45912be974eccfd8812fd778f20267eeee5594af068ff90e9a3985ae834b35b8b7ce4a8a1dc8dac657d6c9aafcb5a352fe2fd36d14bdd4f5a03bff4f0cccc014839d18411b0a4162d66ea3013e927b48c76c5d19116b95b89615e9e828964c3f4bd670608c584d5c8baaeca3dabeae6c4628aab70d3ee29ce0e95f5718e7951ee89c75e4698bf6420028b095fe9f32801d6cb3b21102219e522a02af457d2a7b917f66cff237d36e7c0793094bc249e081e477d82aa746c74e9322dfc50149354feff8b7491c6089659218e1fa09b30878b8bf12218827c0c820e6279c7161f588ab138197d08b212b0f0b77f00759cffddc849425b017eecfb793bb66658319f3767f9bb1f51519af1d21628a657ee0065c4baf1ac1eaa14724dc6f63d9169f46ae5ad8c6754d091a0680f3c1c8e1686d615678de7c6749a8d0e322ff1f8c1941304fc70c89a204f96b048b174a2617435a1e45153a07b827784d62867670c3516c22dfb98ecd0432c0b6124dc34fc625086d6eac8f00da940d859dfbdb6c178fcc9078e7912701bcd3c02a79b0b4d98ca9e8bfe41efee92c544b6fd5fc96d4cecf4b02f1b0927084555d88e1221c7b60022b867e34fa454d75b23a71f63360df7472da00f24f9492eb8b55e9fbdbf31fa35ed8b1ca26030e9a76e87352c4eaed1edca16b4dd4ae955030b70b16eade764357c45df889bb9225ff61f0d1c337517277b0d04878390e0573b2196f32a12f4b76cbd07ce4c7ababd26964f99d7e2242d402bee6800aa1d2ef19fe4a8467bd86edc4fdbd06d3d8c669510b8ca528f83c7e56a0a7e4b65aeb9b642532312c4854d233d8e7933adbe50e055d9e83b291c28891638ed275942d7fd0b61f045f75a9f69be58c6f55c9a1480500545a5c611edfebe7bd815e7edf286622f9196b31843acfd25b85b00a676ac9a1187b12b9400b243168697b1311db9c50b35da674174ad4500d717cdd2e42759cd3eea324396daa7c5794bd187caf0e2b0a62a8e5afdbe31fe263cd8ae5b6090c4164140dd2eb0df48f4aac5afa27232670ef9d35f3e848925ab97f77c4a55926164ad92fb535ee0faba04d6e81ecccced3480a28e9db62648aad7832b93c67e8d218c4251ee018a3addb0fcb6aac67e5cddce2e847dfad85079f08469f67f645d97bdcc6806e00b231644906f6a25d0d46954be3fdda6eccf75e6637284345d21035a9791df79f73e0da473703d2312ab1f8331bea9927b8ea1d5488ed429cc07a0d5f8a14c493a2839d6e5ca39f08d08e0972c7a4b6d559bda3bea1aa17c6d62cdaf163c3cef404a5ca312bad5c4c50d48a3e7cbedda5b7f6b53377d8e99df577f9648e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h14cda1726bac132f37e3fe57efd1c8bc0c182e25b7563501ffdef7cc68369bc345e38e8bb26b45831fbd4a3e404dcb76b54f1699fa0a05fddb5cd5c320b57db3e30e377cb5c273432f9a98ce32fbda9491d5758f42b87519e9e04528d2db37478edfaec112733884cfee6ad68149cf89a06cbb7c707badbc1d18dfee383d385772dcceb385cddcde6f959e0e1a598cdb6f88b3b6b6058f6a581ce3a47fb7ac062612cf4dde35a9b7c0fa625deaca3109ac28baa05a07aade59105e9c99c9852dcc51c108094131e93320a2b63dba0e878be7f3abcfdcdd6684aba9c44a42df013cf69dbd33bb660b4af560041840e1ce41c98a586950a79653e12fd381bb17ce8a921809d8a3b5507c1075be947b7faff059fdd8979a027f38316b3f660c20c7186c2859631606cb27d0aa59199926e79e409e86f1852f4fc1a310c9036d7ab9bd25fb9d59401d8ffa3e2622a2385180ca291d32abbd37e98dc054250a4bec771b2f8b22083df6be83413f99d48e6278fc7cd3464faea9d581dd74a24b8f99b2e4890154e479837cce6804ac4149e94d881e9583b8d3b83082edca488ed053ff8a3c135e2fa7e8bf5991847e310aef2323b91880b527c8f55cae6877024b6b8495bc16c371c8b33eecb1f2258d8732f35d421969f5278f1991ff5df7df1b6057414dea422095717de235b15b9e651840144e67ff108a1d7eaadc8a16cad04affbdda60d8de22252c83c9b4c8e85621d46c74c7b1ef4f856d80a36dd07a9bd4347343bf52aabfed4b62ab815db8f5632a0568a11c0002ef24a978b7ee6ca4a8e3e8b78e5d6993986ddcc92b8f63ff907b933f2b9e3ee855aadae4e26fe4638a4a72e2659111040d9ef46fbc4e260cfca97555cad719005b0b87f60445792b3a36cc3e27d489c2259cf3cef99eb264d2c623981f785501d968fc3fd02c43f7d1ca39c9f8c4881b4909cc6612a70da4f3015c4254f2ddabd8f6ecf4872c41f28a627f63599fa96be5415bea70894a7d134d4ee580031dcc8eded053145fce2592aefcf50bfb626dcc6958d560063f3f683f94c8291b5e7b9f8bfbb2dcd77fa5acc868749ac36707b51a1421e94b6817893308f16a77637631beea0dc727897217da38d3ffbf0f315cb579ddc5de2f8ae8871464d5c98e180cf4a6a3b6e711be7b76d2420b6a0ba68d9b1a237009dc1705983ec1f9043465e9538dd8143f938ef9e2e263f759d3ef01022281c30cc52ae007c1291fca76fda17a659e1a097bc649e7b475e1b77f54bc66b9418c995b589d1b2903ee200662e39aad17161bd32eb9307de34c5152d80f91f6d962decd433d81e1f3ae793005a754adb4f674a38637e8fdb1f77509ed28fbe2bbe259dc1ab7f12715c04f6f2d2c12ab1d9dc8c4f0b13feb3c07aeeaa4eb4f74cbc0310b609105dee98ca3d522cc70ae9875313d04c01f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9c728611a3b49c2e07249042a72c49df70cd3291862ce48013eb9a86256bf23ed3eba6b7ed54de7bda1d986322d5d950f83194146cbad0eb587407d49cdd2bff9b28fbff6e240fed070663c9de2c55bad0897c527220c2fdaf1a78dcfa2594e1692667f50c18883d6cfb5dee533c3877349d1a942e8e8cc0456f4018a8167e15e5c83eaaa14ea8c26fe81f3031c68a4e025f7290881648374e97c1819e3f0bc5745a281cf2646904d55a1624a0b0b1b6565b77d3f83c53bbf7d8e0f0d6bf75ba58ef8a5132ef66d8a7f9fcd0c38eb3259fbdd135edfcbd1f85e16aba88e395001e03756fcbb9e76f343f1d3ed05a6631313bb7f6dfabbfe30b1c2d2074f6bacce0101c997055eded1e0f8f8122d757d0e67612a58fda3692a2a232188629f7918de52defd9452dcb882074f2807fa81015a679f1375a5553e7124729108afdaa904dddcba434aee3f168c438f532e0518a01ad2aefab42c5312a5842797cac39a9786259d3f3f2e5bdbca7444f0f5e908e15a015040e32bbcfddf4e2b22ffffe741df854f66fc21b983c4193055c3d00c3ff55f69a4609dcded64efbd30a5befd403369bf3ad5fede256b3ecbb0279e198d793d3007caebd5a08c42c23e47dde45c5d924e93e638e25eb03ab4d271c4f2b937954abed7f50b5cf75be974cc4047128007047f48b71b7dbfab73b891d04bc85a9be28884c112587f84cc330c2979a74612d3590a28341699d31fea8dc48d90f21dc6c9695318ee755bae7344ee2bc35ef7783ad08bf95591386cf84033602a97c55359aed33e1769188bbc25b423f8a0b7836f9270aa2c55aac1f29b703b756c2ea58409b252908939dd37a26b0cfd94b75812628405cad5546bbf349636fd544bb460e3132cca916f1231ed508c88c87f28dc1c11dc576686150908d57971838c30e9bc9a80cc3048f534ee02ba6faf7f4e552e0b3e06bbb1ab607b71ed86e65b3a7642b9090de7ac047eb9d4e8f1ad4e9dab7468b55a41d6ae65c9ca199958271f8fc7a2f97eb0d2e5c686616d12c70daba0f42a550c0bd54a59a8f7ce025cacb14251def0804d9c60d0b3528251c059b7ba758b329fd593f25ee65685568eee0d8bf08c0853456076000c04809dfc4d65a374024bcc979084cfe198b8271ad1f967f131a47301468700920e0af2a214e207b9250a4fc682df5534abcacf50d91c22eef30061f15af239fa64cca0d441bd73857be0ba0cfb7500531002809656c12eeaaee4747a45a97072453bd8780b2b3cd5a96df1ac6c77aa78bebb14e2a595b7f3a677d5cf7b0815591dee3def02b9dcab0aa5638727782ef04cda1f3cada710d0698a9b59d39771ce1a6550daf539b9f40b2ae230827f11c1fedbadba674c4465d42f936d0c484601bc37ec0e5c8fe8b8e93d3b1fd57972ac05a729600ea271c0cc557b8c4c0415af721;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h309772317cf5ecb0dff216b0d3cbec410fd304128adb9d468ca372194c63703debbc905353e01a3e02a89ada195983f6bda9789e6243d0bf0942803480cc3ac5840e1816aed2753a77590f3de946dea6a66001885e22c2c9388059ddee63831cb4fa170693492923cfceb043d095c973317036e796da3f33758ceb6000e15e1958e427f4868fe6635d7d0a6c3e6c423d7277c64d7671d1d9fd2fb21f4394516ac407f2a052b8f62e93c5837c6d698b8a38444fc042b0caa7d418af02a4f6d7984507ca21b9ce53ab34ec16e4e5becf0441eca9e32f4fc2e72b3931ffa20b8bea6845e76bce15a611836a944a1fd8b521aee2b27a08d30e3da3ecd59e5e838920fa3f1cbdd7f5374630af149a20a921c119c83c779cec4db247f64353d948b74cf4d2d84464bdda87da1682331e776e21b4d6c749360ee53f3076c502f6b63513f50d56f1468d344fcbee02012a3c7d5996d5060e238b423fbb699e8bcb54029c5efb0c5c48be8fa493fe4c2266ddabe6a6574c1eeb299d77f5fdc7172ba07ad16e994a9a9abf8aefa3d431276efdb90375c0f602af0153812c3495cda67e8b22a0c21160a604de4487702a03b8f3db6358b7b66215d15b43dc07ff47484d3c0f9dd4d91e377a105fc0f6c87d7c56abac02b5379b8d38434e368753d543bb58565dc033845dabc57ca6cab5c03fcb6951b081ec87a413a55b25954306e26dcca8287da9d260b0347eae7616300063fa977f0c8568bbebfbed1b42db98e28be9b776a9971b47f1f467f7fbfb89a5a77b7793126ca59de9ecceb81c973ac2edb2eed3f49435572bcafa74a3e03b683f92c941d84f8f33739e84a97b19782052f6479ff2417d861282d2601ba8da872715adeb53331c3911fcbc1017e62fa8185cdf8473feb30d600bf74095176d0d816f99ea104ff39f0d1bf53d316337221b48462b531f83debc4ce5d9a3479f1da993f588d95ce008317db84d0f3987686c9db6f4c53d3778fcf6a41e4746f935d200b8a456781bdea1fd1587815c2b3262ba8b177520ee3e7eb8ebb237a279a665077e6097179a50c6aebc5e1d4965012d6b1448a69be8bed02ac8939f0a910846b63ac1f2b08c871052dec0676aafcebce97e375a39dc42a3fa544070855deaafa857c59db7664b13fb78be9c28469d94ec06f65506a49802cd359e3953a68732b93ea644f9c311af58c9f0d79e0f91376c39e31e3c86269d3783e5c72dff71fa4772fa1b082e648cd76470b34fb73503e56c4b3362c833c04574a9f473e1ed0a829e317fd1402a5c9f255e28a09379dc7b74b6fcaa18c38114eb242e39d905dc171f00cf0567587eebda88e3e8e586807bbc7684531ef84c8c1be5961080e88f8919e1c68cf3bf13f522835221130c7c124bf2c3baa87743062492ed3d0622ca239a283daf8e3aeb4cfeb258fb1e8f360a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha8bd1c1a50efcef58feec56be96969f7cb84be013ed971394e08e2e12708a156c947255a4d0966d8850ede63f7b1e69210134794472aaa4e3f81ab59e38b418aa1d0c75862edfce8f87321e66186805854a9d5e6148cb48f728fcdfc8b5488f3cb9453140b844f2245fa6edb58f2761872c68b9c82fdb56d00f39ff378dd9fb6710ef89df318a666284fcbfcbd87027464cdeafc0ebfb585d16b0d79272679b6adef20fe7f63fb7ef0e9f79eea87df06f1dab0994d92ec2cd54065f346493b698fa070e97a5e087bb15e1ab66dfa6934fd135387b6fca6dbb64c4ff79bb9f492b86367254a2d7e715f938d35967072b2087a1d68e03f6ed15b94595a3676548b68113fddc0dbcac3d71ec9b4285bf4b9a84dbe6dbefe193cea038462c824fa69eb11c2960e284ed49b417c8f3ef34cd37d31e1dbd2d31c590bb4066750678d4e1c5a4ec31d1875857ff33fd6408f66cd748ccfd2743c0a6cce2f1345e881f2bd260f9a65b8f2644fffcc0bba02517ef01e873c52b88c3d50e0f66dcf517798dec6fc07076c7ced16b1ad0e6b686c15fb8d58f906e5210dcb134ced772b71b3eea8f42f58209380f7737398d5b3e473484afe7760587c7ea26bb2bb510d16a637c4ded4a1f49fd2bb81b04e4df9fc6ed93ecf01bdf6a5727bb262553d2e2d75cbef92691fee7b73455a6ed7d7d063dd674a6ef963a1474c6a979e508aa3dd8ece372b3c43b06a733c16373b07f0104246957ce3969e47936d5360135df1afc316c8770fd7cea224f5e2609f6f82869f37f0dcc659e59ebdfc6b065c0eccb950a89bf178b5a7e60e10c171cb3b23299fc407284957fc5fcdfb21829a5087f9e76c55091b484a77b50768fb5440582173117f234d154185aa6196ee66fc22fc7c457268a5abc462c15117d79666238e22114bb6b70912113d8eda71c74f4be7e6a08255d32b317d077923ba06ea14910b9c7587af1df93d7916e00d2ef95eb5adb4c28b104761e81b6fad1e79cb55ec00265ecb9a28e25152b51d525569e75cf9c0f5612b45bd635dac274ab1c8b99a575d0d38e73546725932037805653ab8dcb9909c4fb9ccae1ae2f48dc2a7895dd9d08803da87ddf86cffc66fc01679fc7dac0dd915ac6d85dc724832066f72cf42628725ca33fc8657fbdc9fd9a8c246145a4ebf8fd0d4ab3a5948060a412632bc8afb4c7fb963297544c92d62840bc76e41a6f0eb01f09622c9d146ffbe418c56ef656b1714afbff9554cf0608b13a4b7e2c2ef91cb3f99687b1db85ba5571c362ec14d573cea65df12724afbb8d913843542f6e1ec2d617f78ebe05b2fb9c9ad8d1ebf22ddca266257b0ca64601e7d9798a7811a68f9bc7918c95166f2a33d658a543c1475bbd8c5dddefdd35204bcea641f681f5d39afa61b1e5574ed545c7ac9c3727e4599421a5fa903e905deece759;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha5a6ed4efb5da5f8deb8d06af266e69202be350db89806a4271dc61b116a31c6702ee0c204d3c4126c27d8140f41139540245127a1da0533e87b5b9ae6ba0e51538d3c992c8e9709856d6ba63b43f23aad50da4bd41d3d145530ba69f27ed99ecdb95357f62054d07c861733c16803a69cd49099e0781fd7dd481b1aabb2afe80674135ecf06f0dd94853ff4ac2144240d8ab47695533018da3b2e056ffbb9009512b76ddd819be80eb1666e07c2352dc3c76ca5109956ff067022999570fbdeb5136895fe6b7e8cc36e98a94f9221a8c41ebc4307e952e624f744a52d43b5a9ae3c6fe63fd258dc8956ed1bdeebb8f12be5b00f5fcda3b5beb12afd089b28bc46a01bf64632b5b1271b09d0d17a9f19ebf957301dfb22d47570a309ce3202ef15180534e17b02b08cf2b55d0e80b909922e33fe6c56d5ccd3eb850a03ac79be469fad03581cc082242fb25af1f1a866f16419ab8e5bc1b55ea5eb2eb620208ce6acc349b08934d524037b3c48ca8d58416a8460f501d8eef03391f68c32c73278df9ba8a00899e6b1682b919cbe466d6dff5cedf7d423fba29b3ddd44e72d0c22b1fdbd479709aa288481e8eed31baf778a7a626ac35d9fe1174536d43d5a957c030f4df8840d59bfda0475bd305472481d1fdcd85dc58f5a11323939f1287904fc1dda05e5245b035fa487c6ba68b353905933714279be37142f4d7cd61755dfadece8e881d513f175adacb0c58cb4b35253fae0daad79c89bb3fe636d8058b1cd6a324402f4b00c694acd248cf35337adf997039c12ad7b00eabec5064f36adb122d2e05aa95e9d24b47375331433e0dc5aef0c9c1e60a41dcc60ecca68ab85446c3574de7ac655ceeea1b552a2880a2c6895cf79a9cb1ba86c5efe24ffd2cc5692aab38f1814e4bde2889cf2e89f3c7df1e206c318332d23eb01e66f3e8a7d3421110f1bdfe824fc80e2fd0b0cb0d566f54ee528bf1c9e498d355afb3c0ecafe8fe125f751f4366e882bcc17a15cd5fc7e2abb41692d5d247913fee1136721a25b8c61e892ff4751ff0f878e9dc27f712a167c7c6fe676fc8d7d3d6f6e20e9b1203ec0abc128f23540836228541dbe28b36cc343989b4192c9d2b4c76c60b8f92e7a67ee964f9ed58aadc56ee4d74b82020c6c50e4929e8f0b3414c7f8ce3a20b2bca1a6067ec177042cecc1b125c00831d1a576a27af7f255d68dfe34248e615365d905d63fe99688a3b45d95b397774f49def8acf9c1423ec6a9b439807585ff7877d362cd8fb5f42a56a7e89077019b71b9d7c78829c4c731917e8333674a2e00888aec2d19c6b56a611a37e6a45199a0d5bc8c1b737439252be7fb7ad8cbff985a322b3e0a94e9ef0fe2b55fef5f31428eb7960c5d76333356be82a300f4b7eb44fd44f2984f657fc00fb744852edfd8f5f6b7917c3617dd288f1628;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5272a2852d99e3f56a48eefdb137d1303c9d05505a822651520a40cefbae6b8cebb1c665cecdb7e339c3d59291943c6e16c581f7ae50b595f96f9419df9fafed84a9020afc40748784b2c7424f768633d1284576ea5316fec0f10e66fcba2972d37be5da4d58b4657d74c4860733bbf76140a1c361ffb17082109728ba5b20c5426b4a21f2cf481698333ef6c0d62b434953674c1402239dce4797d240f0c4b73b0c2f2e17e38ad96b635d5778ad30de5edf9ee33676e33f8ee60a5d7d9515f7935ddf98e0fba25bc98e0a67856adf7f192641dfb6cb893dac493042cb21817fd2a187cbac3cf5c08e041e568e157d581530823516db7eb243c5594163cfa702ad7799c32a1f1e41a254dfb4c61e5db2aba0adfedf2a14adbb06c813cd8bd02ef22bb878a75eba26e4ac444f4af0881faf4d5a1c245c5cee36a4c8890aa8f115444820bb61dbe52160fc8c5ffabfc96eef1e6e26759679108b1fc6f07c73f15a081e51de77b2fd78613ef23d6a98aea348fe218aacada53fd3b90098419cef5b1c34eca7eda1461a6dfa827cb212ce18ba80dc1ddb314625da7135ed6c8674032794debe45364d8a51ddaa8e349cceea93defa6217709fc2cb6fbd9507f47218ded0c781d5301db745eb0d68642883e3053c871c7eece8ea5dd0810f2c2473c6ea3c1a68b3875b6f357c3cd858d69a17b6b995bf06495a0f77e38fe83576c8fcfc08cd24fb8b8776dc6e6589777972c96faf3c6bc1a67c091e688477471c1513531eb6d6584c2499c5300d773ecc2c694606ddc152404a87837d4adfc41c23e27b190aba9bc8e006223897bb95f6631ffdc578dfb6d2021fde8f7c0e3cff1fc27c87c50105a5e6f33c6b97f53fd11b50656fd0964fa9108e590f2f9913b98eabe147b9212acb96f5f19e9d555912b2f6b24093de177f5bb51d956710f377b93157a358102e44157e0e90bffe185d48cebffeb7391229d99530f773117825631a94fe94d31f19b0d04e6eef64ed6573d7a2c05f710254365c532535d3c082a41b29668ce578ed427267dc52f1b0b8668d6ffcb5c99f5c3c5fffb6c7c9e915b5a1149b8136721e29c9fc3a342ba781b9de26647559d1f90119d8acde0e42a1306ae110c2719a5609d575ce201fb1c95e1a5c60a1283c8baf6f062eb0b43509e295cf94e46e887afbe1a7deddf444a53fdfda009e76cb13fe219acb37afef1647d7b185c04ceb864808dba2e4d3f8cbe7b22c9da6053cbbc83356c94246301325717b654d15c9e2f3d915156e2f6918de2f7608b59efe3b577e2257450d3bdfd6fde987e241aabf591b04f3657e6098d3e7c8c67b9c7fe72eb651d682252595814042453090234422f48b9f754dc9077fe79cb8785837e041e799b7c790ff967522a40ce2ed58ad340e5c4db51c342e0655ea294feed8a42024dd8c373e5c1f0ba6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7c8388977abc733c29dab934d8280731b19db18e9edd2868c1a4425f9c54196c56f2f113560a3b7ea57926fb731f4099a68558f54d51ae6f91ca79728946bc5c2db52647bb35ea4f32b87b3fa1ba808cd38c7aeb7e74a089a5f74baa46894b69ea15030b14fafc839f33a4d2ae06cb0a3814c5ec4ecaa7225823b39710b224f0b26adb00635275ec570f410da9f9e435bfb64d75ae0f686e8ae22a5e3b13f9a6521c854fbb123446511bb48c3c6ad2460677b6d541bbe0592377daada804a6eb481e472e0c0dad29b2a470f517225f3061b14c4311ae3587dc90cd02d801a9801154b0448bf204e58cf9842a8fd44b83eba01775f6a651193cfc50a8fc6feed940bb4c1f9f743ec4e07d1563cad1685b0e78d2fff56a72d0c25f6cc00a4c3cd2c279426f832cf9784dc0e1920654b7df83fcfb03f957b1312b6622915af395d887a449d46e17fa128b8c232715a776d955cfedc6c940bc7444b16b5f02eb3b026b2612f8db160336c1f48b76861a9938d2e41100804708ec0c7294d9469a13657451dad9208f74dd15b5ff38312f9de9c8fbb8bb4d59c6342875781d96fccece8000d704a689910a2fa441b3aef523e3e18d9ff5296a21d1a684fceb77812017d55f84242e2e5611b219f50589dda0854480a96114b5d4e92bed8e267e77fad0621a6c91378d315ec0e4923dc187dc3cee5600fe57f01f21d94e2c1e2e0804b6b23b7cc3b4cc903f9ed1e0281dd5c347e46af97be87c32964784c8c925449b86c476c82a4cb8d603d6c35b1cc2a6a12b43660b0689573aa86fb38b36a68e6d2d2aca6dfa341a08a60d011a238bfcc08d8b79cf1d9f82d1a60cd7eb09f4c9ed42b4ae4fde81e149294477f9537edb55f923e21a38b40dbfe120c16bfdf430fe0aa5cd17619547d1ab8bd9645b9dd9dd2da53584ffb641ad48edad3b552c660b90c07aa5d9263115a047cdb3eec183e33776afa1b4b00ebe4de59215cf1aa4c3cfd7ab7953d979374b1f3862f0f23c8c18149f4e1547bb12521af694efc9d5af3eb4a17f1c3624ed56843629f94dc2daee9a722ca396f429752adb7edfbfac09c6c365290b99fc44e2771aecf8d0ed361cfd1a9923993b36d3a81d4aa0b92f8d8260e76b8dbc920b9a10680ffe5892094a96d619adf3760e15389fe971f5fa05f8d7c3c680b2b9936b06e8548cc0c28d75fcd002baad2f147ee12d1f155b90c70c8d96db7067704cc266ba388a7741f78afc0a5492b3c875de48403aed3bb58cc880905a9981f182b24dbefd5956518220001d99e8d939d38b621589c167e0cb52289a286cd168d62ab8300500c84cce1c3f09645497274285603b71e48f62fe7971a12580a37bf2cc180901e3106e0ef9a6d4e69fc2c09cd12f49415ea6a1d00368c49c09d70970afa91a3131ee40ceb558782375c70ab637d096b1bc12e15200;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h63ac0cd1e728f05104ac094874fd8e501aef0eefe6a3fa326b4aeeaa43feb27026af400f20f2cbdb2bd962f64ab753929963401d2438a3779bc6e2f5f329cb09c838047ea03fd930c029dea0d9e8ffb807a1a46987d421839bdf73a757b1f03311d4f4fa365ee44e8f653a7fdcbea365428833f193c08954850eca5686e31b145e3ee97cc56135ad5904cec4062c48f9d056844d32873b9ee28fc776201f5a9947bcd3669827f0444935d2b402be4be731dce84ae54b8fd31fdd7b189daae3ec23dc72f528ca7b2fabd7a1824ffa26bbf2301103465131f704935b3364ce6309518d4679a7c43746230223898f87e8be60cf002198cfc88ef450111f1cc37e9269d34a964aeceb774047fa7172a4cde982d4a4c0d5588e827309a068f39916a3f9113e207a9c7b855d68163314167e9f76c29e9d1bbe3e4abea333ab8841c5c9129f66fa0d638115daea481f22114d9d01c6259c7200b54bc245d37e4e84407d2a7ea281b578de3a18b8383563a9a3b3110b59ded6f7be2db7d8de35f385a76de54750f9880ea4c6ad10ca45e85d4ea471603b4eea5b19c828c4a44d661981a807e625dae54e17eda2ca7290ddaad26b4487a4f0f4fc061035664c14cf232b1f31c891d36eb043c05dca270cfb64efc4a4537eda75977e44ae5e82b79c8b78a0201bfc0d9607771f9812845a978d02cca3f155596a5e55528916061553df8f87ff75da485427ac9bb306ec6c48f04b50426fe8ade98bf15435e9311b7c4fa122874dbea019333f92b2fd4f0f53b61ddf344abc7298b02f001181a12804fd4375d8410d5de9588ab2e2d96e96d1335c041521e71cb6fd364ac81600cf556037cc6463525a271ef8e85ddd387d44aba65e7733730fd9f56ebcca9618db32631c95640101d2537c58a9fbabfe6dd8bcad8efeeb4cfbe6673b8930c227752cf8b7f5b3ba598c6bca23a062fa6ade39e91b618127b3e709b24eb83c55915746454f117b2b17aff23ac69500e1b2df048de76cca06fce020009c2d9cdc6d38cc8ba8c98c0566cd34c99452f203cc98c59b4f51b497814cfefc96bfcfb65360631325d34e9836cbc27af0e91dcd4448ce9de24df43a70c295c3162ae4bb6d864e0ce6a44e742d5ba0494e068e2a36f314be330f42af8fa96a786cdf850fa74660e8449f75ba6b0b6e64c08e231146f87f5f582256a3460b53874d947f9900f00f4651c6957b3dd0eec8592d91f997697e5484f3b8b796900180df76002572d3e1703c476490f4507ec6aa9e21df2aac70cc450817200b6400c97f0ff38ec4969bb490e487ac36d83415a8ec7c8287abdb1f01dc7ecebe3a1dd0a3f1a01073644ef1c561076d64866397ccfa049fbd15109819e1f29663430165a3a97809ae649db5cbb9475624bc9b306313852b17ff51f37288d986b0349580adbf9f882cce2f2a4ecc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h581949fd285b203a0c7a1488b788510aef531b16dc1a2329e141a315a2c3ab6a3cc97e081c4caa32f6ae8c275aa8226c8dbfbe67be29e16e8faffaa57f8cbbf06b97436a9d4d521bd8a497e397dfd24d20c189c5db9b72bf5be1122fa53946bd4f8c9e4c4dfc12281ace477f582ec16764bbf3e2ea308141cdb721515b079391ed13b02f5c8ef31bb5882b2d7d53679bb1c39fcdc629ab54f8676c2162670b94a9a70d4c8f7cdbc2162493978eee6f11f965ffd885bc03d0c3732e08a05e951ec7e04ffec70c426c9da290063128723fb896483953a560554ecfc900af11a876c09e533c62859900f3880695a7719638cf6dcb581937e7cc77a702969cf66dc05933bc0783b0aefeb7c00dfacf61ea358e097d084a4c6380632a8d7bcae06ef8cda91b4f96653d2f25fe3f7df5d4160cd0b0660936a03f6d5ce8a6265ba2c2150a59a1cd8dda059100728898e192d8e3fe6a26fa28357c05c91a0f10c079ae19fc2249155ffdca4b96194ef3beb4bf4b98c200bad49b8a02a890e78f58ce076112d05fbb0e868fc92636f0034e9ed72005e6d9d9016d913709f2e15370343e320cb53166eb6d6d59515268d78b33ac457515ed5613f9efdce95308d54e3d18e6dd634496840b677d4d685a01c578a073600e044be4421b0076fd0e73afcff6aab7e6ef652d9a665ce50193634463a61ffd55c0192311886d59f207234835993213d9833eaec64bcb1904c601f5e8d31ec3bcb15e4b226ca8fb73ea42092ce5946abef3cabf60eafe7bda6a4dec074204b12ed3dfb0bd8360688a434acfa5fcae60a37f569e18ab69ef796da69172842406446a3254b89809336b5433cb404edbdc309d2cc743b0c9c22c0e341de298625eabfef2e9ba6f4c79cdc83e04301d0e52e5b78501bb2a87492d89959278bd4c9bcd2eede04372063e62c300be66e1f005784da13466ffa9daff09a1b14e57b02e58f17f4fef7dbff2568f174c512579ce07644e928b1322f4b81f66e012507e3e43c582960d81eb1efbaf5a70c712899eaea7eafe3ccabec3822c8e7aabf56de28db00a9704089a24b62da9000e394287eb2ae6933fa3f8a132499052243f43872ea8bbd6f06417ec4f6e5cb4169856ba5ab464f5bdcf4a41258ab5c67c699fdd62f3c4e683a16ce8fa55b276a82e34079ee00722e3091c03a569f5aebde9f60830da2a48206bff48b0310c00cc6e593d5ff29670c0f97d68f269621b31f4e103daa6fb1dbc5506c27cd8073b2002e65c4e6509107a3e824b76da1a28d7356caeb8d7790a4cbecced35e3901ecff1a920699de84661414b7b4c86e090c8e5cb43c3cd1a50d61582c15702552613c198711951974410d5690678a3cf091df22c7eeac4305d4e2e5b0b25f90bc40a2fdd7b04a3a62e573ee5f4ea4deb69895a3bccaba95536e4b20184c17183f289b58d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6c07c8db674ad2c22b84da4c6beb0720fe6bb50388aa63eea46055f5994bff975736402d3bb215806a69c7bfe7f2f171814f8c8a00d5ec88300fcf93d07d2f8ea52d6342f63baa2047130cbe240023302e0da50bd7a2a08b5a733c419000e0c6310eeefa30065c89f3b08d3359c9bf24093249a98c845084ef9bf94d7e49e04758b699645e60e9d459ea5254b8be03af13f4feca2f20fe4b3a5d0ec0c4e17833c5ff504952ccdcd96d32b20e25ca32b79c5e3a47ae20589ead6ff46eddb130ccaa6437738dc4093daa61022bb4e5d189b800116c5e3599fdab4777a71201cc37c0e621b48b4b4415b68589c8413dc9b3cb9c68f2927555b402b3658a9253b5b23efe1a9ab91b89283e54e621522773a59b942d1018c900c5471f214c74ddba5abd820f61f95ca3739b7da72255083152e635b3e9c4eb703f7ceaf3e7dafdab641cfea4d19e4a68e1a4c8b4656f67d1daa117af0dc3bb7e01b30f0ae4b23bfac9b6320f9f6c1bf3ffad9d15fe42e10a93d109487ec8e0db7018ecbf60fc92eb7e86fc0ad5b4c8c3d4ad4652c9188fa00b8ae86a09b5e00e6f33240f1fddccced4f2badb56d7c801c912de5a59c2797ad5cc6663c3ad2b43fc0910b52c74913f94cb5a45105f7baffd198e39ced5ddbd8cca803ca1eeedf5585b9df5ee825ed37500ed6cd957d4c46921b780ea4c8e1e170492463b4ada9a286b146bcee1f671d8de404855d91b5238451ce280e6de6f35964bdc3b840a04edc70589e0bacd2f4230f4dd46715e536d39c03d09c0c2b9e64bb65743d40da8706137e5f99deac2262770c46154201dfa054a7e19fe50c6c5a66ac1754adbb9f36b7eb107a36c584ae56739f867030d6d5ad07f988d1960eb1f4487d9284d7986fe2557b9a6312bc104a1f4d4565bc72f770a09f46768fe673c4f72bb67ee8f28b02027461ffb954971d8d3b9b05bc682c41aa43b19c6018bca9ab2f730f33dee6cf57fbc243d18ade95d7c7b71464be7621669caa8025a976a43901eef08b58083934f2122a291ee73be38201b30589f027ef263c1cb3da6c37c721d24039f168684e6163811f409c3d3b76ad32342fdd77df90495ee34b16914357353bebb92d5735f09af04605d854e66d35c1ee047c3d53367ea2a9cb12246c09b4790b3888c56892b0822ff7a4418db626863ba9151bebb4c9d1d9cce2595d10ed1f9518cd2794d1878c045e5e091d04937126b595c06ff720264a3255c9991d8922ac78cbceeafa02020b1cb2953c5a526f87a7d4796ffe357b5672915789fa86b658696940d3e496bb7700b0d159277f9f74f5e748b1e806ce24241103703f105ce13171488c223b036d9524b39badc2d0fe7cd78b6f22eeab10607f534accb125a88541e304f7ffcc029f10cb8ff5b92187bed79c02b2d8cabbcc14777326c6bb68d23d88ef945315caedd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfa9b5e2fb2b05b973e00498eead88343e3d297872f651390487a449f0cb87d37a05ac39c57c116a748e655150f64b63e6905bc70c666a8a5f2af49e0692f90ee1da00648b4cb2046662bb82256528b94cdffcfc6f1d6276403d4dc1d8f06e399174e047248b167a9032c70b1ba18c9148b4468c10ed780cf64871739d15ae58c14a973e05fababcd25d2158e4d26bcb2c9b8c47d597cadef74b4d1b8c6ea57c72546fb27a4fd558650327359df70533824126e58d293e8e39f3266c8134fe69841166f2e50c7e46715c870327862c2ac70936e840bc97e5b69fb15e728afdb2cc04621456ae924e9633cd917904f6c092e2c9c782cf12ee6b2e3c6c09f56bcad7c86fd2dea4d2e5220c5507066da161235372393fdb57742dbb7aa2f0a132b6766147af351bb17901b1465801058d22955c209d40e24c6d78a7d4e1f971716d482bd6a7185983bdd1c9554a9ad4765af3bba288a9baa7efa188e72cb18edad0dd21225b19fdb256d4af4b3883c19da9f1ddb674b29de6b2f99da1f53042fe12bd78621332266ec3a652abbb98411fa4af0dfe56eb087af8bcc6f133fd6a01856a6851c2e1f587a562309ad13eaded51225a3e65335c629ccb2d88a47841e1c320e895ac82dc84474c4536c82dddf915c0f1ac8e64f53b030295816e0428746bac15bb06907f337b0aa057c79748042115d3fc7f4ebd55b3f0f1bc159937489071a57e75f5d3bfd2fb1c95086dec53347b09aa1cf4ac48e7e5ecbe5f626e8e58dc1fb321421a9cf408a13bdb834d242f11720a15122cfd3621c0531e275d955aad77dece73b56f7fe93bf87b9484572d36a07ff15ef0b3d644ae142abd3db551df04f25bee28c65934a1ce6ed5b731b8cdce08be135c1a9af44bedaeaf21a40eecd2c42eef6f40243648e56c1ddc6b9bf6715a6dc6ca05acfd8a23886987fa80d0610a07d24f2481817526b9b18803c7c491b433cb353e924ba26d32e36975ff23ac5c1dae63c2a45dc42cf357f8ed5b93e2812a2336e3639b56195b224d4b0e81cc0f779401870bdb603d26b84300b1f1be30fcc8a1c2fe56c2f12cb920156d425c14218a3d2c100e0d2e22b156d050229943caa2013c77d225baa6ba337a9bbfff6288ee8be952499142edfcb42329f126fcd97f5b02e55dc4e14db8d62e481c4bfc8e93bfa847732ae65a9a61ca6dd2b9af5d2884863fb912fedb4995240a79e21aa0eb6efddcce0aa8c3d5adc24c3740d43867c0f9f1fd47fca7534ce224b1bade2e6b80dff92f597bc925e1dca1fb62e16f9f40c86f9f3884d708085c4e49f00baad9df7502a8baa979eb66006530086fb900e380b07821ad12fbf812685bb9c4a0a6e6fd49330b6282e9f20eefce1e74862e746302630a621cd64df1c7ae06c532a3c1bbddc5dd4dbb519d2f5ac64cda37923ef5eae7fe4f599c81a864c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h80b3f3fb53a5c0c41abecac6b89edd46038590632025815ae4864a670ce011bec0a522f3b84c478262be63baa468f00dfee7debd404ebd059a145ce32291a2af2655f05bd0ee2c8ae506e3bf11ccd6f85936757bba9c3fd86cda909cad979917ba362b33e09b21e3fb4f61c674a45123da5edff7bf1629d0b66cecabf855814becc95d166f5037b9bd4b0925e60c1580355475e5b92905b25652cd3ab49c83191849b32b8dafc052063804b89faa06f5cf24359ab73c87cdf42d252538035b6f218ec13e1a516971921db8e8fac111b3a3d3d1fd47230fdb3ce35822e333ade102297dd75146787db34527c4dfc74c555d4a71812594cf12fddcb4b66c99b12c7647eaa75647c3c0f77872dc7d4661d6ba33ec0d947e722e2864c1438a10820ebb7c82872854eb71f665802ed804ad0293949a38462e904f96d269fba8a55d9c09d80c6f28225f9c150945d47c1eb27240fb3abbe88d9d1b384bac623a73686304d9cfbe20ae6083d317990321fd78876c240a361bd12f4f082ea4eebea7b1b62a9259020350f4dd79f83d7195535ea08135efd7f3c3e1c8c7dd2bde624413a2fc62cb278980eccc2d28eb6e9f51a990d5f6f47260131d5d8929c0328c01e37cd325ee786cb4ee995b911d47ba6c4df26cf8b879aa24d094cb3f1153b5b053d7a4b7dffe748be490162aaeffd0e7627502b278f2d47830993af4e42a4a82b77f137c71a652f18ebd764e5b9cdf53465b0836128bc4cabc4d52a554a83c98a2e959c4a7abd5ac0140b57aa1d93766621bb579b1ac10909051285b95a347299bd0b832e56e81f2cdd775bff51156c398ca256183dba921e8caa0cabb18ae9c9efa9019c7441e6015b54398d71603cd7bf94fa96be71032b01ae0664f53c303cc3f6062531bf64a63e95b62e6e25fe91a66ae74ef606b316fe0f9def98feaa4843793d32f87c00998d9f80ff12ba26d5b86a07dbafc2789305b75677703f566cfecc9f75e67f01f2b41002ef451d2ab3e7ac48d2e974a6cb3929a1700db16fc24bd02bfd955101b4df2ffaed80fe46debcacae5521587bb7dd8a6ad0046b614d4fc8e4ad0150eed780331c7e151e272c31a0087ae2ef374aae8e5adae87f76dba691f5b612d3fa2c429a9d215da3dd49a1a37c74a55c617c5022eef868f79f9631b55836159490ae2ed7142338452728b75d0338f6558c056d22b2bc47aafd3b5aeddd713f8c8c5526eaca33b5b02db71f220212b0df56fe118cd8883ba03b3ce4b2fb2ecfd9695e6fe35ff592ab42d70e3891cceca27a745f05d4c73024330997fcaa2e0932594ac825330fa18aaf37e9ac8838f1f5db15525a26b3e28dd5ab0c688a91a85738c4a3131a5aca271550512b72465d6671802cacd8e3996c5665f1f32b8ee067e1c38196c5583a84b3254a7e7a80a54293d64b31c80ad61ac592a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h72503e4c33a9b55b66f6eb6e86b3093f719a14c0f6548d103b3ad9e8742fd536039bff4ee48bd1fbaa67fa65cfb20010a5fd55293da71960f02457e27c1b137e084840fb49869d5c1472cfd92ac9d816ce85573c992a37381def24cb6cc304332f3331c699a74e4174134f261f381b9f8c1f603176d5e047298da919076c53f1e5d62d7583cfa7ce6c314e72d89a6606e82a8c7a643b8ff69cf0cae7a6732bcc0d192a6b9fa156e013e3a1ae31767a13eec88a4b0b5ac627a250e3a632ecaf1e9b980ea273873360c7e815bf664db52fd9d8aae5ec49900d3b5bae6b317c42ea8a5c9027992c8c45d74e11d6b78b1b95438fc4e630567a88ba849cf08bb4aa9f3fc119e3005a8dd867198c4da6c597d871fd7917b0e9ffa4648cecf7e082bbc449a6d425baa1e73962d6255d28caef7c77b0ccd31031b6dfe52291e5164725396ddaa3597d998dd13dafd74f64acd5d0168b03d3c500c90050bc2411dbc7fa14c6399e6f296223d92cc06781846366b5bb48e65e3647f7b8dfc5f7ca118dee8d917e385c6cdead54fe3a6cbed925e76adca37608e11843fe7a22fc44c849a9169e53a8c85f93c557d7243e9e5fb7e6e1d0e1b54295f0ae0c306715bb99808aea305409d1a0e365690b28b979f3e1c453fd5cf06c24559099d10fdc15ae7f3c55ab89dc6e2f352d62af4a47a7c4e90024d07569b88624e45a2f992db596fffdabb2ba063ba1d70c76d2155bfb3135afbed082cd9be6c4b3a9551d279666b2f2c3817dc0c02f0cb846f4f122351e95c7659b1efde2ba03a951a0b0254028d823846c445c0bf5192832b3764c9cc4e260a71e872aeee6b51913db4a84eade4fe7ea776f9d584e2416bdd274d30481c9f29c7e1ea5c380aa76f6998d23b8f3323d8a0aca106d50d19eaede2ce17ab34d8b3539766def8726d2e257ef471b85a2346242e14d2307f99f26e4dab1cca5e1fadbba240b1aa9477b8d911cc09fb0074fd18609a800eaf4323c096a01dc1a2628c028bb74342dd0104f25afd447cbb9a38024375cc7d8b79a7473fb4b8136bf281fd7453f8f86a6ba498a45b7fbebc29022be3a805f2e453f7ae171cb1d0d8c5b75017a6598b236823b3ca78f5a1e3e3d42ef660f97bc2ce654557cff96e08cc4851fdd08ea21f51dc09625fbb9cd2c7358bc3a216cf6129d2eb0279329d07b0a79cae435ca04005c9ab5f3e99825e1a6c4fecb4a3be1d8b250342b7cdad539b756a5934bc38b2ad31444150d944e0e4abe6a93c8aa7cfc43e886f5992b664327c40b81e313a4da85510cb04a81870e0d8ededa32b1bc300bf94c1cbdf799b9237a94565a8ae4a1bcb2a8532d1524ee8984ccca25d8faf895988788ccd3b25a45fb2a04af9611b654859fda81a5afd1ed8195a1c028d0ac2f0cd0364dc3667efddde97035224808bb2658a1388b52d23f0c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha704d9e072752564720033291ddf250494384e70c31316737322a8a44d43cfab8e3b3d48f546f7cd885cd51d65543b3a8af8b47a8b866f3be038c6e59fe6e055011ad1c6269412cd038a295e5148a0d17a1c32c0882d081202cf31d57a5877153c7be34b4c789e813d96d21e5ca0ecd294d1a18a1f804c4a74e1775b654ca4ae321277846286e6d95bcba90ae6a20c4ef5e86556fc4f6060b42f6d3f918e6cbfeaeff4379d821937b39373b6302d8d39b80d853de78ca19de507ea5ef6b8d27b0fcd853ffca42a563f43447f0970d0f28163486c6ca4bf0f2425eb6a615da4adf8ebae88f99f44854f235beeebb888e068ce0dfc3e2322b866b244244353f275ede828d178271d2dd41d8754dcc36abe8d8a91edfd93144dc054d3ab9d37f413804c45fb4a5df15bac96c43f9078ef655950bd898733e4f4a1223168695e4e8f78a4ccff8b5ce5ee28a9f737f1db7445b6f4e3211019255fcf97452799f70502f823add1051135cb4d8a7cee0d5be5fad516d120211a2c2b1e50a081cb2b85f6d3b6b615ef11035fee5faba698861d4b0310994552d809158c231036dd728bf8c591779ec5b9cedf770e81829c50d8644fa76986a6e8a39697cffb39589638410181c89666c34efa3f9493382e9658209987e4b7a5490db1dc076b782bd0d03e0476a808ba037277ab552ac145d4a26b12b8f979cb557f579e1d85a04f6ea77d95cf875ec5915097de0736d678f471e900802716bc87ab9e9f67ceb9f90d357f99540a39980bafbccf6617ca38d7206372e105ce99868e9fccca144d5bf8e2a21b8496aaf34f9345b85c29b5073d5bbeee9bbbf0e94cb2cd870f85d1ae5064c891cf8e4919bed300555de725515e9473705e2117044d762b39db9a52d774adfa23a99f886bac46ed5fad68d43601113f6575160ecc2266a5e30c47426c67e04f02cfe8f3b09b9e169d0a5d6e9379b2cbc078eaa67ca76bb879bc94fed6f23adef5cb9f1a92e30545afe1f31b447fafe98c7e67820c6d412a53e8bd2bdd02b00ff3c63413a35267cf79afd88fd62bf0b570e8f1ce409c321b4ca992250e657fc3fd54ece23b97fa9b4c5d9fa7500b12b974d02b04315e5aa1acf2e8f5d3c3d23adc7cc4efd577a835b6a90e5604b7dfb10bb82745b8ecef74c5858f47b86da1e682b09bd47df7318aa9193078f8410368bbabec10736a863714a74338c02b193bc7e0802b67de386659a0e1b3d21c74ed63176163dec848db55f10af3e85d85807053b6e0f851bdf37772018586ff073609d376b0111397d632165b31077848e210e59bc62818a343a893a3e249f3c128e3e6733a9ca0c374af1ac6c40d0631ca5c63d3742801bb54d4ab3aadd145e71989317cfb1e65bc5e96801792a19f1db509763fd4e4dfa40c5e9902ffe3b17a944ca85eba8bd76dfd60b50f35012236e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5d40bafa6fdfc2e39c79035b654cffca4a88b87e90ba9315305e0fdb55c0faa404200764d889b956758e6d3cef5b7c4922c87c8d2414f195730d7396760b1488d8a204567bc00365f8d8960f20703d5ae31e4549f37073a2de0536979347124eda5b19bc2eced802269c3795dbf27314d6c19c7e0bb3a7ac72ad5680b803794da0a5ad7b5111489cc8ce099462d8989925b3f9901ce72a9615f020d6a1cc83bd4d3d80a95cc3e1438b2c57db6e584283381ce273f047a6aecfb45a022752c909e15765e915be600ac2f1a75b7c9d0460b485e2b331afe9cbef383b781198fde6d2359946d59593aa485c4859b0feea88143b158df47877753f1e642f205621fbfdb27d7dd87fae64ea6697badb9a7f50ba12de87df5c8f19362fea07cdc46250a510b4a578f1acf0d13d5bcb1c1cf5acf1b59730bf5b4f54ee80e45dcf2fde33583d0f4577426b86a4b6a30ed6ce99105b97233ff485470ef1804da939c59abc51364e148783bb7062a720ba180fda3e211a1cf17d91546a60d3dadd53e4574c1509f8b0ea77291465955bcd3699c1ec0643d63777f50e113d7db6bbac83a6655ca71f953977659891e55553a4311e92ef9d46e680bbfcc29c32932da48561c1fe4d406477aeea29c9ef2b4cb3b1527e98f056fbc82570bc4d2ca85cb5c596008dd91334ba21103de9455b711ba5c7ecffd816bda8aafe2101e2b7dded2546cfc176865a0d319b3a1e1cbac93cb8a9015cdd2c1715352c5f8f688f0aa8bb6fd78d9c339ef2dc5ca9df378e11d0860623a779a861de793c1f5a40b9f72a9b7dedd0499d048f442c31b6d0fd0c41fb5903b55aaf4f2cf04eb101599d244219b35279b932eb49e172434118d901d35002987767862d20bd5720df489721ac61c6c6528159bd3b0cfe5fa62e1ae2da7b20cceee1a9e0585a11e9a75be94edb3e9ac0606410c84736d8630d89236113284f5f15db11ec74ac1da062e3ac4dfba42739708dc9dbd616a71bd323234df26312ab15748ead99734f035d8fbf33e4abab1c8e10caef6d19a9dbcdcf2ee60b27f5425b21a8e3b1f62826976ab10c12f38434330afc434851ca8f653667f9e74f61a22121b6ba036bdd90d7ff6818537c53cd71658b7a57313b5463e91ce05417b665b307d8c2d58f2074cffa8fc075b4582fe02551f14ab78df8dd243a5e93ba119d505538b86463549e7513bfb265ff627a09cb58087a2d0aa16df8b6bb3959777106805d9278f1f1728d981970c5c2c7a609600e25718ed106d957791d6e96afb76d89f36e4ceb41ba1457906ecbe09f8592ff57d495f4d22436973c654f866d025a6ead0dce49b8a8c9097ad2eb3bd4668ea1050b14a3623b6a02f418b0e4286ed6cf5a8631104d775e15e780aa2de5c495ba5566b7dba1d9eb4fe9183e1761a3176c5b42a7261b8cb98e4b4db84e9f5f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h341708ca41c9e6fd41c7dc42e16e47edd19ffeb1c0f56af947c5302d4dd3e5be42b6ac2f657543f030c2e224747b36bfff11c46905441a09691b31b9d6c3516e190fde1797fe4259e7e9042bee966bd60dac25df7a599dc0e11477c974402ebd1f5264fd5f08b9b1e9435f86720cee7682f5cb9adb272995bc22e3d9bc30685a6dcc17b1bdc26e5b00ec0605767fcb26add85d86627e01f6e45f4321b9c440470d41c242b4d6e883d8000a4c985f6e5ff8a8351dee55618592cd3d05424c8eee520b708b10deab504445acde42885ae78147f6eeb5f9e391a8148043415a68dd6c337f13e579bc0344881b3f0e3333c7fbce12c0df26829cc919caadf1daf8bba33e81c597108cb6a56cbd1584b7915806b80ccb95df3eb71558f1ced8001017213aeec6244a04098466071e0eba96d6fc1f0b99c5668833411a39131f61ef5bab9768d3c6cba1b45fd87d8fca011b7df03a2392633ddea36ac7d98fef637666232804ba2216572c4531d8b04a7ec6abfe5883151a1641b402b07d40d9c679a7eb812b807e43de1e8f0cac7fdba44a3c3ba6949bdb5126ad93bff5253fd7daee6975488e1bac2d796378fe0a5df101304e07da79eae874f5294923d201a96638ee885cb357488ec42ac188d610f33fcd4b9a37f906dd52d8872e45ef2e5982e90c31cbc35fd109b4507a116901e33e49fb19c52c2f022272544cca72555adcc8e7e15932e860c873f1ac4f110040dd163f2ad6e449b2f35570a5b84680d68bc577bb3a1a114893d4c8bec7c076cbdbfb4f4207d8764cf0994883d004a4d05593559f9e2894a7400ad13907bc876d2865f330a2b7af88d54215e18dda5c016c75c0737cefd511780a90bc2f77c1122d11aaad0adae56171bb4ec870cb67ca30334ebd054a9e6cffb9bd22ac14df2151af6ce35b956dc77456de365356f1b99c227248124074df7b0c023a7ce9615529dcf984d9ca434d0ec57e901723cbce077b870a1d61b24832dfc3f83fda1389b5b3daad7490354b005830f4d787b7346de631a18217024e14eacf498a0bd39f2b8975df40525ca10272d70a2abd1bf1098eced9d12abfd592d65abfadeed6baff8a53030433a0c886f4d5811ed34598f6dfa223420223e4266a7d6403947e2d351aead1fb1982ceb8ad40b3f6967799fcca19da0ff8886ae76e779d2e36aa50ce3b16330215b0c25c2888d4415bd1deb4d7efbe1987a41e52c3b0f548b541b1f98c2b08ec32562ae0c35d44546d015a2ea3971c8b65bf1bba1ef3ac0a4602f865a00576fc24b9f5adf4c796969d50ae95475ca77902df322dc55714f459e6ffd39a6373fe1bc8af23e92f73583c01a0a0e26c14861d7ba42b87bfdbcf86ede6ba0897e17c86006018ec42422f729d486660f539781b65fb31854087d93ce9fe59b3fc1e97bfacdf387808a57e3fa4ec5dd8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h96b552918a99eb05f137d62893327d33fc84759362d5241a3ec8ecec5fd2f3941487b9afce901db86e26112abbda944b6b41371f22acc49cb7783d57db489734ee0e8cbb1be483ddc96588071e7fb66330fede91817efec052551be0ff2b05b6478e94f84c4e0e1eeef14b17f00fcefa04cda7f2792b5a4e9b2fcab019dad10ed80d6a7fda43519b132cc22ba0ea00b617bd80acbe57de545bbf8426fd7f32c4b0a3e008ec39fac5395842770b19c19dc51963af773380e4eb598dd1252d90515422e0978a86b5b71a926d6941c31f214b125b0f1ee55f2e1f3c41196b5b3163b772acfba5a0aeb94852ad5e3df92ccee33fbb5c99798f7469cc1e0d5738aa573c645168c1022b451d9df6c6e74f489d89f379663e9b7ed5bc730e66883cc30338f042374d8f9e6473ea76445d839c22c48200673def85c23a67fe719b12fddc1458aba9e64c0b7438b6129f813973108f33691d46261a7f946572e20740a3d04d313c060c020024b1a2d27213c8b3e9e0649291c542c19031754ea707f2b9e9beb4683a9fa177a0a7e353de727d0825032e45bae40fddac380f88b7341497a0e57a1fb7479bfafd92338964b1537097cbeca115f166f6af05b006beeaff9520ed84d23790c42b091b684e2beeb22eacb303664b814054e2bf7139a284b531e0cbd6f84bd5832cd8fc496d035e641f45479e1c1954fc7342d7a292bf245add16a6027beceff23930ffabd414fd7ea5c6ef3f2d40e48d925f766c156effd66200296cd37d3311b62be8232898b698c02416fccf2e7ba6f8f1058d8ddb18849a422ca8a23a27974f7cd1321f78ddae5626a7ea901fe12eee27efc1d82e2e84cbade45b1b4caa9f4ef7def0355ae8da9feafb3ec761bec04ccfccdbed3102c1cf6b1a90545dd86de5bbd034252d27089ed905c660f6381c618c29eed8aa0fab87c7fc1e3fdfe84a3666908ff2360998439e8028f3d493ac6420e1c381ed26bc13bd682793d73488c24b4b589c26d4285fd5f17c820db0f06ac3060543379c2104526b8ab31c899393e6fbb1f9674ce0059c245278159c017548fbd0bab00c08a4e099cb3c119b7f27c4742a4cde0cb91cabf17042b2402b1093825e95296007433be7b043eff8d5a4a37e95e13167666adb8fc31af88fbb073c30b2bb9cd24d696b8a06d7e17081d95a6d6a3dd4efbe4bde1fbf5c6b35bd35ba80082b4ac8854d14dc92c01c770b55c04889bbe93fef2058eb84f30eb8f78ff94796e2ab4d183bb7c3bf4d3de025d4985d2e2218d31d80554f98fbcc25b744a126e5d2c7a4476ba897431485911f06a1ed557d337da07391d09e2129f9ea58efcf0ea9901ba3b407b4449e5d16807338008e24b08079ef7f21774fc06d98753ef8ef0f2245ae8230cdf488df31062c37acd2e116206c449588fa018df493b13e03f8c9b46c38978c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8dbfd113a9970aab4030e942f6772b817ef37c9137029320102b13ecadeb79ba3794f9db20c2e1038182b43f31660356f80a91e9932a1f76144baa61897eb34ed785aa48f7222fdcfde95dbed0f7079953396b720277495f231ad2e79ec53cea2b82afb77aa7413ce32b6f7b3070bcdec47daafaeff7ac51392af3c3f25939e44cb765ba6803a5c54d21e94e1187d5c8786a90cf0299124dff70c83a86bae9e1020e0eaa4de7f6d6f9247c4b9aeb224b7f80814afef5f775e25971396298968cc0e5b57205021975d3449fda905ed703a1dc5ac5e31fb0b8d5ce9615536c80ead9a27fdcaccc76085cd6e37e8b4504540f1e316d885669f36f27f086e1f93e025d39e49dc3050e4ff05c9a7aff55ea22602b4dd45806fefe6fd50a08fc6633b9aa228638ea3d2d38ff921b0f3c700b21cda58e1adc27ba479009af4bf81424adeaa857b8729ddd7ce9deaecae78e6066f0b609f06a2d93708fca6fe35e276bfba26f4dc7fa2405b0c64b1b18977716088ddf1c8735ade7e0b3e6013085832c13ec2956daa28a4ef015773efd560bdc19984bf62559000c7102149d3b42d89badad0f0670e02a94ae9282c3caa6974332ce5b66976a7b6f8f45cf6ed62355ba3813d9a08eaa687ca5f83dd01a00f4c27f444b9d5cd8864a82d24573a59c9bd920ec9be88d8c80bdeba2b7529291781a1cd5a5b4b34b4ec1cdcc6b2905ce554224c166cfe78dc44b6f0bd617a091f75735e0bb3d024c30603ce7805b7731dafa4857b4eec56541cdeeee19f6d105e2e0048f7c489beea53dd383931f27afa47998ade4ee30eb31f694835b232ec4331925fd34f375e23ad92f00b4ac0f9d044d87da852e741fd969bf18338c1b367bf37e1b5a468573143521ece9224d4ac2d0fe3badc9ba9920d50295de5c0f20ad0318aa7822b16ca792568bbec52fdb0047a2be2c829c95e89b3b8dbe16f237c1aca7a4b2c79399794fff04004ee64cddd4604f03cde1b9197783658d16d42f5922b074c20007aa9f02022f5c8a99e3399857eb0c3b68e044bc0b8dbb0fa2b6c31a16f0bff1ad20af6fbba590b28bfc82b45c3e71977452a24da589903ce622fbab52078d0e26eaabe5f4999dc32d27f27419c0059f53832391ce030b4443d1e1c02068ec2b10ddb282d38feeb7a564a07871260a16458d10f2a5d39bdd19a690fac785ed022376f2cc1553b3c7373616918aca5ea3335612333a665e0191ffd1df7ed836322ecb8a93b2c83845a35cbd6e07bfe674b0d4ed8abc3963b50253546b1baba4a8075c807c618855c06b879f0956a1888ebac1fa6d180e07218ded50d9b35ea8bd6f19f90b077bd58c6c6075572aaf0a9d368ed968e2914ece3dbffebe284099f11015ebd8f71a6f0509e9797584db6df7669e23b4a5f9bbafb24474e9bd4bbe5440e2771c9682b5b57c772997d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h307f237fb11abd2c6dd00b178b3cfdeb7491155d6adb87193bf143a1f3ac2421e4b9e0cd4fb069c105dc4ae57446a490e88f708a75e1a9388b614dec8f5d5c0f4a334f438a776b33c6d2e859f941cec00e931a1d1dc7e33881ca16d6251985667b4ad59aecfa8d22ff5482ac2e3bfbd1b67bf49e393de6361e33bde84a96e5b333814f46c4491aca65b39d86698074f1afc0ce8fb7607c37a9ca10aa8d3089da4893793aa72ad09b526d09ecd456f354f3e7eeb1456c7042b4eed517e0f0a363ce463997c5cfde2d463cd49d6b9ebe75c2dee64c9d8a6585007be2893d3be710c1ba0d8c84c12cfc64b24aa6b48a068f83886652d11b179647d6074144e09d4b4fd6f6bedf2838d7e8c4ad75f8921458c18c5850bfe71cbd544efad9dd5c1a0a79c4ac1f3f84439faa4feb323907748f503967d1fc632da153679129ad31151a16776ed6c103a29f761d3df795426d52558a8dcd16ea2b4862681870f22f5e5e4541bf503c31b3b69ec049d83d22b3c60f4f46fbad90d44b281b56720627264af3d931658aee12cd7c56d7a08e7e769992bce06cbfaf8d1c8ab08f1da79e832d75c44e0f31828a9c2acb6e10f9f906055087a12e88e98b3d0915c7324424e1b60a95a7eb1da8e2bf199871a84fc05322ff93c764d59107945aac58b214888e80a37288e748e32a3fbb5dea570556357381a5843a00a4edbcea38ae75f6f822852c767b263c2c555f6f9e4d4d6dc91c84fc41fffe67f0805ee9c0c0312e5f638693c220235959ebb2285bbc67363082c00ba5e563a217c8c97e07ec7d594f3172c64f9f5a4841a18e923b04bf710b2abf2702b86a8212a7da82ab3f73d5790fe3989355c26d79b28b152b75f658807a475df3f2a4998d90955a0831e45ca62f299e1df5f512ce3c20c0b8e84f05cd5b3078236b0331962480e2690b1dcee342f8a0a7a5a9d68abe51a0de6cc0eb2869c7fe37f34ac687d95fb9738ec917aa2c8ebca23ab92a3781a663451e147df41c298b3ae89b59edaff8648c8fcfff88b1a4c202ddbfa057ab1c6e0582f66845f1f85995344b5386668a1c941b6d9f5794bbbc6ae756410148ae63a5aa85e3c0eccb0872dad3bbae5182e94126a8300894e27e528b652ccc03ef9cde0a2a4773a0e7ed405de5e001e8ff1dc8d67689d9866b65d693cb5b87a392a0f6fffc0192e60401ff4700e423f553ced2828f8dad9b1f6d9cdea667dd3f61e1d5ec839e8871b4c73d79ac38b6221267fc4c812f1e12a27397be4dfb8a54124e36dc3c290329dbd9f689a8ad2a83558aa8af2138ea4313f1b31c8c0e058fa266350ad2fca50edff7abbbd8402839c1d8b2872fbf88c14e502c5df956b98ead81339ee952236922af9c9e37e6de1d9c507c31282f508bb726da9a01010f1b5eed33047cbb141ece01baa9be4396f880446de4a697b624cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he8e702cbbd662a698ff302bc1b13ccee2493c910a29f4c20866a03fa55c6892f3eb625f810f19e0984a47eda0a88c4edf1ec9a1341a2b1485ccb673e29dc8882200364128f6c1b3558f5177aafc8f5f106e48efd64fa35195e1310fcafd4ea0b63dcc0a12d67665936d5f89012cb25c8c8c66b3ac46630f53388ff88a24f2eb62138ce52c809fa9eaacb970a47f8f4e73ed6302a360fce99640e8e81efd70994b14d627610f96b434ffc0f0dd89713190257e6d4f08e32f093f522b758c684ebaf1741e61052d3b6ca598c3c76223b02940164898f6605192c616d0a0e1a18205f0f5c04837961312f60ffeb5238104115b5159ae468c8dbfadff175f50ff81eb6d15f27eb1ee8cd1a43cf6fac7f397f27ce301220cf2c07707c0db26f35317ae4d2f97f6168df22b0745babb2e0ee4524e87e2e101e86e5beeac9d54cc647e256330cf11b5205f102f5ddf6e3c79f2c5ce33f300882d7ff2eb937197f7a0684c6700dffd7ae66f7c9180e1e4e859c3143b6f4e2d747bf921364ed2a400dede692ca7a38097952285338d1b3d57076838673ba5d5c06fada4b1f9a0e990f064f52c6b3adf51a40c8329ca9cb4a5ffe608cccda044908d42321b81ac994b0159d86564ab900a250638bbeda1a572e8bd9ed395f8d274392fbb90824deab6f68515a17ab7d99b9c5bf7cf3c1c867d0654c32a8f6a7a7fcad374908a779e3b713e0eb676a9c081a9153ca80c139038ba0807879b87a24dadc7852056b0e65d3110525683cfc008cf8130d77a41d4bddbda6cc431f57b306a52b550ca4be7a779b021f2f0e4d36ba7bc0bf9a7a1581c1ae41842800ab3b3bed003924d84209f10c26c21c718be453e238fd39cc54a3c0041bae927daa23acfeff9fd527ed85c149a110812d4b5e78eb9b7d3e6ec3c42914c8cd1d4acdd9d5212e5131af7fe7df442cddfaa0e747bf3d371314eaeb846c0d04a19e833111b55f441a3cad0e8b70f9399905d94b866c601843dc18ad8169ece02f3b8cd4b1ae4aead5ceed0164ff7a07ebef35bfc3dde567431dbecd2f04ce288452f1a6d065d0d3789ed0f3fa0dfc69bae075f97bd0f4d8ff5d2deb904c5f2ce1ccd4c79e28752397994d4f43778e032bb7f136b94ed89b9717ec7dd404a3fb0398d5993f5f7d028eafe809245af214a578d85305c1ffd4c35b9c0cf59841324c0099e7d3284800fda815ab845db81a43690ed06070fa712c8e1995ef041a0521e64c70cd44fcb544f2591185261fff3b477ff257eafd6d4f4fc0352c1900cf997c93e37ce8f2fd3066429ab308b069ed086f1dd911542c21e8965bdb3c0c283c12b981897ba1f55c6de872e6c171a67c9669d96c8e920a7fdccdf44c2298e45b684e40d72063cea175fea3bb61c28f975380657c921d3c000e9cff0d5b51a92f2e3f9fb3b05768db46c0c41418a35c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h918b1eb892304c4c4e0e9b93f8b96f90046fcc0c1817d195172c1180c4f60139a65322a41a872655eda3d7c18b8c8d266df16d48c1a5fad4fbeb0e4de9c85cff39848d556572f87a3da60fc79df46cd72a3cc762b95fb177d046e207913c22779e513ac291a5d70f3ffaf67903832f3a489b89714ea7d75b6d0c81e5213572d82627a958b094ecddf547be701c394fb377992fcfdf5cd035b171b8af2e4ece84365fb47e80d55787b28aea761b71903dd75e22178d6ce6b81d9c587bdf90e6cb85e3b7e8b20b7187212d1231046aa3df05a6ae7272f3f533631f3c31bdef45b043bd2c13f125de03813880198d5d581217e6d270e8a79303f3dfdfa4e6a4596d2fb780b39e49a20dcd2145b3252a10e78771537336e62049cbb50b886f68678610eb52011407427ad84f64ed8eeef8c0e02eef544dc7a59b150d2313763b45a99a79a66c5a323d7059653a40b776e045b1b351de77e3f44cd9a241750c300c51c9cb1e519e9d1e3795cb710fbecca1fb48066397861d23bf6dc3a0218af249094acbb3d9c8a01d5e7dbafc20bc865c73f987c3869da1f08608c66424baddcc7192110efd6151d2a652f1ee9d4d30473a209240db3b99a4a6af1e069de75b9e5e5f3f184079e53685b7954f197ac39eec2f73197c4977602a5c6af5e33b20366eb209feeadba81a0c97733e4577e0f151de3b6293f219c664671946d9cb3dfbdd356ac290b43e1b9fba3e204e16574142cfe960e9edd5452bcea3d561431ff10cf83138da2e732fffbcfde9f6470064845c1d8e5921181b5b502e480f13ae2d29f440318932149d5c9510c1406782d48e167a6dcc27737a8e5c7c7f9b21c78dd730fd3e7103dce6e89047fdb13ea0d4d71c946ffc16bf599200314130fcecb7061e8da4d8558ab9876afd957dc687db5c06609e1c1d7f0d0fe4d56dda7d809f1eefcc11b4506026ad933cbdb4ca3099f68461788b22b0bd20bba8022207aff7d49562bb7abd878ce92af2a31ddf8297fd4b874a1f29dc3877f3568b15740591db36f34c82535658c3d85a6034307bf96183d7bad7038b1cc83fa6b32da25bf7c5ef5c370c802701ced84edda8354cbdd33a2f6765fdd21fb93b826d0dc4084506e488cf95211c645915515e3262c7d70f791db4a8ba5a128a13b9cb0adf5d0ffa8a36ac73562dea5d37cd31304680b1bf614eefe1d6044bd610a0089a5df3ad8a6e3263e9b171f0f442521c17b2349a31df9c507e7c46892752861deaef006e284993357fed0eea626e8b852393b0900f548d7d705e728b9410012928656119e323c86b1100ca8ab9341a9fa33f9774c9d23c3435aefc46d35119197f0131d3d09ac4eb3f2cb2fc8ee8b700e66462e848161507b7a1eedc1323c6da39fe1b1bc8710bbeeed56b2bfd03b619ae9f52d4eced4be37a2a1a9e303f4e535aaa74149b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcc28f925d8776c53e639a8dc505691bef8f1aaa0305fefa000df0d8094ae508c3636a335bccf7efe70c197392a9118a671e64744870c87fb109aed1b60a50bfa30e6142a7a74f2e1eff3cb5bec7912a2bb7a35ec438c8e1bf7bce84cb179b65c6c228f4777bd6494d6e7e7826b3ecf369f351803b2ef2c732122678468749ec1e6a14141350d7da35cb9b28bffa2bb221a111cf901ab5388119e57dd62c6fee8869debfe1a9cf1b2f7281ca2ec34cb1a81c1ab8c26c86b54e1f9e1eb745ad4a645608350afa82a56dbbd5a4fc68cb71011b501cdf2c620ba3bd92b1b1dbbd210634ad04ed325d254d3e8bf35a6affa796278f52e8cdf8696d1482711ab6bd24bc6519679ae8006a80ae8152f62d7ef1a3fec0769b3a4c86d7cff87e78f221d482cfdc23ddf38a9852619a9cab737d8ae4fe9d1b9ef4216d5ad3f7b47862786f55bed10b3d4a6d82e2ec9d1e9839388b5f8bfaf0af92c5794c0251019fcc8d27f1908bee7ec37968bc4100917710cb5999f6e20699f45ea7ee4ab1f21ebfb7345212bf206f1e363ef0f061965a4a91f1e4922cc061ee0898fe6002ff67224438df78c5a4e8fcb45c55dc8bc0aeb24d6e7cf7f8f5c820ab7502b2ef8a9dcbf43e0ccf0753a3aa78683208485b90030cf4ce18ce33b38282e75bfe133fea76bde00619be8561eb1aa306caf5d88f6c098e3c28aa74dca356c42ec815b366be84e6f149d0975dea0fc1453bb35b26996758e6225c24350b023ab67993743d86c8acb97d5f814cff3b662da6844d06bad17926d9e900688130708a611687afff869a31be55a718b00574fdb84372f45f46ffdf3c3f884ba3ed6631ed2807c7a78db474decd23965a99aa546dfded4cfc61a646f01bacd16a5971cb26da0b2397756b0dd6a5480722bea40a426e19fed03e90f2b717a1846192b0a357f9d45aac092b1ebe4fc604ffeb5125e3ce4d573e68732be233823732d22e573a42c3228145ece27ca46ab2c89c6ece3024c3b26d916bbaed63b9e4c0b6122f5cd997c94fdd87728c34779bc94ba91d454705344c25396a88699eaa92a129c4f620870ac4ac97d3159a6df4e51635c72fef4bdf8fe7cd9e1ea78bd066959c77ef39e55403c03d3eeef644b1b61132b6cb657503a22157bef4dfd5d5c775bdee4957a3fbe587761e7b3ccefcdcc4f2c2eb7a4de6edf232d6724cce92724ed1b1b52e97ff1276fa1d512a83bf8e6533ee466340933c1ae96d527f570af48757e9b38dd220d5cf38e672928755d7151d8d3f97dc4ac59f150d0a1f9027e0c3d15b2bdba4abfabc741d12f8ecb1c840af183aff41c51483e11fbf1d7443422b3d2aca5c81f8949569cac1344b031789b7786a228fccaa8ef48ffb719de848ca4c47299f736044ef0207aa642385dfda03e30c15b7b1f9f3907d57caf0091b85670f3c48aaa1adc9388;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9161f065ac1ef927729c32738efa76575a843db38fbd1b0fb9a841464f70757ad8642a3601a4a35d1a146d4e2e58728babb6d322a18ed1aec92a257075b4365eaccb1b42467458747e4ca51bb7251f3057c3160a31f7bae0f3b8fae3297e7c9fbc6f63c19758be2754fdffb35be3d2f52b6c51fdf167520d3daf9173eda5120748159dd69d25e6000af0f6f0beeaa72dfb539f223fc4a2c0e1b3a67e4fc779d8996754623a616a53c21bb86fa617743c43e79ed18a99798e28ce668f7d82e4af6e38e020df6c13731d550978752e66ed036cca9b60281defadc4f8a11df4dec237542a14b522ce2b78ca664991cea107f661e83bf3c37694d7a307f95e3bbc79aa13e54954512ebb6d18996496b9dd818391d85b8afd4cdc31456a882f9b8e7f6bea21e6fa80309ae61bded308f73d85c882480c53275718c0ba78891b7aa3b1c27ea2332ab1beba1b534609ad8cecf0399298c762277943d8085d498a03384b62213b10fc4ca9258a4c5c36eb312b1b8d2c25ccfbfcaf07eb34754631cc1a639ca3389471c1462bc7e848bfb74c53dac0407b328c0fa56866a7b471da640752cf4d94f04a933b87da9a1c5bd2a6612cde80a477f82b0348e9b5e8d9ca1b01d1841a880e023c259efb5892e26b604f3b52bee3ea999eebaffb5d5fedaed63eb342fb13468a5ac4087a3ada80edf51caa2101070ad308a627fc248e546b424e69aff593c8ac4cf12aeacd4f726c702c04dcf9b99a843c8447b17464a6076e017382a6b29a81e974f4c48942c6450226c3933582436c0eb4ff3d4fd38408589b3339d08f7b5169c40c1f9630395fcb4b4d25dabc9d6f59e86cf8ad5b5a791fa3cd30e81c9b25d8f6a47fdb67b5095890d2ce269a0749893ec49241039f97fa3da991c1667f32c45e0d69a28070c5f2e1b49e7e05a07abb4e242160292748fc0fbddcf2af8905a88b837ed72f1646893bb2107e9eca4253e6fab9cb4ff9783f88ed943e9caa15fc704f571eb5609c0cb2ac1a454571d0a178c484f749af171dfa5f0c9ca859952007ac4362b22520679de78ac02a2dc279bf2a7635fd74c90cc2f02639baf8ec7a0629a83fe50ce227d61b73126396864e565008a38045f1d50ff33711cdd3b64c035f62ce75aafe20a403834db37604f6b45319bcf99474bbc94be4f6b30b43f746acf2dda9f5c4ef9730b766ccb080038f0e8d27c9bd26350ce634022d980190fd73e9476c68588905da42d38cc1641af15d019b3e109e5f936b069b2282decd96a06a60dd77eebfe621f9934374dd924c46a3dc100249c3d0061b8198c446c346d0808e6d2a70782233633d304d0f20a3f724db6b4bc988191999c60100afdd9e715eecbe3a9fe2bbb00fc7442f0aa7ce339c3e9a57177905f082e95fd0eec7dee95ec1c1c3a567b716162e571b9a2ddae27dec2edd65bc6850;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52ca129fec83fb3df15eb3faad3f4ca32c6507f4ee4da2758706b8dd8787157b7f063c81159475073053b2936085891909058c95ec3753480b8a97954f340805f5d1c4b33a5c67e0d84f460927362f474ed3c6ff24c235b148d9a0bccd64c5d301301fff3352ab3a8d3eb32db386a4d6a3321e0ac7c7871167d7f142bdd4e16281d49b9509d92f211168c290dc1c1b0963286e73c6009969345da0dbcfe2aa03a571799c2f2d2704950ffa7d18f78dbcc665c473730568f37a4ee2ca1f6e7a87be8e8c1dfb1ea21c8ef63e0340f63b7e06c473a3884691db85f8b5efb75cd8dfed8d44a862f492e0878edb7442e4aa46fe8bd46be7f85978bc19be30cb806db743a1f8c36704b3d8a0910112a5f08c4c35e45207829cedebccf02993eab9ca33372898030955500203f14de1f10bbb907b19d2db8f99a2fdcfdfed202f108566a7fd3c011a81ba6d8209a300ad3b1841aede1ddf634a85fd01fb1041bef655253e158bfdd61c67637d5f4d1c7bd252e78a67ff015a280b1717f73818f64f238692457646d27c6a9c7df3eb99f2623c668f8cce2c34b3ba40209cabebb93886ebad64d770ef993413cdbbe25bf4493716717f1f30bc0a821b5d82a054cfbfe36b64befc84d1394575276a857c5bd44c3c0d0bb4f1547eda699f29d678460c650bb51f2889344693ed86b2e89879b823407156c81867b9e328769f646394ba7b175b07cfee8bb973bace9fa38e149794a5353f90f7d56277f9d010d91828af66020bbb472047fae544ef785ce3ce10fea5c20ebbb4b15683f5394ac8934371669c98bdbd0b959ebd0929d4db81c5cd6274f09802ebf197e0bcfd030fa9d123bfd1dd9c763d294314fbdc0d908d860a4a09b47b299d2e90f9b7be27cdd8b6b6949746e48497a031d2dbbc1b922c11b5847b3696008ba0e060eb02a391e6470f1c61930c0dbc789809d2ef550f870e5398a1e18a75083f2683641464537dffd3b4d534c2aae55f772c3daf38ad7dffe1d4ae224f33bffb11497ec37a03af1731b8d8631099044007ae44a169e2e9b003f245c82ab256276572896a67101ff4b5fbd77c129f3a19fe1a355a53d247e3a9cd46a3c49da9628e24b490acf248c5870c6513c9675c14f26bb7a26f46c76c76cd891e025e3a5d922965bac1761e301a1634be46632ac38fdca0c629553d38d0864875447f3ad3d0be664e350796edebbf202e64f782fdd585061c5cebdd8a53b411ac447936863a554578e3a845cbf9b05bb3788be670a062402fd1fbfe6648293b3803df2e25add4efce3208ba05bd759ac67b99def27e1207e198764d0bd6cff7c3c755de93883ec7cc9b7dd8c70093e34270c0a6bb880db56ae427b68d84198531d26f75106101525216b33997a931f0c8d230261260da41d26433a942d2a54f6f9137debdcd3a52700e5d33ba6be42;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6ccd88ff2c73a4076d1f215da54e726f13ea78a00f074cd6b2dad29044c8c1081aa75c07eed1ccafbcd38b7058d272be707cfa0b8e9dd402e5227e26a9424d02e0ec2f8f795b87438655625af23a9ff9d1b49d0787646b26ecb46fa8a6a4d928d79c8553478edcb555d58817c26277b2c4bf162daa848bcdbee84e19446af8b1e6e9c8909fea62b851b00139a15ff01d80c441277ddab4b2233f8cdf1c22b808fb9fe32203af995f9119a2431dc8b9ad2c777f344615c5c1f3af7599118c182292da89bacb1fef126549779d8a41e31f5dd8b0215925a8fb2928dfa3cd40e1441b312d26278023a68cc37277654df36fa85dbbb1eabfe85f6796f5e918482b03408fbbadeef656b33a497fc7e3c4fde9c2976678713490ff4a53f71f0dd00be4835aaea24bdc16e3f6a48f0cd47572d618b962a6dda3c09480b2808876e9b08a442451c60f03772503be97daacf38b601d800b20865bd8c694b86924c06c9775c020a87b9213a95474de134f6011de47188cd9634e4995e16c61af1d2301f09434d312113be759eefd8455a6b4073c46344c145ef7cf8d57fa09bc86bc4a3b9985897de3c699fdb459dec8594a66f895662fe0428e8e3f6e4d5fb2f79e35a1258cf7a506594a6f418b306b674a9b692a007f602f3ab9b42dfe1dabdc34e3c8f9fe9d3e303e9c2675c721dd0d10d344c1168586cf91b6ac6a19e9c4edda421dc067ae8f723085a2954f727c752825510e1cdb6341edbb75c3a98181d6b5ea7e498c130302d53d255a2cdc70125498ff59d9696421cc4b3d1d912d7c065bf16685e6d9a0dd68486e8b0d7e085325edf3a9926f58de01d7862d1220fabe9116ce57e1f0a4af5277133f9d45e1ca3ba2ab9704972427d4b480546757c82b2f072a53e47e10732e82b2575202be462fda4a85a57752fd5a8abcd46c180f57c9c118074cea783416080e174c4278ac0e02721aaad2d57cd29d3e7bc261d82591012280a5702450e6704a86ecefb69290176db6ab036fae55374c59250f77390c26476824b4522e452b6c6310e78eb1001f733bf99dc99f79b42212b77671f27421297009985aa0c8da6aeac636b3485883c7c3a97d2b1c47fec371be1e920fd3f5d1d1e179163b3cd0713535f6b0433a5f67428553e2dbc91be2cc1178ef971c22aa456b04d1f26d848de67bf6bd4e9dfc51762f3af3163338ff08f0d55db8153fbb7cbf1e87ba64a35a74288bc4428037e93419dc0a517cd2a18f8af6451d30c5e36093e8ede8781568f7f10597ceaa64c62feea48699516d98003dbfed3236dd3c567627b4fdd9ab522f8fae671504ad42272b1f2bc876d517c4d4f177e5e1c5339e199592ad066f09e06923ce229c40ddf8dc059c9ea0efc4dabe8ef8c9c7eea85166b7a2706cc538e59e01c44e1da625490d509762162c75f0ba4a55962de87f1e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h50445031fad3cb6f29855094b5266f53b4e5510825d29a75636cec8e957959fc5297ee10d44de8b960e8f2d77be691e688bfadfc454d5a995e961cc1c9be10c2b7f34c589d7f87d4995a070c766311677230046f9f4da04d15b1d2e0447db058df58a32d65ccd8c16c3473e2bcbb161ae386ade8a1484d7b3cc1281537a205238bf3991b7738d68d9be55b58c40ce64d983f5b6a30c10d45cf2a98b548d38090ca6e6f79f4e4ccfdd6c404f0005432fa4c8ffb71ca01e7a7cbc8401a14c79349aaa449ff054aba77e5f7711e6c18fa9926149596d3107b2c68933ed0b9cba4846dee46567cfa179e5e56a533a041eff742ce01268784c1e18d60d9223e2cfa6bf63ce97692ba5a9e57db0b707ff4430eb52977055b369a715ec7d26e96fbb5530e976cdd0d241dcdc8f554f5f59dad64328c09231dd280e9a661f1662aeda82c64cd1d66bf2d3959a3bc064f7c951b56136444d222817fd20dc83db5d70c9626e9cf589404a4096f9455e95b804dbf7e49814d18595f823d1f646ca33bf5f2b7ff08662ec2f540a9b8c229b5f8294d54aed14114101177718c60e7a67db0f4a2b81a04b7f1117a26bc6f2af1646299441eba92501c0a705479e3554a5ba6df54c52428daa3efe6d4cca224b4a4a3eac898ce1c4ab11044aa487897682b97cb3cf47f358b7d8e1a3956dd91d95beb78cba8f7be45c7573d7012a383e5ef389839f64263064e28cf7a2d3e0f93b693a808ceead1e4c22eaea1bd19e2d9621b418cbad8e7b2b32d9e731a2ad5a37b476f05c565c34f73f551e5abbe5ebb2554f7e75aa87f28467d38da016430fc1a4b8a3bdbf007ab5d79cfa124d6394b75b9d783570a0df5603dbdb0f6b9bb44034c3e00bd9fe6d8e42fb6a3554771a09eb108e610867a9a5e8158177c0c2b02091b555e5dd9ed8a84b32bd60c092ab91634b79457d899667ca5beaf7e3f8d8bccc0e98a2819459df1fe3f48309b073cd25d36637a2462dc902edec37c0e312f13f3d405b54b2c0480f26448d85cb8332ea0b1f5e3bd5ca17d84fb5a7b7bd94fb3ebf9a9c5ab2fc3d9f67b9a142b7cbaabf5c1512873d35d09d6c60acfcb51663c6cea5ef6ffb227f1a16bed421e91efba40f5b483292f66c194eff3e707bbb3260a5b9e2c64f841149b680b4f561b47a2d911e4c515c59fd1a4cf3b23dfec2b8e47bbe20415957fad7bf4eb595af43c07000c239626d6fb9d65572fd971087e7a1fd03e2308c1182b95a16bbae712705897e3fbbc46cb03ca0b84f36f9bcb1292a221a05a639c3a6542f521196064a64a071cb075ac35c6d10cc68977f08d6a0ceb10349edd16193d77135dea714ead7e6eef7fea9ef9e493105f8084b8316864c21b0b2dce25362035a5669c48aaedafd280dd53d6ee23fa96d8ec9b0225aa7c399f6082fdb56c5b26f08ed0de13642cd4ec10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd5ea193f40806d6a99ee4242280a744cfd5f908a12a09139f13aa389c290e1f0d3458cf749aaeb20a69d64756119270b579a409eb031a44d9d378d6b16678702461fe6f2b7c780024c98808405c15afb5a32b5ae61b667507bbda048af9ae155be8c4ccd25789271b384856cb8cd04db2db9447049a28d36a84913aeba367ad133de75a4c94d725d0f4997056adc0aa2f8876b70df3c1e9568659d3583322c3bf512f61e42d64400083a2a6a4b76811d1b0a7f71ca62074fa6a67d8ffb7adef6043b7461eed12a9cfd6051969229dd86768cf8304f8d879c6efb026f7b8fce27c8af3ba7d0eaf0b60d89c60ce8eff087d5fb5dab2195a041e95d87b82a56e3ad113b9058144fe36a10f0a7560950311a212da33a6e7d57412ccac2cfcfe91b55d626f4e984fe7e4e833aa8950858b1d82d711b5a814a201958ba5aa871edd7a632d04a643f4215209fce6d92bdaba3672e7f9ce28e0a76e30516f7bada4a9202b64f2faae441308ac46ea76f6214730f5f0c2f6b1423c95f6f04fa0035b2dbd900dec4adcdb8801d49fbd96c077706497a37825f9fd6ea68951d0d7535f49fdb4ca996dbbddb0bec55a23a2c1f5e849be14edf6996e55bb89a7c735675353e21f799938e846efd349adf9442e8194312f659e2bb12c3fc4201b1b88996a8e411b202ccfb8569b69e43088be9c65a1f36cdf59a8224f86f8b812a3e0e6445911153b2e745e5ee2ac6d7f2fbd2cc6baf8f486ddfccd6227ac3e802ac3ff1b27b8b878579cda581dcbc7c69dbd7de3622c1c2042a2585c16144246ead9156e3017b915aa55697b815fc75726bf96d25048a445a4585711fb5d498d4811b4390fe30c47351304938189c0d31488e51df935f87ff1c429938ed19917e5980067b0060bacc3b679403cbcae356ebe89c3b8c154deccf2d2f4e74743d4ec1e7e4a273731127b9d77a840cafd9d7b2af573af15dc833929cac1a91993fef5fe26c631a263f2310cb9dd72f78121d64185c04ca8db22093bd7da24fe51098e0456c1c5d95685954a4e782970a587f7d40207e546beca431e928b7ec072bf0cb5449f84d3f797a5f3fe3c19a26f089e94a07dd535f8a6332933e94bd830b1167a95f22b8ffcc0fb5a3c6c0e8c5ca427b04ca89e3ec6b45ea6c7c101c6306c9f98be12ae983fec312316d7cace8b8c5a5160f5fb891f121184764751ac55feea0c7f14cd382f25b54204ce6640ed989f859d100ae6d9f7a29663f94184d9fbb21d281140c501af99bed59147da29cc6f54c6d3a5920ddafa338eb35a223c469d21457dca1b47bd330e2b774fea3e5fe1c1e0da6b6b8ed640861ddcace0ce506720f41991333b9a9a8d5c5d3d543e22fb965271f71a029b0c0304d498ccbd190b06d3428fc501503985ae9f2fa44b38d57b6e2e6c90ba534c4240ccc93f286922ece16a46aa2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9acab342b4d657a7399a9828f297578a52db999716e0a77b1f4915e29a6972315c7312f043e979ba826e69ea6c241c42d51f883e1adc41c56615bd2207f227594586511256909ed8c9f7ca064a60ab628b4535dc596969676359865311777ec7c80463e7ac2309e32c1fef3ac09bfbc7c433e0c107f1d5df9f4d2b7c180baccdc03a83941fd648f4e04e5ae3b323c77d17201fc9b8d2f459015213ead87ccf07dc6715d72c5e79e5281fb4f7d5c2e894481682ddac9cbfcf3d31e1eba4972e30c7810538e93c78094a15e92b46f15f44cc6df4727593336a5c3902736bda9f25f1f1d355f673c3213ef5daa885eb9f9993d3d103df6405e18b3fe7c84bf0fcf21905cfc59e64ed7182cbb2408ca3ce8ca4ec6e277da425a5474683aa349d9070f4a13069606cf80cdfd34bc96b58ea1b330111667098023100b5bf78aa95f4769ce34b80156e568d8111b934ae836ae55b2d66e36ac0305250cc92d3672db1825b85c4f859eea8d9c7ad17d46880662322396227f346ccfebcb0d133b52f3685347f09940012b15066a76b678bcbae7bdd63e367c09324b158fcc7ca8fd7afcfa4180260a86c90de808029cfc42987852f7f780aa092312d7b1bc784e6cfc7741fb2ac307e2e5c29f44986599aea0e98f819667a84047306cd5945e268a3cd97b709c9b14c64e9b06df04c037d3aaddd8e3a09b3280fc08de69948bbb74f911b0de723c12b20351857fe8689603ec17d30fce86c3b639bd1290c43e11956c5addbb66255392ad15a20ecc049d976b5fd4e6a81da1d6107cba502352ef94d537bfc40455c57382fa6f854be7918fc9564aa1d6913b9519cd2a22c3cf0f060dfde42d946c8554f7f49488d73c6d87c618468e33c72e9776b026a87c08e6ed69d9802feca82589df0f56f67913b8469144d35457557b3a968120bcc3d383477634fbbeb681eb49a6bc913e831abb47ec428108967cadb78b4c27c5e8394cbbe0c5242d40591cac2872d911380eada3f909f4ac642791ea29d2825590bb10a875803e29a3091d841f16b58fb842548f339b2eb76117a65d9f7c5df6c3de2f604b14e094896c70a2a5382e8514ce305151c17cdb11dad653815131fe6935fd5bac4485743ae1b00100c9875c2876eeac0c9f2bef8dc58204dab3a36136d0d15f035a891ad15bf3f3e472f17f177246145daf44e47e3d3efd66d37aee6201823479a77fd76dd12d7908e38cbb47007dc89a34d9d80f4d77415413650c06541f8798b327c46e720c58bd1dba5765dff42e812a0464ac5ceb48b9cc959163fd3ea790ca0b09bd17bd66b7b6211887926559b210e8f718ee97ff7087ffa1327606fbedfa4c4502021de5e9a568b5820d2df9fdfff3ed8392065f7acdb2a772dc15b3382a897d1e3dd5f8aaf6a42a5fb14378a7e81315684220c495a6acca183f898c035cf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h573b56f3bb82d5baa56531c1548c27c17c6eec8b50962aecc22701b75bb71e943d017f2f9f8c7177f1e2380de39471d1916fcf6a80b624801780d7313c367f5f42f9afb2e62e3d524f59ef8dcdd64fb6a089eada143abc4b280c6251f19103fd8feb2e85515c47bdd5c16ca73e7e0eae96f5acb240b45bad6c4d372c72053c73776f26ad2757b0d9f37e795a481e4ab3a5d7ab0d82cb325f5493b93723e5741974015b7dc5a1b2a2de4aa2e70206ac2ad95d699b5cc2a801c2ccfbb74cf75eeb9c0f625a7654bef4b5b377fb41d0400325afd3d3a8b3e4b5660f538246307ce290e5941d04504fc819260274fc4f9b786f764adcc23f09bc9e94bf2f59fc71c2694627fe3d1a61f79bcfb190353ef3f6fd04f47226267650c61a9c6f2ab0e4533967d971ccf61175c0881863960d318efb993d9d51156c80ac58b1437671d7df816e4f194e76f4af15d5d23c478e364db2277df21015533701006cde51d6617b6362854f41ff79097c5d0de23ca595254b3ed99f8e7154a84dfd0b86eb4a2ab8418960d4ff5e2f97a3877ded73f6a5a47bc1ecc0b3ba8efc1cb6347d7af05149de028055ad640e2d2f75a1da48a32880a8821945d9b5fd85fe262219e878cb7ef1ddb9324bf263b4f5ff7b7071167dbde4146aa036c837e554800a36848378fddc5610f0b6444a80b78fcb8f6bcc7f91e6ded1930ae642147d5ec3d0289117a090f695956cfd2116f8a51a5c07fc6216b508ed2a23903267bb317124bff5f031c1a05847855fde9350b19a7f37d517b34c1db43d7b3ccdb7aaac28cf91e4a5fe9e9b21bf818adac6c11b3d7473b85513f6b793d97187e0b171979ba41d7819eb491e82c2094c993c96b6c5b6a022f60d096fb1f047c7be7027c5a5b9ee7c088d3e952b0a47c934f6f0f9bd24c2d0e59d356f11a7c48aedb8d8edbcfbf8bc4f87d859cbe7489e9e0873392fa7f8de54bd8008edc86a242550d8bd3eef6fdbeebe8ccb452299201e4388a7a627c0976ecb29fd62df9410073e5d2cd462a422e25943cf00ba90bfc2220b9c0a5d27472b3bcd308a57bb7ad0fc485826a5be103a50eb3be60aafb3fe6fd911a4640fb965e6c5b85a56f03f01505715cb75ece5111a1591bede7bd5fdb1307cc1acaca63abc9d125cf1b490ee7cfa4b423a4bd2a03704a9daa0b2a7bb158c7b26c32163965b9cebcba2b39a8584a35b125504f0d5e98410fc05a9935f7d94b29e6a0b6d18d9f6af7cbd4eef819c938506a7cc245ad53ce8cdd09dd1009dc317d6233033a38771febabeb6ecd845b13c5d315b10c01d9dea243669790bba7005b5f9fb41e025faf2680f29b106b3fcf0ec883a54eb056eaa11600e7ba1bc44cf90aa9f9bbff73e7e7548269aed55cd99a91567e686a3725e6d7c8c5e2c986c7a39121a7e1499b79c2b8aeef5b3c06bb07232cfe65096;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha4110eef497bb37862d2a218de146ef7136584cc8553df141f52e1bc92739455e8d9e5cfa751d5138cca8db9741fabf967d87356bfa952ed82e34470744b0ced84fb951e66b4f27d42febab003576f8b90944c1daa86e5ba41b4a2a178b23131478b8abad9c55c41c5e23c6fe9733a8a80ccf2e3243cdc10dc105de97a80699317264c917051ec08edd23670e8a528c69126c50a432394ce0f034ec2513853596713e5724041ba905916fd17961042dff4f95e62fd49a6b2662c1cc33d005d75172f24ff697ea24bc15398fa687d3e4d3b997414326f1bbabf82cdf4c1a5de0079ae0c895efa59aaca18182001e0d18abff9397609ed4c61b920d92cb4ac889a7578c99c36f31b8923304de3a837ae3be6e85f6e0e2a51f4d4baa45bfe6aa434c289c8976654f8c4d8fcec22aa58bc7c4388449bb7768dc66a127ed3ad04d4331801a70e03efac9979794608148d51f956823725daf2282084be9e6b0d351ff867a52ebaf265fb217b527ec6cf5c87c188a399ec73fa33cc44c1d0f710276acbf7d11343678f575e77c1fba9235a4fac912f95d2f46c5e882043e26356ba0a0e288b3982e7dc606a6febf8526b4f22f1f3878e5a635c1e281ac44f4da2ebeb93fd916af40dea602c4fa5044d5a07c4a2a851ba961e85607e29cd4720d3f0f7edd1d0a6b42ed9e0f15dd89ff06493e5fe46f94772680ab08328c4f8b3fb4e40007f8ca1aeb34c607828697f862787ce29911311b493cabe4c56e48729387515a2f0572541d1821d2fc9bad239957d25e38d7142881aa29a1f624709ecf139e1b49bc59042bdc577a8bd8efdb0320102a220bbc84fe8851ffe07fe67ebe3faec15225fdc4f548575e52078d480e98e8403912b4de0cc525b7058c8e8485f117afe2dfc85e44e62290911082a18cbf134b8f3caf493f77c41020a406cc4651e509f5deac0bcc67a61ff4c9d34c85a760e021fc077714cff6a2c80765dbcb2b1a42db828b480d07c21323c6b74a344cda2ea2442af305ae746119f3bffb957ae6740d1f69ec15baf3c236582decc12c1653aadbcbca483f2a58a4191f444a2a205d43c346a86fbd4dfd4e8cc611ee7e2ac01381cf59c93011f17ad76d68cd3c754424046e9f27cbd9afef572b7c569ad6598b55586b3867f3decf8d86a4f00d8cae4bb6c41af4e7be43b43c8e4183238f0de58cd4ac6b48f4f0fb27a4fc6a85644204d623c93351cf7a8a09a3e7f5d489a98bc8f0c9a6baf007224fcc26d07d51a034ee36243626456bc02a1fa2f52c25f9fb393e4aa0566555663526148b30d30ce35928b084be5e800ccffe781c70d33b0d9d85ceb1b460e4587608c961cf01888e61412fd22ba31effdc916d39737552ad46ad64d225c99b5cd10e046b43a2ede86032fe937c25a4ca5a8409ee98a0bfea9210c2935cd1d98fc9bece55570394d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe6708f2e43addec9e3ab488c5068088ed91758a7e7093e376144a57a069075766cde0c892e8ecd4e39bb5df48c4f86b28bbcd4815937ce04eec872e802dd7e92cf0f22160c3c5d7f24727e6d71cc79835171ae334785f2624a270ee98fd4cc66e84662c72eaad21c90dc837cbb5e59f0d3006620f01863705fb5576129af41d4e61c2cd2f580974ac04158f81642aeb2d3daea91b782343b854b16173bdabef720c0722baa5179d950268fff71d8d1409ec35e81d34e2df7840bb896224c76205653f0c052f81b65de519a97f6ff176f4210a76885d530d5b55c35634dfb13b983912e04de672b998c3cfcd6c4f0acf6469c54e73fb3609b521c6ba33347f6189173292234ff81f6290d33a8e32d639f89d5e39ddb5e9843272376272706199e5c12ddab739422acb45a9edbfdb942a490b721e7310b3f69cb3b12a4dd3aaa4a9380f845692ba396001d09ea25bdd111d3012963af5fc02f64eb1a022e604759bb32115eb2f80c294ebd69ac00c4d02ce36461ca4f44193074bef870f4d8fa419fa7fb65424006f87569682d9e07c1f0de84c94fc38b53f3580141bea4ddc353d530ae8dde2a2675fa554a71ace2454813a125a6eb6df56085e53cebadde8a18279d4ddfc228deb8a7e63ff545555a39ede14176743e1f98cf5148c5110e57a9117ee55725b0921898ce3baab3a1e14e56c77c8ba99d91d877f914260936a74e4f831bb27ac92f37ac58a997701dcf72ca5a6eee28f4d0a517abfc3d2fcd853cd5272a66f7aaac75f69cd82393c1878ca52f21a8b8b97e38ed94dd243ef33721c4002bc49ffffa2f7c8e33e8933ada3dc319b907dd7c71ea2fde2e9cc55f5db509e0ced05f6f6aba18a5920614d8666898ecd2c2d183115e727431dd4789d40a3a8abdd09eadb8d2342178b71d86e83b6cef9b72b40ecb016969ad9fb2fae6cc1469c20f2e792554bd2edd9791bc00b8dc57b017aba2477454d10639d2e372470f0569d5b34fc726de4507639d0c3b7cacfe5f3b40fde5ab2177be9ba0ee35fd282a734f90811d306f45235a00cf9167bc5edfa79d667b9f232ec70f13488b9fa5d789c60e8d675b2b26c924139fd29be07af0349662ad844ae0a783877ca33877f8d62bec4d680f20518e94788f030ffcf780bfcba7932333618b27f3f8b86355cd6bd0b8938498ae5acdecc8c24c0f5c1e72b8beac533b544aecda2c1579266fe9eae226d4ff60918cb38975dcf21090aa20ca7ad4acc7029a234a9118dbabece889a664faaee6c0d000c5a9309f1d64dbef1ad5d20de6a4b6851b5dfc7ac69f349501200fd14473c1ebcb63a51b078ed6ffe22edd8e9792b9b3b596e98dd1441ba3055e85be9f787eb396c0cf4424d956e5b9d942ec0b9b6a3a4bb53d07c397e5fd623e81ee2fb833677985ba2b097b325d5e1e4058d2939cd54e4adde21;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h78280a5fb9e21cc1d5b69af29c27464a69381eac2f6755ad4400dc0d00a702face353f78fe31990d54cbb4859b03b223e59ef2bc465d8499e4250073aedbfbe6d14a7668c58a267dd748c32e72647ef56063480b3a91f312ba1923b81c84b9256e38cd8622f40027fe4e461cfa8649accd12b1c0dcc9e0e7d7d17902defc118e2a267073c261a07ae5dc316d0df511603fc94c1a301bbaa5d0b2396ce1b119fe64915e37daedeaf890e2066fe97aa62cb90084db85258ae584dddc85f1a93dc6fa4e1c8589039d9d5da885f6cf76080b7d4cbd083852fd438f8bd92dbaf6a11f3b1911b490e788fecfe3a5038e75809acddbe27972af8c9cccef7157edb0705332c22d790618bdf87a26941ac9d703a170275073ec8c373f533971ab3ae74314ee009c01a7443b1b7846b133b8c865cbdfccd4546eb828082df693e11274e29a47e2d05f4de6f1433d24314d2c15095bfdfa7c5858886971c76662363e489a07eef69d3af54ff4aef107a1d65f656d02e4f581e47b591a94a00a010385d130bc4fa9290cbe68f7512180cf3cec12f1316687d21498dab48f2871f549690e88d57300cbb2f8c5a06b9a76d759057280278e2945fd43cb38b82f89645dbdcc458dcdaf006d83c8c78b631a5564f2cf4643209109e4c25abcb94fa50c2e53e8c21c60190e54029e1bd6beb3f2808bc161ff72aadbee3c407267963e483fb91eee346f4e7569725d73dff9232e197d32e9685f3bcd4a87e112132c6d572b4aa8081a0e97981fa94cfcf5b19304204256e6c8cb6ab32577239d3a99c87c75b290e3248a88e00e58c1200c903fe5f657d0f70c28aeb971b722174379a8a939fcf171bfc4d6ace453fe0c894f2381c1b804505216c1f6c39384d21c9ef77d9c132ab343cf6e5703a4f9b29efdcb49955b5212be92ef5ff9fc966067680b7562c13f3b54e4f1eccee6f51dc994a9655c51157b8f1623dc4cc0808c1ab7c05beaa64790913e03757b63834807ec64492b4b31565bee574908e69a43771ff7b53862f95ad7fb1cab1b61cfe769d9fb09a6076f115aed819ff34cf58572a95d612875e7313f7e012a816fd1f07f040bb5f4e065ec30134543cee330f6fef38cb79385bdaa92d421baded2c5e369bfd4f8ea5a184334126ded08f61606535e122985f01984ed80d655272995a9da3f1257d05405a43f3806f0493003a831a311490f3c7cfb2312a46519ab0d6a896a2c66fcc49948689239521a4bc9ed7d921e5e7fcce7a3549c75073d9eb5c54c2a8de56e9ef1ab56c2fbe8e611723a90be21b6a746c3feee39628b083b388f103bca805c199e050023a06742e9d507f7c60cd96c887417a7029f571cf3c5587d536d1a480b70ae75ee564a3bea36ef768c6809c67c7d67efa18303efc1140a23ebb9983cecb741cc1cba36ce375f2f1a34452a68b2d71672;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha77d8c569e5e1bf729e53ddee2f4202f1ec6a6023ba2a9ec57db7de7f8ee6d1ee34411ad3524a3f4131e4bbd038aa37b68056a83119be5e4fb8895bad1f73650887212988cf2841c43fee27616d488f5af7bc745ad85ee53b31faf08d25c138700ad06bfb7a7f9a8bdabb9acd48c4dae91542b4b89d13cbeb921784d28f8db4d29d17b10ee098384ebb25931db1c314712f5b7a58cff401ae30ef3911929dbb4b857972790da6fe7e23e4f9d536f121d2661a697132d0da15e95be312ebb52803bbe5dd35fb57f24ecfa522a66f4239672d6f83c0b3c932b9289336630fb86b4411992ea78b6f83e550edf41121784f1856d8f98e7706359c7311178a8ce5b3ab1b29965718da8a8e3308b3f59bb739bcae529722879e0901d42418834aec09ee752899311252443b5d14484281025231e68f27b62840b9b4dae2da6a808d47688af1815fb150a3a3766ca7cf177fef00cc8ff9802b6d941e9593f3c23b4670dd598feb1ae353779c8247f4376a94ca4261e4e610c241745faaa4f67de13dee57c61e06621cb3164e49624bc012008423d5f030f53a5211d91c35178e91d9d1c123a1b28166d1aa34566019a624e24aed6a9f05af83504126f2cbe73a4a42b849bbb913ab6a6982170ba6c009f0db3f62fa446d85353c0ab463f5c23c25a8f5202b990074a53af0a40ff9b04689d08f46454355f28c6445c2f461f45950d57d50a47c530ab782db07c9dd28dfa0114910a5f0e5a32382382ba50c64b7d49f91ee30f42b15bc2b6b836597caf906719c348435b058a11519183d014b10637476adf28e0e80cfd86814bad4421177f3ccc75e7d6cab5b8c3e433b04a387f5b30ff83b6d12ad26d6249ca40b6006d53119460152a287d2293093108f6f65d67c6ffccae816d35873a4662e6160d98e7fb19860102d00cbeab38cdc989c9d67182566a2ea4a56e8be8e5c9e5525f9623f4740eceb55284c862cf4634c7fee9521fede0df2a659f390551cd55f895c40e3bda476b74bb3007242aaee81d838c3657b34b79b67d2702820c21b904aeaa1b1fd0bb328d1b928253ffa8c88cd89b0807e9db3697c64036e7b405fdeeeff1acbfd9b9186235ae5963e84a060b8324abae18322821497084881dd0da4b912bb2d87cfd74fe8e334e741040776048bcad287ea2b0837b58f54a0c2a84af2807ec85e23fd31ec47c865294f4b7dee71ec76bd1282e871ba1345ef5048da44443aaf9fc47b5f0f87cb557c70b8a90cb203de329b8b0b9e273c2ddbf5de0c616447c12143b12420210b0eccbe72d43f37a2610685225718e2019c9ed36adf189cd534fc004cf2e5914da74157c82b711feb145fd2473f5c4f59c2816681be936d50f5e398428e4c9deca8557d203dcfe60d596bc62b6aa2aad06133fed40c3121b34bdf08f397d2d951ffbf9f56a747ecd6f2d12;
        #1
        $finish();
    end
endmodule
