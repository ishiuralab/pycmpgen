module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [8:0] src10;
    reg [7:0] src11;
    reg [6:0] src12;
    reg [5:0] src13;
    reg [4:0] src14;
    reg [3:0] src15;
    reg [2:0] src16;
    reg [1:0] src17;
    reg [0:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3])<<15) + ((src16[0] + src16[1] + src16[2])<<16) + ((src17[0] + src17[1])<<17) + ((src18[0])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he736a888cbfbc061f7d22c205;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec79793d6adeb163e2ed634ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53a97216fede3f60610f9e0eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb85cefaf1321f40eb6a4ea11f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a86dfed5ff4942c8307eef54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30feeb2059587b4b84494d15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f9a9e27b725bcd99d0253714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24a3379622ba1f3c262d8cc15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac609387faeb8a1d81d10129f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccd15ce385794ce171270a23c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h884ea8fdd179f6d71151689da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had44c57587fb647cabe11910a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83b18f41f810c1809565c0d3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h644fe0c0f9459ef484eeee60a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a08775901fc4b4c27b19daae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93891122696de2edfd55ad2a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24bf0f15b71a2c6f9d69c8117;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8276a81fa8796ff11e6fbe38e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9235eea09ce04c4eacf1bc6bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d0a52590a420e8d4490a504b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a918e86faae947c129bb8755;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77e7e1cac526fb9f092a9b1de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95ddfdee46431b48510deb4fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc67b2c6cbfa49ffb7632576b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ba0bb56442c246d8d74ed06c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45ac44c26991bbb8e3555adc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23dda11eb0db25c45179753a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha31e4e2d8a4ba1ee90abbcf83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb6d9c33c48f001d09b8519ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h607aafd8e69d758785054c84c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h353860fd8bcd1690356a7e31b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17e687c9d52c0868707175801;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h131d0b62f21e4e654469835ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61125099b544ef3152f930ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde205ca3e249cbc5e838e97e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12dfeb5a0eb85a5ed8c4b3b45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6309ef6b2ff0bd6b3548eed5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99e1f54f476845b5681994f72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd058afce3e09e2e25b0b6a5c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h730ab224aa42dd4579139f622;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cc9be8ae528da8e2efc0a081;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h890a57409072594bd4eaa9b20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b70f92a9ce1c1fcdf3414f33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5513d6f565e952454cb24df6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5c2d6fca7f6656c1347c97cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bbad5287cd8f5e8a5e8e462b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5057bffe0ce076cce1707567e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39dfb70eaba0db55983c035bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf583a7417069295493b479bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fbd1417c32b8b4fa6e0266ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6834f91ec63b8e351e505bf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7f5ea5ba092d5ebad99c4379;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e6a093aa2134a9ddea36275b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7b4ee4188a1f7ad6dafd3988;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b2a71ce41a6908a75a491336;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a88cc6ffac36323dafe5d49e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20014890681bd30623788f4c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h272869ae6490fa3918c3594f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h503874f0b309a22512642404b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8627adc13e238986398dff838;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7912b2f4b5e652d3176c9da25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73103fb0c6a2bcec3dd78919b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8627dd439812221086b359c5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha015d6a966458edcdc3ac4c28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b136cf2044f1e56f2fd511ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2f6aa36a62ed787a22cdbadf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9faa2cff2a3b566e41327c245;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf69d0bfe7d5bc895246767a53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf86553e96c80885af3d42a69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h285f00a7f7ba4810f7f84cbae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4df7bf58e0c7c3d24427faab1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e7c4d0f65443ff6850d712dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4d985f1546478c951baca4d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22644dbb3619e5fdcd35f27e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h529c6ec9ada6d9974240ad529;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6c70694665ea7c2d0c672df8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbde894101e5b30cda67e2fd3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h320726ed86cc65caa62edaf12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89d2be67a134e922b5c54380f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49722c949289d5de88d9eccee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2542cd53650ac034bfc64cae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ee725467fe03c2893f9334c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6df32d18aa1e048511b5c5da3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77fab18e1a0361cd9563d66c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb90e3b512f77522464d9a0d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h664cfa0e2b71d74628ea68b59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f4d93d42032e43f07c48a3fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d6c64dd7729f1b51f8c98968;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc21ebc08980ced9a0540dd570;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1edf61ac45eb35ecd9c288a0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc3a6c44e5c3bb65060a9109;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7312ec6c26d3b706acb48c3da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfaf853f73d0336b04bbaa0355;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1687e6464bb1d05fbfa49e44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc80bf70b9862b84798141f5d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9aca1aaa7b21f9c353ef5869;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31dc86feb7cf5bbb7dbd02f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h261f592462d9bf9336da55da7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd18cd0da4588757396f4f6cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha53f388fd7b591a7c690f826e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5345841a53b6faa0f795706c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16a1e4b14b067f057d0443d34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bd2a7170cd01b7e6859c07b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h402390b1fd7909aed6a2e5f8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h770d90cf279fd577120c6a184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2badeee9f0faa49ca5f420306;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13b9f719cf6c4442fcd100bb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfebf063a49c94360556aa6d7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2525029717943eee9a15a3de0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9217c7adcfea93f22d141d1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b646b22a06cb7d1f97e85798;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he19a73703a69a30728a7a2f26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65df336319efbe131a84b8392;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h446a2903a5da469bb9f4dc1ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2bb07dacca4f84969ef5234f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a1c0ba162d6aaeb17106aba0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f7f50a6fcf62d73b21ad6ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2f7b71bf9ae0d512a43fb957;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2ab87a6d78d1dccddb5c5f9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b75343fb6ddd4a87fd1e8df3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0f0a00fa5141ac012354d9d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf05b932bae5fa2b74e8d1938;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h969fd63ffad259dbbacaf0764;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f86d3fc5e09b91c745227656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dc049663732c7370d007377a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8cbe71de9386dc45cfe1d32e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1c911de7a32c6dfca9b23d9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h844ba1a0656a2423c50215beb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef990b5e1a988e2b25829731a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h829a08fcb9af54195acbae68b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f67fef94bf566eac29532f4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb45c9921aa071410ccce941ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1387c2667366d5e6cb1f51b90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ce1263e7514d39b4c6a1814e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43ff6b67588597d8f9ed44a85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc85c1edf8c08a17b9d3f3af6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64cfdaf1de14e2041db76a24f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fba959fa8530f1881cb10876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9df08ad553b3af17d63d580ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c199fee4e79cdd477fd3d913;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h988b0a48b0cc272ca83aac879;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfde63ae5b151d6632b462b56f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha70bceb25985ac50d03c97701;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ac9f1eedbaca6c07ed003ff6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdf249363ec8b65c5823674a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6a83af9f78bfcedaa52d5a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h335d930f3f3692c8444e5fae4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7270cd9a4cf6b662bc6f361e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1006d5a5e79e7c138c507790f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc577ca36dc7697fc025652238;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1da455bfd880cffd12408be92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f18d92f7bbfe6cfd690dccf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf25d3f08d814ecff650862187;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf48bc18fd60c34cdf731cf458;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h376a330c9472e036c83af7845;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0cfe6231098bf09b160fcb54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf487c7ea6b43dd8760715889;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb40e355beee4ee876a6c51928;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b978f3062a5e7588cf24a4ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbec10ad6e20b2eac2f1808e5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h650c89ebe1296757222859d70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde65b48e26a10d1e051f502c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3ad0d9a1874168fa5b295021;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21c714a4b0ff5cb0feadef44c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca796e0a61264c8fcb25b2bd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46e63e651aab9586e216c16d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3ce66fb233adfb54bd9f3248;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44e9d180e99f599fd03c8f07b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb345fe71386e0236009b4e26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60a214b95c08173620b375f8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaf2df412f89bcc5f768b94ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42e4e400bd9315eb0cfa82761;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18b2b4f3c3e5e154e28a0ca28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8bb44d877a47846833df84d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc713de01d1e46199b72a8d6d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ab142de50dc7e2f8a415182;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h136060262225842abd31d6be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1de037149d1552913b2ea702e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4486efbc1fd48eed89dcce987;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadfe11e9eb55f7e763756c0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f9fd486372d7d9ea29803a2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fae91f5a08a8f43c0e27cfb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3c7fa0d7c0b2b7d9d556b321;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1faab277b526b8ab32e5d3e4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha05fc7749ee2c249949dc238f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fb95d7c4f453fcd6139f6965;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78cbdf182ab8b9bb3f99ebedf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a187ad1fd3cabb203d0c4325;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc89fe474dacfe4e8a6deae7da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9901f757ad127975ce4b5c9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h161f181bb6b9594140bc6efc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ffc0e515c00353962e734b35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fd4d33a99e6c0652653d30d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d9e80e0ef28ffffa81b94b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha632f0f33b49196f18ff9563b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3f12f09f987e8ccf96b58d49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbe67aae7b0fdb51f2933da74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26472cd7a1b2b06665cd92c3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3563e8cbe27338f84dae16a3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4aa1948551e026b4fca5a1061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4124e1ad5ec781b3c0b63265b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c6e25cab41f6df3618f5d5dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1e7e43f2929f6d976af3c1b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b178f4c78aa1857f2b1d9ff0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haca37fd13df138cce4207e764;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0a09ad78d3ab2e40ecb4be9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h312d258cfa91942f6b7d3d44f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h252c768f3654c5464497482ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha28bccb7e9dfcbf2b736ae0a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6544934b17e65e2f9a3883462;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ed74139a52a46d93650adacd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h543039a1cf5b8613f7ba5059e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79ed3c1f0161fa9440198856d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ecddc906401a9500a7fd35f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82c674fa2d5ae929539c8323c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bb5c3e6bebec249dfc83dd7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1096194692cf34455665a34d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha25aaac803697c96e17be6d19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bce38a8033e8dfae9a18ec0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e5949a814930c196ad159412;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39b7ffe6737f26cad598a05f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hacc47e175e3b8a51d21b41645;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ad67b1994c5c70cb145a90c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he44d5bd5ddceadb48894047e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2f626462b4477dd69b57efff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7adb9bb2458a8f9ed82f8b7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h344f171188967107c3933bfca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6529f248b267d8e4766ea2c74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h853f4da706c3149006c204a00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb99d3e288c9ba8a7a9d9c6a95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h229e1a6642929bf625f72175f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d8314974be7657750f5b6b50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0189e89576d29197ee7c57c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4ca3d28d5d5ba82ffc97087c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc74318cceccffe2fffe4968cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d55dd975d21abb1c39baa85b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb0d4e35de59850f0661fd37b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e1f204ca63acbb31562902ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c89f8741e310c7a92bbf581e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dbc76816ed621f2b7edc66e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca4c91b6939ee66585ccad03e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a300c4ba01e8119f6779396f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb14ce0bd2398cb79d7a41c396;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ef9151baa8088ff8d4d0be6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95bb21ce2a4c2c2b13deccaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca65dfc33eef738b8678d6ed1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc8b99841b228d2134a60d4d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h172084dece7bf1c4eb3851b1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7584fea7176ccdc19c04e570;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d596c9f7828135de1dfb6ac3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73b14a96b80ea2f69e7f09ab9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbfce23706783d4e11a4ec57c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7dbff1628885c805c069af41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h347927f6bcb15637e58d56cc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb24b826bffd92727bd9af218;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he24b2124328d034c3f65f949;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc5d43dcb9c2448d270a035d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cbe13ae05e2779d6ba57cd47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he41848e6fb69bfcbbe0ffc51c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac80839441d6b3598c079a94e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h346cf4ad6733ce5dff17c9b57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb52a9cb4deb8a601f61005cb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0e3a76609caffb45cdc43929;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff5d8e5e61ee9b1eb116ea2f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bb1e50d7b5b69106e489e566;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef09e55ce6c4066b8f46ccf50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h722b20225dbd84ecf352d4faa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4c7f9c53c39314d08428f4f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30be76e4a1fb6dc8ba12841bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c4727c3ccf436ea5dfb218f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1ac62f9f60f957e571115b91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da70f41fcb9a61767a67b011;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bd6663f276220655cb9e152c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb078cd159538fe648d7e6d9a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6590332c19772a722113c44d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha72b8e255f5bc071f1d1a562;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0c40b8242aa1ae07134d2ef7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5df736b4ff91959d0538b050;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb65511a4807e0ae3e1b431c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58359e1da761ed35216b43cad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d438988c098400a703405349;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha06aa0dceeaf21076e837b127;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fbb4ed006ddccacfcf3d82e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55918beda5b799ee1a7a93d39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he24cfbc6414acac3c6d498667;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbe6c106edf556c0e89b90561;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab0c52a5f20d9b738755be72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f40f049204901cc62fba51ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21da323e1255ff91778afa14f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7af42fe16f304661ea115d658;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeeedf15e22639b47c32df0d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c44fd4e38c4cf67ece992a18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37a83f550a987bfd0f33ccbb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h568d895fefbe44d904335b3e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76934dca0c90b966a31aeea40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h505343e16db9a780b534269ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2558b3102d63c4d74e2e6f660;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he64437073f21d5eadce5e3b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd615fb50f2dd92a8f8ca94a5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ff99dc805f2798523bbeebef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5aaee74d5c7e3d62524274c2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he30b3ab919fb9091797bd982c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55689cbca4c0ffa5eb2246a12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e022c63d432e12aacb7c5a1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6d179725a20329e6814eee7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h391a753d43d1dadf8968ec7c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e13821b8f74e6af12c550e0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf41e30504dd13b2c25a68d28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f910aa2eb105a5dfce09614f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29367971b271428a2a42c8f91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3de3e811a63b61d57ce26c6af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h780602aeb0d4df7b361b2fd84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6d6de063c9896ee2eced689c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7df7fe8a3ca6c59244e49bd51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ba4110ea3f9746b6a4f3e7d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ec106b905dc71a7db93fac1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8c77aacca31dcf7e4e60c1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ec5ca8be2c046001e3a9555a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e9a5d51dfe5dbf388bd8e8e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5e584b93ca85357969641377;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bf281766d3836812061cb187;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92dcfac9fda8500edd1efdb6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0674dff90ebbddd6029df68c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c033022dee3fddbe1618813c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca2d625c54bcd23858f336cb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff4b00b794dd21b92444126c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f5a8142a424a73d6f667e103;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6995690b41fd82ee578d639b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb02ec712c52a9cd09494d93a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bf6f4d0f21f030d3e3a1de69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25831425a395387213c1d855f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he709946b12dc03de91f6a808f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3847ad615fa9bde14d789ddfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e4ec12c105ab39a8aad6161d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8695def22c21491b1d4ba67fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha865133c4cf91b4cf0d1c1eb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb03fc8ec0cea6fbb646be5d1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59903f4267449d323620a5a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f62bad15c620a290481d82d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ed974841ace3205857049c9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc743fc159c041589a784946b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heef4e493625d6b07469e2c3fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5bd1cd2531a371bf200fef06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e3aa5d7e77068ce939210f6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h234768ce0648e54786603fd57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ec27c2e56590f0521b9ca091;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h925688c6cdf8a1a82c7135178;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69d5b85f47e76c35d1352b4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6aefc2e2097e83456cf1b2e76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e1a2778009cb2f5a0811e28b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb065b3778f74c90a25b88699;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc9dce71f920da8eba37a4598;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4478ec170edca4a0bb4c80d72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb27ec527de850855966934074;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e8d28fa804708f357753b1cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h694686a23d1782b09ea9a1b07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haaff7df8522ee6d718d26e990;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9626df11dbf7be120c4a234c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4ad0267c72d32c9b48723a63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75cf0c7d367cccdc462bff8eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5722c6fac07c13a7b624cc13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc622673ddcbbc0f3616a3fdf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75043869a691dbeb91bd621dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d835c6bdaf203caec5187d6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bc8b2074e5ede2d487c088b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2d4a0a7bf9abc557db7a8ee0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h923d4ddae085b327211889799;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3eb17d6bcf882bcfbf14e071;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he62762d8119ecc9cb89273510;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5b5b37a4393009bd0a169886;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fb3422d9fdceff65f5776c10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64eb91272deda118dba916017;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h303b04d940051ac342f7033c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbc94f5141915187bdd774d49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66f444e62f9d8dab1d90294e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62f282184018f427f7f107221;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb15cabea7bfd352bf03c645d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2c17fd2a414551aaab90f316;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8d7844bfea819deb8c2a8f84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde63a93d3f825279456a9886e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bacd5377b4e1fb301612f05c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24ee127260e1e86e8a22468fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he592ea9fb0ebc40ad80bb7298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8763e8cd1d8b3920b39885e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cb4efccd3927895a5608f064;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4573290c3a6c923bc6365d77d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb32aa88c4fb3858b39906b721;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb8386230b57fc21e00395a98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8225fbb1d02a157f77bc858c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b86824af232f1f15ca74b953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b7908b80a049995942426a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2149bae1f0e577e25b549ec7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd89bb79fd7342c8b3b5058a33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5b6b92f0280adc513a504e38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa0ffcec4c3bd71c34ece8a95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7dfdf9a77e459eb7a8923b41f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h675afb605ae69321ab0c95a9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec261a3df0a28f0be74020112;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47039b823f931379a8e50d0b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2353d1e5b25ceee052871d3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h497a87b65d697be008cecaf52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebb03769dcebae13a433b2c6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h743413000c7a7660cef9d990b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1e64cdb8913e0e0f7828e613;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2de91b3cbe0b241adc15536f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he048f2a6edee0214388c4a9dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he76462478669dd4aa0f26ffa9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea4ab36546f59abc41118a731;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9fd3391d3664b497435c5756;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4180b071a64779a3abb3ee376;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd90424a5f6af568801fd76a96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce4dd788649d247e40b5a714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h308d8b4b97dbb6709243eee41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7c560b1ca5962042515e92c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6404ede466dac16f03c80cfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd285ad4cf2fec59d6bd94fd03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58b78786ea2c97bb796aaae75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he937bf83ed4f66b8334af9c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce74de807d3bd251faa3134c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7057ac807262cee2ca465519b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h905fd5085f5745c5ccf9a6f50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h200907dcb2dff1151c1589ae0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9271c185de00f69a611c6e5fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e01dca3b6b5a6554cac154;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h911accc48324fcaa5537b4dbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7231040eb393d827ae1e55d85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25511a2ec1fdff9d6e4aa73bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7270da17cf60dbff8c262681;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3353887dd7eae7722e28ae911;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b6a720588d6bfd215edca7cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he94977aff6267e686ef2eb279;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h957e04fb68ea01a2904afb96f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34063969b84eafaa19cd58020;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h908a97f9d125d51f7b5f4a48c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e7f282673922829847828208;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he16bbc408586a61f0de8392d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea53819e8a6f53bdc8ac9ea6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69bb04561f21a78ad8a4de179;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he26a1c61187fb611b96165f07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3246d3e31473dbf39adbd2931;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24162bc2f653b285eef9c4f1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d47e5160d42dfcf31061e0c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65841071c6f54b725b3fb9ffa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c49acc3246b3d90873015288;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd973506fb5012da463c184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68e0abfb05c1b3bdb2837d36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b1b01207fe94e2658012377b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haafc0ed81dfc93db79f3b33ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cbbfc79c38189e40ab987c1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ace7bcd8c06723477ecf1442;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a8d49913c963fae1422f35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcfc8c1812e9e7b7f0bc9b86b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dd636e1d17654a689b7c839e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda76857d828bc6e5fe077c51e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5936a59b042d5213caf6e4cc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65679c691c988257de0ee07ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h738d049b08a3f329fb9d3f44e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ed513eee13b998c6e33ddd19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ec66f0207a18d492cefec596;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98cefd9a1f2ce0f5e8078bdd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59a314b355f500983887b7173;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4175025c8f041bfbe214a799;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb039b1061d9a890901bfa5bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d56a84adbab66ecd7ff3599a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd53421f31c9ca6a4d616c8352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24edde65416a91152f70229f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f5abbb0c64d5d8ceef7539e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b5a233d681b146f42e9bdd5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h287bb0de3dfc6532cca904deb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1d03c9bbe279bdd9d6ddb6d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74a412be92feb17518c2589a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha31b90aad464e538b9df1d91e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb40f71cb30c02ab8510f89061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e92ae1840b2f1b8bc5a41e15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0c054623ef4397b69361146;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44ee759ff00f41b19a1b28888;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10ad23022312d772cf487086b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80d6dd11f666baec01a0c1385;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9539eb12ae713bb0064a45a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h328a99fd38450b94d4796b083;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46e52150fccf574f5e7cfd6fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0dbcb0b1d96e6868403a567f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75afe8c7c5379a39ab60f5500;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b80b648cae5d33acc199338f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85fbfca167eeba65c4317891f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d7366a91fdaf29ea4ddc18b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd64a7ae99cb62fa92a721bc2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dc14fadedd072600f0e5b966;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4ad4b14ca9735c7b68aff5a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb46c72810ef751ecfee964e80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2026e6b2bc8d304421c1e579;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb60823c31fd8c6164a1002ed8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h653663b189bb3614a0fd569e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7c0b6f02e9794aaa3ec370fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h467d9da11d1d19263bad8aa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a314a2991bd81088b404a8dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1502792307cecfb777857fcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb46b9fbb2725625f691de18d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb40ad0ad9f5d21c3f3c747c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bc1f647c8b59335cf83b0fc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88645daceadb2fac7aa9171dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b63d5a14513e198fb9a3f421;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd449a7697dc1e0241247bc51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef61eaa4bce1aae35f0990ce8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h771180d179e57cafeb1ccabdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ebf403f9f196ab7aef62194a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d4bfdeba8e751e2680952313;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc51acb78fe75e5683b182465;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7218508053b0298b81e15dab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3430427bb0c06c1c85ae4ce5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha72852e5f49acfddac9cb2c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2385e8d525f0c3c07a7a5f8a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5316b0b9feb7158949e88344;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h247ea5e3a39d8c09bcf97b3ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6181bdca541c993bc1076c131;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52ced7d2b9067ca61f2ccb129;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19b3dc58164c8b0ff150422fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc753dffd65fca0a67e00d9290;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa054f6c59ad2334ebd22688b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h968d07f5fdf82570f1c2b50c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0b07ef741aef27329c745de7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6879727b4764eac7f7aab3c1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc830384c7c3d97d2fe6543ac2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9603bf2bd1b34dd2539cd8f90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3bbce5c4c913199a9b05e2d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7455a3cdd166ba9c3c984deb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5152c693ac4d002e4b62909fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ed4757da53fbe1d5d4459446;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58400dd96f6c27d6b6c7d87fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc77b3ecebf554b285d109256c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h771120c25214025282bb36a7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'headcde70fb8b6836b944fe228;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bb7046e79a3beb6763163f46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc85a75c3388c233de6f8f1a86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da5db4181c94618017548f86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f48ef2c533387dd4776f8068;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ecaf5f5b0e0b5aca7429fce6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3814b0166e75b3762aed795cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91d8421e235a8893e9d62e6a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha528c7129ec3b5bf9a925c7b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17b05b4ad7a65d9a949c6e95b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h315a47d60063b0f19e37dfcee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1002b2fd5327ee44e547bdb89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd566b741993439920b1a443c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2a721d82d7f6426da881fa0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5fe20d38dae504a69e30f987;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c5f0689aea937f5c36571a04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc38f288f51e854792d382a2e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0691f2f5d2070481af959979;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e9d5ff6456b7d6c388d08e55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53d7ce335f6272510b8b2945e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h498b58f7f91fac723ae9a7fd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dac08049603599c34030ad8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h557080fb43a76aeaa2164ec8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h192f703452be5e79962de9e8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h187402e6b53400587e7f6acfa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef65bd538d7ef007a62ca446b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ecbe0909af45843562da2477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8f9185b069aa1c6a438d67e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he22503bbb9b9cc432dc065416;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97e0668012b71405ef9fc0bd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f818df81dba5931adbb44dcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb680515db7c0095341b6bca8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbcf6f6a2418272a3ae2d8286;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3899ebf16b93ff9a1294c8fc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cabf13290840a7f9582f8f5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he220984230ae0d92a900664b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8bb49c067bd2e9deea0e4081;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ee4702ca4749cce5c87d49b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73b223d7d4f586e7013e1e4cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f6490f737257d55d56eedc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54a6fb863edf0594269b4eabd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b40bde58459c16824e155bb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d8ed8be5e94cbf8701decf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb55eba44cb4522c48f66943f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf00211251aa67c480c9953f91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2f7bc0d02ff0bebdd0f2c184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7540a07d8d42c45acd1c29236;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6028745b8f84759b1090fd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0a33a4da77ce47c9bed6debc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2bb7f21fd1d1c5a46ae0a2df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h364ee91c0fb078d162828f101;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c843c85dd064d3b49440437;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc030746a50223b5da33f7768f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72797184b01d2377518c5a0b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha047b2a32759347afa33e11e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f575722eb80fab1dc4b017ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e5578f0ffc6a7109d0a02251;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20992bc542127dc90049489a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18f1f74a9a423103b76b5b047;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccc4fe1b64f766fcc90d38fba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d637a52958c6e3182f863f55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h737f54265cf2296659b795690;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h555b21c2421ad14619fae132e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0c5365291e15f4272077da3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h540b5e60af87f7db8d1f6b062;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d5202a78583a07906b751e92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h338adc5c573f27eba217e7523;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h448424653a091e7a38edfdbd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h937ae62f1df25b0792747cc8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac5b7a569eadb8d1bff8ebdb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf8f2efa1e6fb13953dcb901c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he46a0660fafe40609fafc56f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d9e69ef87b67ba2a8abb019a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8c936d7d54d4923145d34294;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50a2e44a6a93fe580af299d67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75aef6be7f55acecb9973f3de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f4d3c0662ae416cc22e0bf48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h951eb70a39a8b0c6f79d2a24f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37b9d860de114cb884114de23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9685596b9f93bd8cf33118119;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41b3f9e68a32031b58b5f6ac5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h669de302ef087963f140f1cd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5197a98d0f228244f30936a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba20175272679fd0bd1e7aa8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab62aa874e51a14f34dbf5047;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95feb5d0e447f3ddec4c29607;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf11f2bdc2796dabb7486e9083;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe48e5ecd597e273099f09ace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9b7201e74ba6485a714be2b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb0e8e4e76a6957d5c8e1ec0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6743b96c2aa087fa98e8996a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2e9f505c0bfcf5e62d15a614;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb91144224d5afc6fe62aae335;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb92ebd01a657ee7fee0be565;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3848654ca01b90c8c821a7701;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1257c8fc47e026a15cc1a103;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d4c545a3725eaf006bd02dee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53bdea1fd1e73fd2d3ef9e556;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfd94a1f6dbb79bc028093995;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf266dac62c0948ea942f6b0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h821665e4e0eb07d934ed0d677;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64bf7aa526154b9f0271c2073;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8585b60e353dbfc174b799856;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ecd89924886d82d5dda9ac6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64c0f170761c2b8256308fa8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha445188aa439e65258d9adf32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cf1d28bf37113e7c8845daec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a8b03120cbf789b97c0281ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9605028dde2709acc23badba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4297be18110509f1d0ce07b71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef30ff639c9629bfcbbbeb9ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd157322324aa0a2056edeb520;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde41d6c6ac751ee8409745771;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68548cc8645af09cafc4ed233;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcddce9a3d19e9f2d76794842;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d62e8cc15db0b0fbc4dfda91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbee0b50bdf7d143bd58fd3657;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h796de57bb47b222983f2ebcbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h798df0170c43012f3970c1e2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5c18311d368387b650411411;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65b013d713bac0ebbe2d4822b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h750f0eaf7f040d40fa6d0a0e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26f5ee4b29bd1d9082a34d774;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h898fc03c51374707df8c64476;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf826c5698f80bfeeb82ddd030;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a3c9d013149735a892a88550;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7459c7b842bdf88b31be131d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0ff0f4ae28d8e9cf35fe26d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he92da4e0545728fd495c6fda0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ed3b94d164512b296498a223;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e8c2d18a9f15f8ff761664d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6d068187487fe9388ad401df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c7d4893b74696bdef8994b39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79081db5132b9d43c2b66c260;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5ba339b4bc5fc44787ce97f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32d28600ed0711615bb4bf299;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c33fac80f9e9acdf067ceb5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc1416237ef2155f9e31913c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44ab2d6383c3852f6abc8da92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63fd7f680f1a8ead87fb689d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1884382e5512fdf2bf2c2ffdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5567cbd216d01916d891a857;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a158fd1c15f81085c2f79405;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f5bb1d54089b494efde7c181;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8631044e1e2448751b92e40c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7e3cc5c873c39008aaecd38a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b8e82ba43cef51169fd54e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49f748bb5d9460d200e3f873;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893e687503945539d4e311724;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87782e855c314e14339503c97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9600e002e167327b84508c2ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1b6afaa0339160ed7e0d37b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e18a75de9f6e955c378fdb9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d502c439cd747e8b6769fa84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17038867923c3625b94617710;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d6648ebf09e808bb4a51f31f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habb67ef116f8e2689f5460048;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b50802bcc10a5ccb6375d44c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b972ac8d92c743635bc759a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e75bf29f46f29814f0c023ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc77becf6658c1566933c970c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18972f2dffdcef2145d652b7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61058a9a79f9c4e3d72431394;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10e5d62ad09cd2918c4fab565;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fdda6141084bda1ff2c89ace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f3dad0d31b2102b676812dd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1abbc8d815d0ca30bcc5fb4e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f04acab371e94d814f780b85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bd9f4c6e7f01b840ca26667;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h148e1452453408b8937da88b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec238b03883fd1d963b25ecd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30ae9f90ee6f4c2c35a03d5d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha79422107850a3a59c592d1d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b1909e0f35a153b52a5b47b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cb22c0776e8f2f1d60b85ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ee09d3fe7515d03919015520;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84452b008dc61f5ae0b91c4a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4899cb17c70ae3f07fa89c3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34105a16733d0383611151d74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed6e5dcdd9d1005ba52428bcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7332d68b1e8c86abf1993b1aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb6315473fc7eae4716be6ff5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16f3611e3e0887c0ab833b144;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4c81882e5007e97858a65970;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h285e7e26237ac87b7b43e9077;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7259007d95fafaff1c2d78dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f47d5bc87dcf52bbcad6b946;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3de939cc8ac71c7c0bc494ace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f905750ef41300c8789a97fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba1c5a988afee64290ce126dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h290226d91b6e02cf28836d5c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8d5bcb91fa763c3ea983b98a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bad5263878fcb0d3f8f0541e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e919ca10d7bad7bd14911890;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34ee88ae8977ee937da766892;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1c9283f0a1b6f85674e54ec0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha76567fe92d42480e4dee3e35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4280f4d87139db8e22decf07c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cd61950ab82fa9a7cb6ff01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc93da93aab00860a005964a58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50c8171583958aec29cbb6c47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba29f71e3827f897aa590cd75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc21f73f3732b9e1f60be65eb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85d8199a213eef3b7263c0847;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecc6591049e64d11e37831c8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heef1681b105c5602b17e444c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86197149a679f7e17f9a69d03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29b2f7fa8e7a4b36aa9bbc33b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa033b736986fe55b5603d5de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h743e5f7352ced55a6e28fee1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dde51f7fdef671896edeca6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he89cb7e678a573f019779c0e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cf3e4e377234b7087644099f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0d605e689b95135e218635a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha73ebcaf12dde3c3e134dd05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8b25106a0810f637d191e4c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ec0f2083112c4443de1ac732;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb93b201f1e1ce541a9ceb0b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb2414093b97d458f8c8c7514;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd451ae38e4025456b386f66e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6dfd2287797ca25bf851bfa7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf469fd461ab483ffb5690c24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3aa8895395d9c31fe0747e62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfbe70bb09df0bbe34e3d11f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha35af25f4946a56e58c8734cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h476910f0385c46f8a7d77e78c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20f1adc1eca6c01a052df5e1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2856311d5ec2e5f91b2a1256c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d408032f8f1b41de94d4e9c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h168a201ceaf7f94870d5ef3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc6839a448c80ebec49cdf661;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8473e3920bb600e99f6cda6a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd78e34602a6d4d35c4fb84cb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1961a2f009c073c44581298f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cf3a31e14ed7a4afa2763794;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c149d2eae060087f84c83fdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3551d170b700e5e0b4b0509e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27458fdc73612b59e267d042b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8d666abff2c7d7e78c9036ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14053b598da9c96ec3c03f858;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5992fc24c98db729af917adfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heef0219d9f039ff8cb7bad108;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4aa73c3c08dd8895618435d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74715fb4ceb879b0822527c47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e24b352f67c01942610326be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a662bed662d6892e91f9fbc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49e4aa44bcd067f13e5168ae0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc67205aae166c69ae7911edfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he39d237f7e7995a71c2ab9a6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1382d8c6c2e2eed13e840dde3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafa88ff740ef0971f4cd7b8ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5890a80c2a8308d0613d296e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd08c451a1b5c32c04897ee66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e7a1eb7ca435d27a0037d8e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f19230da4ec38ebca3734671;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha89513a243c40318df892196c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha55cdfcdb50f0f96d6386027f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec60cf339ca1027b03cf49f03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81d84e485438bf3b82bb64e8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54fa87b69fa09f01de33371a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56490e356999e8689adee28eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd741c5753fdb9fe72ec696134;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedfebc1269957bffc0f5defa3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14eccf4f41095957f1bb23526;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e822a46a7ec8644374ffd656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf87cda37ed619cad256971627;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a9fbf80776df9f4ce67449c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca12b8ddc7fde165b5d7dd353;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf938e81f84da725caaab1277;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he85a78cda4b664f22617f0cc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18155c0128de7eda9c24f1e15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c3730aec5ce6fca294dbac5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd44ec9eb969606d158ad3f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbe51fb2e69713d07ba9fbd75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b6c17835a6c8653577652960;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he929164ab5d44202f2e8e2a8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddf56413629e0c5be6d275bd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9163b1d278f3f0f6a1bcb7c54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc2c834834995ea9520373acb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0e62716b0c26f14926cf372b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc4d65cff49e24bced8a4f054;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h506ed758dbd82b4837914ac4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5600c8108ff752fb64024ba1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c3ce8e558c29e05f1b2480e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa3be419596db22a469d8fca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h865b05674ed20011f5ff9e172;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3ae1100dd877dcda3f315025;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdce965f6d07116689b9ac3452;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4294dc43bd81264921a261fa6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcbc4749a667eac299e6a6114;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a1a0dd67b9210342c810dc5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h313c62d592930cb490016ebf0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h290ed83286dff359180ef61fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc07e1f8dac6e0ba4af1135a08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2a299a0e20574f36bac6daa5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcbe6e10028ba9efd5df58c37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf9b19744c5eb9f1bbc0b13f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa96f91cedf34d0b38d2f3123;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0a6e7553ec0458da1fa3665f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1cd460f9240342c9a62178203;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38b5abdf90203ed1aaf94d9c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61eece4cc5bf3f31d3d833afa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a2084f9354cbebca3168c416;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73bcd8d2621160405d920c2b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9578b2b175171c8a95f99b1d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f2d02d82b3a04ef71779b031;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fde16c541cc49cd2e182c173;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbcf17b0b1dc54291a1c33eb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a608107506df56ea46686cc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b2dcc4a4bb7e9e49a9835225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf25b58b483eab10f8743a727d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he23d70287cd879a7d5a493683;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb496e58c35e13786ce4bb4423;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h550d7d54456ea2c64db781ef0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d4214edb238b75b348cc03ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc253642951196bc69a38e5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he77285483e33297d14de37d27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bb2aa77b896fd48d8f60f388;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3e7b137b8d4cd9a347c63d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc855eda376a24065d7b183281;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f4f1fc29a8fc3bc674d7c1f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83d63535f8bf0cbb1abf20c19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ac7327357fd758fc64a5c392;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb168a2804f4ea9819995959af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42fd5e6ebc5692f97076b5d99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96849ec46e01ec64449b604bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e8ac181e110d654895cb63a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8841a5a1e675e9424b8f42f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h726f72392b79a142e82f95af8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57fed2ebfa29ffb6a2451109d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedfabf434b1a0b4c661bfa266;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65574b33d636cac2b53c976ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93d3682deb951b50534b47a51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd33004268e3b0859b390f164;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3b6ee4246dfc796222d23332;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e498a6418d5ac84f95f8213d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd705e0d8a85c66439a1c0a1dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49bee82cc2e5a22be37f71bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31f848948b8757cb07a2a154b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21ff172db85e956f04214329c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf97a47f7da70c105abfef936;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52584a1a5a29d3d20ced3d214;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5996400f82c31040121bcf2e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29c4b2e5372dbf6c69b500a6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf63f4840f1a79e15a7675cac6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6794c0dec9ecdb0d95c0777b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd23a387745852116253d1a90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9e5fb92951d575cf53201c42;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75c3d06a3c98e266ed9de075d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h124021a0f4f640bfa8b274985;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab363aa581197ce18a3e21a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc44d1b79a9753eb7618308b62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h392338e02713a1cb84a1e055f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h738a94ceda2241df36dac2714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had67386840a54d3877d515245;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c08dbf0642d298223f211d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94874e3bd4d44fbb96107d1d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e5c29dc4f360301965b5ecae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc6e585c30a4344486287a331;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha52860b327f21d87475b30d8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc3017140bc59d30a0118bc40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96a8ac5b7660c91bb01a874e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec2d96b6a9b05270ba11d1987;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52c0d51553c6acf005f985511;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3536d01f8e0be7ac8e83193d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb26a7e3f54d861f2a20db773d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96dbca3dcd0b28edfb0edd14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddbc8a96ff85047b0438bb26d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h203bf91c0b5ea97db5e89eda0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h163c281551c822f3b2fe4e997;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf774b0162d0ff235b6f8c47b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbda7bd85e4f2024ed6f3e3e3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17fccd95f4f0f4e1a7e96be79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h441bcebb285a6d654b909bd6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha200bbfbf6da6f4a143ce187;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4a228459a182924280eb63db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68636569991bc2a33ac255313;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd30682aa74753486148c174ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0acfc15a85563fea27135a80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h575dc686958f9fda1437d4503;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b465657370638848f71b79f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9a144e0b2b65c0d836b82f7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec9466cb3d82bd34e46666e7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7900dc006fb6feba15fecad7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28136f1d3d228fdc0ec22cdf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde6a3ddc2fd590b57e840d339;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61eda6f0f927b6c7e0c8637a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb95d162e61117c7d885930e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39bbefca0951dc9767b4d849a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5ebfff6ff3f47302fdbc2d5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd43bdeba4f3dba0cb47cfd202;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23bab524891d759cf14a0ca2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fba9fb2ba9d7ab77990558ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4641e9bdfe56f37248b3dceca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5658ba185391f97e5bd1ba8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0229f2636ae71aa5ef795702;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd6e5082bd8b5558caf08ce3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb527540f2f82d940ed6bc697;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h184936b1bb7c0b6ff7274a7e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea365e9fd0f1715cb50786df8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39c2fa0bcabd76b90015016a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2e30f98f2b0861816a20627a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f1e9a54b017232e5b58c3eab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89f9a69353f29661e4d6ec875;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8b11c89b7875ba3c95e6a24f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b4cd000b9d828af479871ef7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8e85b0753e613e859256ed41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc297037a86edb67dad6a344fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb2e18baf56bbdad7cb7651d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13ccfa0b87e1bde53ea21cce5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6818a1dfa9d419739679ea969;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6aaa87d28e376dd9adb12befb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2ee77e88dcce94885280c71d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28a549ee8cf399890d446c537;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6ab86fd3b76087279145d548;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf746bb019801c1ed82bc2d60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfa4b6d0746b66d0069bd8983;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe935cf85eda514d4987d4461;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h321c2cd3cac779cbb9a77863b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa8c2fe9ad32b8204e99c1e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83926cdb79239dfe53418023e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e09fd8215497fb763186210e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56e7e06e6ae46159e752d39c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b8b9c4a50f0d3e5f75e76dd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86bd9ee96f05d351ac67cac31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2c5c5565ec8eb4284b6f3a95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20478ce1ebd9f6f4aa1ec8a1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34f0b269566d09a876c1f53de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h452df700375d92ca6b38ac86e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67e0cbd0f3feb1eed07640afe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e7233b8a9535386e6c45f65b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab7a767d0be12890cb7bc187f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0e9eb92cd5d30c2372b98840;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe4c7dd4aab02fc5ce572ef56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88e7f4bd1f294fa1f13cfb02a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7916bd5d94b884bbc125b3fb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51ebe33d67da0a343718632b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h824ba02c1345e9a3bcec6a1fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5267e140a1227845b97f9646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7d32738bbec21f977f6fd589;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h191daf7ec333adfa73098cff2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he720c9fbcf73f25012ee50818;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d91c9d29f9636200a01f7945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcffc54a107faf1d4b4aad4fde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd96041b50175bd47848050f54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11c5ad95eb7290230958f96e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb26fc637056da0f88818b2c26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d8bc04e837b39457c27aff81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h406f292d57deb067f2e603b12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h102d6566c147a535b6ca7e7df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18f1db5534a978b3354e23699;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b73e58a6bf82d4539b115fef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30592f8db15a5325136457dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68bd7a497e2c7ce3d2010a5ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c6c80b75d71787f0868a0085;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5604c299a61afb8f696ce7767;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86b3ced644e8d0ac2b1a0a479;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha408cd72c3ff5887aaa24dc06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6365731030fbb4a23fa2032c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbf737a2c77510f6e58911d0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25f4a0e6850455f26a66c2182;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e9b752647fc800eef4bd16c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b88ca01650650179a706ad16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78f30dc270b6b7e727a9f170;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5503831293a22e239cb86c3b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h372a3cc9f2d871db6a6acebeb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he23cd20a9922d10971708eeff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7b48755ed5885dea203ea812;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49fde7c69a4d392615ae99a6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab2b890221570fdc71bb0876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16f148190c503e59541e93c65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77416bbd460ce3d460701846a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3b658256186478910ffaab4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66d274f70294d51df51c13dd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbda29fbbeaa774f8c2488f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h269722569d610ffd526f83ac2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab48d81c13dd4e72e82ed8aca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94836cf848fea06204c1dad34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ea845385a5d3c9e68181edd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bd6f7465fda2eca2ba78e6aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h267345e3cb8eb160b7fd3f0e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha19c4f8308f79bcf0c80d6e57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h197ead10fb92f86adfcb8b27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1aa414cc47a3ff290ad235129;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91afd7baf02c09045ab51c1cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b73ab0d98cced590ddcdaa78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79b37e78c204c438c2b7d515e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70e9ba356fbf0934fcb249533;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h176e6bc4f4260280a6cf40c2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h359f03cafa9193b2a4dc60cdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a30eeebb178d76242991763d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3551e22fc8700d84f136cf235;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h220c8867e8d3fa60504622db7;
        #1
        $finish();
    end
endmodule
