module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    compressor2_1_512_64 compressor2_1_512_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
        src32 <= 512'h0;
        src33 <= 512'h0;
        src34 <= 512'h0;
        src35 <= 512'h0;
        src36 <= 512'h0;
        src37 <= 512'h0;
        src38 <= 512'h0;
        src39 <= 512'h0;
        src40 <= 512'h0;
        src41 <= 512'h0;
        src42 <= 512'h0;
        src43 <= 512'h0;
        src44 <= 512'h0;
        src45 <= 512'h0;
        src46 <= 512'h0;
        src47 <= 512'h0;
        src48 <= 512'h0;
        src49 <= 512'h0;
        src50 <= 512'h0;
        src51 <= 512'h0;
        src52 <= 512'h0;
        src53 <= 512'h0;
        src54 <= 512'h0;
        src55 <= 512'h0;
        src56 <= 512'h0;
        src57 <= 512'h0;
        src58 <= 512'h0;
        src59 <= 512'h0;
        src60 <= 512'h0;
        src61 <= 512'h0;
        src62 <= 512'h0;
        src63 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor2_1_512_64(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    input [511:0]src32,
    input [511:0]src33,
    input [511:0]src34,
    input [511:0]src35,
    input [511:0]src36,
    input [511:0]src37,
    input [511:0]src38,
    input [511:0]src39,
    input [511:0]src40,
    input [511:0]src41,
    input [511:0]src42,
    input [511:0]src43,
    input [511:0]src44,
    input [511:0]src45,
    input [511:0]src46,
    input [511:0]src47,
    input [511:0]src48,
    input [511:0]src49,
    input [511:0]src50,
    input [511:0]src51,
    input [511:0]src52,
    input [511:0]src53,
    input [511:0]src54,
    input [511:0]src55,
    input [511:0]src56,
    input [511:0]src57,
    input [511:0]src58,
    input [511:0]src59,
    input [511:0]src60,
    input [511:0]src61,
    input [511:0]src62,
    input [511:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [0:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    rowadder2_1_73 rowadder2_1inst(
        .src0({comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], 1'h0, comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      input wire [511:0] src32,
      input wire [511:0] src33,
      input wire [511:0] src34,
      input wire [511:0] src35,
      input wire [511:0] src36,
      input wire [511:0] src37,
      input wire [511:0] src38,
      input wire [511:0] src39,
      input wire [511:0] src40,
      input wire [511:0] src41,
      input wire [511:0] src42,
      input wire [511:0] src43,
      input wire [511:0] src44,
      input wire [511:0] src45,
      input wire [511:0] src46,
      input wire [511:0] src47,
      input wire [511:0] src48,
      input wire [511:0] src49,
      input wire [511:0] src50,
      input wire [511:0] src51,
      input wire [511:0] src52,
      input wire [511:0] src53,
      input wire [511:0] src54,
      input wire [511:0] src55,
      input wire [511:0] src56,
      input wire [511:0] src57,
      input wire [511:0] src58,
      input wire [511:0] src59,
      input wire [511:0] src60,
      input wire [511:0] src61,
      input wire [511:0] src62,
      input wire [511:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [0:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [511:0] stage0_32;
   wire [511:0] stage0_33;
   wire [511:0] stage0_34;
   wire [511:0] stage0_35;
   wire [511:0] stage0_36;
   wire [511:0] stage0_37;
   wire [511:0] stage0_38;
   wire [511:0] stage0_39;
   wire [511:0] stage0_40;
   wire [511:0] stage0_41;
   wire [511:0] stage0_42;
   wire [511:0] stage0_43;
   wire [511:0] stage0_44;
   wire [511:0] stage0_45;
   wire [511:0] stage0_46;
   wire [511:0] stage0_47;
   wire [511:0] stage0_48;
   wire [511:0] stage0_49;
   wire [511:0] stage0_50;
   wire [511:0] stage0_51;
   wire [511:0] stage0_52;
   wire [511:0] stage0_53;
   wire [511:0] stage0_54;
   wire [511:0] stage0_55;
   wire [511:0] stage0_56;
   wire [511:0] stage0_57;
   wire [511:0] stage0_58;
   wire [511:0] stage0_59;
   wire [511:0] stage0_60;
   wire [511:0] stage0_61;
   wire [511:0] stage0_62;
   wire [511:0] stage0_63;
   wire [118:0] stage1_0;
   wire [168:0] stage1_1;
   wire [220:0] stage1_2;
   wire [321:0] stage1_3;
   wire [250:0] stage1_4;
   wire [216:0] stage1_5;
   wire [179:0] stage1_6;
   wire [339:0] stage1_7;
   wire [238:0] stage1_8;
   wire [362:0] stage1_9;
   wire [152:0] stage1_10;
   wire [317:0] stage1_11;
   wire [218:0] stage1_12;
   wire [184:0] stage1_13;
   wire [255:0] stage1_14;
   wire [257:0] stage1_15;
   wire [223:0] stage1_16;
   wire [217:0] stage1_17;
   wire [241:0] stage1_18;
   wire [218:0] stage1_19;
   wire [243:0] stage1_20;
   wire [204:0] stage1_21;
   wire [200:0] stage1_22;
   wire [298:0] stage1_23;
   wire [234:0] stage1_24;
   wire [210:0] stage1_25;
   wire [188:0] stage1_26;
   wire [211:0] stage1_27;
   wire [248:0] stage1_28;
   wire [220:0] stage1_29;
   wire [232:0] stage1_30;
   wire [211:0] stage1_31;
   wire [414:0] stage1_32;
   wire [209:0] stage1_33;
   wire [267:0] stage1_34;
   wire [190:0] stage1_35;
   wire [330:0] stage1_36;
   wire [302:0] stage1_37;
   wire [276:0] stage1_38;
   wire [196:0] stage1_39;
   wire [229:0] stage1_40;
   wire [276:0] stage1_41;
   wire [228:0] stage1_42;
   wire [243:0] stage1_43;
   wire [268:0] stage1_44;
   wire [188:0] stage1_45;
   wire [299:0] stage1_46;
   wire [277:0] stage1_47;
   wire [210:0] stage1_48;
   wire [241:0] stage1_49;
   wire [216:0] stage1_50;
   wire [226:0] stage1_51;
   wire [303:0] stage1_52;
   wire [186:0] stage1_53;
   wire [262:0] stage1_54;
   wire [225:0] stage1_55;
   wire [256:0] stage1_56;
   wire [179:0] stage1_57;
   wire [242:0] stage1_58;
   wire [293:0] stage1_59;
   wire [199:0] stage1_60;
   wire [216:0] stage1_61;
   wire [372:0] stage1_62;
   wire [294:0] stage1_63;
   wire [111:0] stage1_64;
   wire [56:0] stage1_65;
   wire [33:0] stage2_0;
   wire [38:0] stage2_1;
   wire [72:0] stage2_2;
   wire [253:0] stage2_3;
   wire [92:0] stage2_4;
   wire [111:0] stage2_5;
   wire [120:0] stage2_6;
   wire [96:0] stage2_7;
   wire [172:0] stage2_8;
   wire [104:0] stage2_9;
   wire [133:0] stage2_10;
   wire [135:0] stage2_11;
   wire [127:0] stage2_12;
   wire [71:0] stage2_13;
   wire [114:0] stage2_14;
   wire [114:0] stage2_15;
   wire [109:0] stage2_16;
   wire [89:0] stage2_17;
   wire [161:0] stage2_18;
   wire [93:0] stage2_19;
   wire [87:0] stage2_20;
   wire [111:0] stage2_21;
   wire [109:0] stage2_22;
   wire [97:0] stage2_23;
   wire [84:0] stage2_24;
   wire [122:0] stage2_25;
   wire [130:0] stage2_26;
   wire [85:0] stage2_27;
   wire [79:0] stage2_28;
   wire [111:0] stage2_29;
   wire [99:0] stage2_30;
   wire [127:0] stage2_31;
   wire [117:0] stage2_32;
   wire [108:0] stage2_33;
   wire [127:0] stage2_34;
   wire [117:0] stage2_35;
   wire [119:0] stage2_36;
   wire [113:0] stage2_37;
   wire [99:0] stage2_38;
   wire [107:0] stage2_39;
   wire [139:0] stage2_40;
   wire [122:0] stage2_41;
   wire [81:0] stage2_42;
   wire [110:0] stage2_43;
   wire [137:0] stage2_44;
   wire [131:0] stage2_45;
   wire [92:0] stage2_46;
   wire [107:0] stage2_47;
   wire [153:0] stage2_48;
   wire [115:0] stage2_49;
   wire [152:0] stage2_50;
   wire [87:0] stage2_51;
   wire [127:0] stage2_52;
   wire [96:0] stage2_53;
   wire [123:0] stage2_54;
   wire [110:0] stage2_55;
   wire [131:0] stage2_56;
   wire [78:0] stage2_57;
   wire [84:0] stage2_58;
   wire [139:0] stage2_59;
   wire [110:0] stage2_60;
   wire [101:0] stage2_61;
   wire [144:0] stage2_62;
   wire [112:0] stage2_63;
   wire [101:0] stage2_64;
   wire [67:0] stage2_65;
   wire [53:0] stage2_66;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [14:0] stage3_2;
   wire [51:0] stage3_3;
   wire [59:0] stage3_4;
   wire [54:0] stage3_5;
   wire [66:0] stage3_6;
   wire [54:0] stage3_7;
   wire [46:0] stage3_8;
   wire [52:0] stage3_9;
   wire [67:0] stage3_10;
   wire [60:0] stage3_11;
   wire [80:0] stage3_12;
   wire [46:0] stage3_13;
   wire [34:0] stage3_14;
   wire [50:0] stage3_15;
   wire [58:0] stage3_16;
   wire [43:0] stage3_17;
   wire [63:0] stage3_18;
   wire [45:0] stage3_19;
   wire [57:0] stage3_20;
   wire [62:0] stage3_21;
   wire [49:0] stage3_22;
   wire [48:0] stage3_23;
   wire [34:0] stage3_24;
   wire [51:0] stage3_25;
   wire [51:0] stage3_26;
   wire [41:0] stage3_27;
   wire [69:0] stage3_28;
   wire [58:0] stage3_29;
   wire [38:0] stage3_30;
   wire [41:0] stage3_31;
   wire [55:0] stage3_32;
   wire [62:0] stage3_33;
   wire [44:0] stage3_34;
   wire [56:0] stage3_35;
   wire [55:0] stage3_36;
   wire [34:0] stage3_37;
   wire [68:0] stage3_38;
   wire [59:0] stage3_39;
   wire [45:0] stage3_40;
   wire [56:0] stage3_41;
   wire [53:0] stage3_42;
   wire [59:0] stage3_43;
   wire [84:0] stage3_44;
   wire [39:0] stage3_45;
   wire [48:0] stage3_46;
   wire [73:0] stage3_47;
   wire [36:0] stage3_48;
   wire [64:0] stage3_49;
   wire [63:0] stage3_50;
   wire [53:0] stage3_51;
   wire [55:0] stage3_52;
   wire [52:0] stage3_53;
   wire [62:0] stage3_54;
   wire [46:0] stage3_55;
   wire [38:0] stage3_56;
   wire [52:0] stage3_57;
   wire [48:0] stage3_58;
   wire [45:0] stage3_59;
   wire [52:0] stage3_60;
   wire [56:0] stage3_61;
   wire [40:0] stage3_62;
   wire [71:0] stage3_63;
   wire [50:0] stage3_64;
   wire [32:0] stage3_65;
   wire [53:0] stage3_66;
   wire [14:0] stage3_67;
   wire [4:0] stage3_68;
   wire [5:0] stage4_0;
   wire [6:0] stage4_1;
   wire [8:0] stage4_2;
   wire [21:0] stage4_3;
   wire [24:0] stage4_4;
   wire [46:0] stage4_5;
   wire [20:0] stage4_6;
   wire [39:0] stage4_7;
   wire [34:0] stage4_8;
   wire [13:0] stage4_9;
   wire [28:0] stage4_10;
   wire [33:0] stage4_11;
   wire [19:0] stage4_12;
   wire [27:0] stage4_13;
   wire [29:0] stage4_14;
   wire [22:0] stage4_15;
   wire [32:0] stage4_16;
   wire [22:0] stage4_17;
   wire [31:0] stage4_18;
   wire [19:0] stage4_19;
   wire [21:0] stage4_20;
   wire [26:0] stage4_21;
   wire [20:0] stage4_22;
   wire [23:0] stage4_23;
   wire [23:0] stage4_24;
   wire [19:0] stage4_25;
   wire [20:0] stage4_26;
   wire [20:0] stage4_27;
   wire [31:0] stage4_28;
   wire [23:0] stage4_29;
   wire [25:0] stage4_30;
   wire [16:0] stage4_31;
   wire [23:0] stage4_32;
   wire [33:0] stage4_33;
   wire [29:0] stage4_34;
   wire [23:0] stage4_35;
   wire [37:0] stage4_36;
   wire [15:0] stage4_37;
   wire [26:0] stage4_38;
   wire [22:0] stage4_39;
   wire [28:0] stage4_40;
   wire [23:0] stage4_41;
   wire [28:0] stage4_42;
   wire [22:0] stage4_43;
   wire [39:0] stage4_44;
   wire [25:0] stage4_45;
   wire [24:0] stage4_46;
   wire [25:0] stage4_47;
   wire [21:0] stage4_48;
   wire [27:0] stage4_49;
   wire [23:0] stage4_50;
   wire [26:0] stage4_51;
   wire [22:0] stage4_52;
   wire [28:0] stage4_53;
   wire [30:0] stage4_54;
   wire [28:0] stage4_55;
   wire [28:0] stage4_56;
   wire [24:0] stage4_57;
   wire [15:0] stage4_58;
   wire [15:0] stage4_59;
   wire [24:0] stage4_60;
   wire [28:0] stage4_61;
   wire [23:0] stage4_62;
   wire [17:0] stage4_63;
   wire [26:0] stage4_64;
   wire [22:0] stage4_65;
   wire [14:0] stage4_66;
   wire [16:0] stage4_67;
   wire [11:0] stage4_68;
   wire [2:0] stage4_69;
   wire [0:0] stage4_70;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [2:0] stage5_2;
   wire [7:0] stage5_3;
   wire [8:0] stage5_4;
   wire [20:0] stage5_5;
   wire [13:0] stage5_6;
   wire [10:0] stage5_7;
   wire [15:0] stage5_8;
   wire [12:0] stage5_9;
   wire [9:0] stage5_10;
   wire [19:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [14:0] stage5_14;
   wire [15:0] stage5_15;
   wire [13:0] stage5_16;
   wire [7:0] stage5_17;
   wire [13:0] stage5_18;
   wire [13:0] stage5_19;
   wire [7:0] stage5_20;
   wire [10:0] stage5_21;
   wire [14:0] stage5_22;
   wire [11:0] stage5_23;
   wire [8:0] stage5_24;
   wire [12:0] stage5_25;
   wire [16:0] stage5_26;
   wire [8:0] stage5_27;
   wire [11:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [11:0] stage5_31;
   wire [14:0] stage5_32;
   wire [8:0] stage5_33;
   wire [20:0] stage5_34;
   wire [8:0] stage5_35;
   wire [18:0] stage5_36;
   wire [10:0] stage5_37;
   wire [6:0] stage5_38;
   wire [10:0] stage5_39;
   wire [19:0] stage5_40;
   wire [8:0] stage5_41;
   wire [19:0] stage5_42;
   wire [7:0] stage5_43;
   wire [25:0] stage5_44;
   wire [9:0] stage5_45;
   wire [10:0] stage5_46;
   wire [12:0] stage5_47;
   wire [17:0] stage5_48;
   wire [16:0] stage5_49;
   wire [9:0] stage5_50;
   wire [9:0] stage5_51;
   wire [12:0] stage5_52;
   wire [11:0] stage5_53;
   wire [16:0] stage5_54;
   wire [17:0] stage5_55;
   wire [12:0] stage5_56;
   wire [8:0] stage5_57;
   wire [23:0] stage5_58;
   wire [5:0] stage5_59;
   wire [13:0] stage5_60;
   wire [9:0] stage5_61;
   wire [7:0] stage5_62;
   wire [10:0] stage5_63;
   wire [19:0] stage5_64;
   wire [5:0] stage5_65;
   wire [12:0] stage5_66;
   wire [7:0] stage5_67;
   wire [11:0] stage5_68;
   wire [2:0] stage5_69;
   wire [3:0] stage5_70;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [2:0] stage6_2;
   wire [3:0] stage6_3;
   wire [2:0] stage6_4;
   wire [6:0] stage6_5;
   wire [5:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [7:0] stage6_9;
   wire [4:0] stage6_10;
   wire [5:0] stage6_11;
   wire [7:0] stage6_12;
   wire [4:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [11:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [8:0] stage6_25;
   wire [4:0] stage6_26;
   wire [4:0] stage6_27;
   wire [3:0] stage6_28;
   wire [5:0] stage6_29;
   wire [7:0] stage6_30;
   wire [2:0] stage6_31;
   wire [5:0] stage6_32;
   wire [7:0] stage6_33;
   wire [5:0] stage6_34;
   wire [4:0] stage6_35;
   wire [7:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [4:0] stage6_39;
   wire [9:0] stage6_40;
   wire [10:0] stage6_41;
   wire [3:0] stage6_42;
   wire [4:0] stage6_43;
   wire [7:0] stage6_44;
   wire [6:0] stage6_45;
   wire [6:0] stage6_46;
   wire [3:0] stage6_47;
   wire [5:0] stage6_48;
   wire [9:0] stage6_49;
   wire [4:0] stage6_50;
   wire [4:0] stage6_51;
   wire [7:0] stage6_52;
   wire [3:0] stage6_53;
   wire [5:0] stage6_54;
   wire [5:0] stage6_55;
   wire [6:0] stage6_56;
   wire [6:0] stage6_57;
   wire [6:0] stage6_58;
   wire [4:0] stage6_59;
   wire [6:0] stage6_60;
   wire [5:0] stage6_61;
   wire [4:0] stage6_62;
   wire [2:0] stage6_63;
   wire [5:0] stage6_64;
   wire [9:0] stage6_65;
   wire [2:0] stage6_66;
   wire [4:0] stage6_67;
   wire [9:0] stage6_68;
   wire [2:0] stage6_69;
   wire [1:0] stage6_70;
   wire [1:0] stage6_71;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [2:0] stage7_2;
   wire [3:0] stage7_3;
   wire [0:0] stage7_4;
   wire [4:0] stage7_5;
   wire [1:0] stage7_6;
   wire [6:0] stage7_7;
   wire [0:0] stage7_8;
   wire [4:0] stage7_9;
   wire [3:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [6:0] stage7_13;
   wire [2:0] stage7_14;
   wire [1:0] stage7_15;
   wire [6:0] stage7_16;
   wire [2:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [0:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [6:0] stage7_23;
   wire [2:0] stage7_24;
   wire [5:0] stage7_25;
   wire [6:0] stage7_26;
   wire [0:0] stage7_27;
   wire [1:0] stage7_28;
   wire [2:0] stage7_29;
   wire [3:0] stage7_30;
   wire [1:0] stage7_31;
   wire [2:0] stage7_32;
   wire [2:0] stage7_33;
   wire [5:0] stage7_34;
   wire [6:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [2:0] stage7_38;
   wire [3:0] stage7_39;
   wire [1:0] stage7_40;
   wire [5:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [6:0] stage7_45;
   wire [6:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [5:0] stage7_49;
   wire [2:0] stage7_50;
   wire [5:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [4:0] stage7_54;
   wire [1:0] stage7_55;
   wire [5:0] stage7_56;
   wire [2:0] stage7_57;
   wire [1:0] stage7_58;
   wire [2:0] stage7_59;
   wire [4:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [4:0] stage7_63;
   wire [2:0] stage7_64;
   wire [11:0] stage7_65;
   wire [0:0] stage7_66;
   wire [0:0] stage7_67;
   wire [3:0] stage7_68;
   wire [2:0] stage7_69;
   wire [2:0] stage7_70;
   wire [2:0] stage7_71;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [1:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [0:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_2[7]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[8]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[9]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[10]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[11]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[12]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[13]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[14]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[15]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[16]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[17]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[18]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[19]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[20]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[21]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[22]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[23]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[24]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[25]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[26]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[27]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[28]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[29]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[30]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[31]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[32]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[33]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[34]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[35]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[36]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_2[37]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_2[38]},
      {stage0_3[31]},
      {stage1_4[31],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_2[39]},
      {stage0_3[32]},
      {stage1_4[32],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_2[40]},
      {stage0_3[33]},
      {stage1_4[33],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_2[41]},
      {stage0_3[34]},
      {stage1_4[34],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_2[42]},
      {stage0_3[35]},
      {stage1_4[35],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_2[43]},
      {stage0_3[36]},
      {stage1_4[36],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_2[44]},
      {stage0_3[37]},
      {stage1_4[37],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc1163_5 gpc45 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_2[45]},
      {stage0_3[38]},
      {stage1_4[38],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc1163_5 gpc46 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_2[46]},
      {stage0_3[39]},
      {stage1_4[39],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc1163_5 gpc47 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_2[47]},
      {stage0_3[40]},
      {stage1_4[40],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc1163_5 gpc48 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_2[48]},
      {stage0_3[41]},
      {stage1_4[41],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc1163_5 gpc49 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_2[49]},
      {stage0_3[42]},
      {stage1_4[42],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc1163_5 gpc50 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_2[50]},
      {stage0_3[43]},
      {stage1_4[43],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc1163_5 gpc51 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_2[51]},
      {stage0_3[44]},
      {stage1_4[44],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc1163_5 gpc52 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_2[52]},
      {stage0_3[45]},
      {stage1_4[45],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc1163_5 gpc53 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_2[53]},
      {stage0_3[46]},
      {stage1_4[46],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc1163_5 gpc54 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_2[54]},
      {stage0_3[47]},
      {stage1_4[47],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc1163_5 gpc55 (
      {stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_2[55]},
      {stage0_3[48]},
      {stage1_4[48],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc1163_5 gpc56 (
      {stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_2[56]},
      {stage0_3[49]},
      {stage1_4[49],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[50],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[51],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[52],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[53],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc615_5 gpc61 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_1[307]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[54],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc615_5 gpc62 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_1[308]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[55],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc615_5 gpc63 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_1[309]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[56],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc615_5 gpc64 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_1[310]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[57],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc615_5 gpc65 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247]},
      {stage0_1[311]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[58],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc615_5 gpc66 (
      {stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_1[312]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[59],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc615_5 gpc67 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_1[313]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[60],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc615_5 gpc68 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_1[314]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[61],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc615_5 gpc69 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_1[315]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[62],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc615_5 gpc70 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_1[316]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[63],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc615_5 gpc71 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277]},
      {stage0_1[317]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[64],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc615_5 gpc72 (
      {stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_1[318]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[65],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc615_5 gpc73 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_1[319]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[66],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc615_5 gpc74 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_1[320]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[67],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc615_5 gpc75 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_1[321]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[68],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc615_5 gpc76 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_1[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[69],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc615_5 gpc77 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307]},
      {stage0_1[323]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[70],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc615_5 gpc78 (
      {stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_1[324]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[71],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc615_5 gpc79 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_1[325]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[72],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc615_5 gpc80 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_1[326]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[73],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc615_5 gpc81 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_1[327]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[74],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc615_5 gpc82 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_1[328]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[75],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc615_5 gpc83 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337]},
      {stage0_1[329]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[76],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc615_5 gpc84 (
      {stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_1[330]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[77],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc615_5 gpc85 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_1[331]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[78],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc615_5 gpc86 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_1[332]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[79],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc615_5 gpc87 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_1[333]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[80],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc615_5 gpc88 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_1[334]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[81],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc615_5 gpc89 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367]},
      {stage0_1[335]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[82],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc615_5 gpc90 (
      {stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_1[336]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[83],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc615_5 gpc91 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_1[337]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[84],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc615_5 gpc92 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_1[338]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[85],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc615_5 gpc93 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_1[339]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[86],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc615_5 gpc94 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_1[340]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[87],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc615_5 gpc95 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397]},
      {stage0_1[341]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[88],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc615_5 gpc96 (
      {stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_1[342]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[89],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc615_5 gpc97 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_1[343]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[90],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc615_5 gpc98 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_1[344]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[91],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc615_5 gpc99 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_1[345]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[92],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc615_5 gpc100 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_1[346]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[93],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc615_5 gpc101 (
      {stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427]},
      {stage0_1[347]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[94],stage1_3[101],stage1_2[101],stage1_1[101],stage1_0[101]}
   );
   gpc615_5 gpc102 (
      {stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_1[348]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[95],stage1_3[102],stage1_2[102],stage1_1[102],stage1_0[102]}
   );
   gpc615_5 gpc103 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_1[349]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[96],stage1_3[103],stage1_2[103],stage1_1[103],stage1_0[103]}
   );
   gpc615_5 gpc104 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_1[350]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[97],stage1_3[104],stage1_2[104],stage1_1[104],stage1_0[104]}
   );
   gpc615_5 gpc105 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_1[351]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[98],stage1_3[105],stage1_2[105],stage1_1[105],stage1_0[105]}
   );
   gpc615_5 gpc106 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452]},
      {stage0_1[352]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[99],stage1_3[106],stage1_2[106],stage1_1[106],stage1_0[106]}
   );
   gpc615_5 gpc107 (
      {stage0_0[453], stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457]},
      {stage0_1[353]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[100],stage1_3[107],stage1_2[107],stage1_1[107],stage1_0[107]}
   );
   gpc615_5 gpc108 (
      {stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461], stage0_0[462]},
      {stage0_1[354]},
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage1_4[101],stage1_3[108],stage1_2[108],stage1_1[108],stage1_0[108]}
   );
   gpc615_5 gpc109 (
      {stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_1[355]},
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage1_4[102],stage1_3[109],stage1_2[109],stage1_1[109],stage1_0[109]}
   );
   gpc615_5 gpc110 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_1[356]},
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage1_4[103],stage1_3[110],stage1_2[110],stage1_1[110],stage1_0[110]}
   );
   gpc615_5 gpc111 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_1[357]},
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage1_4[104],stage1_3[111],stage1_2[111],stage1_1[111],stage1_0[111]}
   );
   gpc615_5 gpc112 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482]},
      {stage0_1[358]},
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage1_4[105],stage1_3[112],stage1_2[112],stage1_1[112],stage1_0[112]}
   );
   gpc615_5 gpc113 (
      {stage0_0[483], stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487]},
      {stage0_1[359]},
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage1_4[106],stage1_3[113],stage1_2[113],stage1_1[113],stage1_0[113]}
   );
   gpc615_5 gpc114 (
      {stage0_0[488], stage0_0[489], stage0_0[490], stage0_0[491], stage0_0[492]},
      {stage0_1[360]},
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage1_4[107],stage1_3[114],stage1_2[114],stage1_1[114],stage1_0[114]}
   );
   gpc615_5 gpc115 (
      {stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496], stage0_0[497]},
      {stage0_1[361]},
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage1_4[108],stage1_3[115],stage1_2[115],stage1_1[115],stage1_0[115]}
   );
   gpc615_5 gpc116 (
      {stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_1[362]},
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416]},
      {stage1_4[109],stage1_3[116],stage1_2[116],stage1_1[116],stage1_0[116]}
   );
   gpc615_5 gpc117 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507]},
      {stage0_1[363]},
      {stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage1_4[110],stage1_3[117],stage1_2[117],stage1_1[117],stage1_0[117]}
   );
   gpc615_5 gpc118 (
      {stage0_0[508], stage0_0[509], stage0_0[510], stage0_0[511], 1'b0},
      {stage0_1[364]},
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage1_4[111],stage1_3[118],stage1_2[118],stage1_1[118],stage1_0[118]}
   );
   gpc7_3 gpc119 (
      {stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc7_3 gpc120 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[0],stage1_4[112],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[1],stage1_4[113],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[2],stage1_4[114],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[3],stage1_4[115],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[4],stage1_4[116],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[5],stage1_4[117],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[6],stage1_4[118],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[7],stage1_4[119],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[8],stage1_4[120],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[9],stage1_4[121],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[10],stage1_4[122],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[11],stage1_4[123],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[12],stage1_4[124],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[13],stage1_4[125],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[14],stage1_4[126],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[15],stage1_4[127],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479], stage0_1[480]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[16],stage1_4[128],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc615_5 gpc138 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[17],stage1_4[129],stage1_3[138]}
   );
   gpc615_5 gpc139 (
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[18],stage1_4[130],stage1_3[139]}
   );
   gpc615_5 gpc140 (
      {stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[19],stage1_4[131],stage1_3[140]}
   );
   gpc615_5 gpc141 (
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[20],stage1_4[132],stage1_3[141]}
   );
   gpc615_5 gpc142 (
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[21],stage1_4[133],stage1_3[142]}
   );
   gpc615_5 gpc143 (
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181]},
      {stage0_4[5]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[5],stage1_5[22],stage1_4[134],stage1_3[143]}
   );
   gpc615_5 gpc144 (
      {stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage0_4[6]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[6],stage1_5[23],stage1_4[135],stage1_3[144]}
   );
   gpc615_5 gpc145 (
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191]},
      {stage0_4[7]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[7],stage1_5[24],stage1_4[136],stage1_3[145]}
   );
   gpc615_5 gpc146 (
      {stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage0_4[8]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[8],stage1_5[25],stage1_4[137],stage1_3[146]}
   );
   gpc615_5 gpc147 (
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage0_4[9]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[9],stage1_5[26],stage1_4[138],stage1_3[147]}
   );
   gpc615_5 gpc148 (
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage0_4[10]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[10],stage1_5[27],stage1_4[139],stage1_3[148]}
   );
   gpc615_5 gpc149 (
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211]},
      {stage0_4[11]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[11],stage1_5[28],stage1_4[140],stage1_3[149]}
   );
   gpc615_5 gpc150 (
      {stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage0_4[12]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[12],stage1_5[29],stage1_4[141],stage1_3[150]}
   );
   gpc615_5 gpc151 (
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221]},
      {stage0_4[13]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[13],stage1_5[30],stage1_4[142],stage1_3[151]}
   );
   gpc615_5 gpc152 (
      {stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage0_4[14]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[14],stage1_5[31],stage1_4[143],stage1_3[152]}
   );
   gpc615_5 gpc153 (
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage0_4[15]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[15],stage1_5[32],stage1_4[144],stage1_3[153]}
   );
   gpc615_5 gpc154 (
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage0_4[16]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[16],stage1_5[33],stage1_4[145],stage1_3[154]}
   );
   gpc615_5 gpc155 (
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241]},
      {stage0_4[17]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[17],stage1_5[34],stage1_4[146],stage1_3[155]}
   );
   gpc615_5 gpc156 (
      {stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage0_4[18]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[18],stage1_5[35],stage1_4[147],stage1_3[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251]},
      {stage0_4[19]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[19],stage1_5[36],stage1_4[148],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage0_4[20]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[20],stage1_5[37],stage1_4[149],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage0_4[21]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[21],stage1_5[38],stage1_4[150],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage0_4[22]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[22],stage1_5[39],stage1_4[151],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271]},
      {stage0_4[23]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[23],stage1_5[40],stage1_4[152],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage0_4[24]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[24],stage1_5[41],stage1_4[153],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281]},
      {stage0_4[25]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[25],stage1_5[42],stage1_4[154],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage0_4[26]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[26],stage1_5[43],stage1_4[155],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage0_4[27]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[27],stage1_5[44],stage1_4[156],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage0_4[28]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[28],stage1_5[45],stage1_4[157],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301]},
      {stage0_4[29]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[29],stage1_5[46],stage1_4[158],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage0_4[30]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[30],stage1_5[47],stage1_4[159],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311]},
      {stage0_4[31]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[31],stage1_5[48],stage1_4[160],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316]},
      {stage0_4[32]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[32],stage1_5[49],stage1_4[161],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage0_4[33]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[33],stage1_5[50],stage1_4[162],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage0_4[34]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[34],stage1_5[51],stage1_4[163],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331]},
      {stage0_4[35]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[35],stage1_5[52],stage1_4[164],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage0_4[36]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[36],stage1_5[53],stage1_4[165],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341]},
      {stage0_4[37]},
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage1_7[37],stage1_6[37],stage1_5[54],stage1_4[166],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346]},
      {stage0_4[38]},
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage1_7[38],stage1_6[38],stage1_5[55],stage1_4[167],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350], stage0_3[351]},
      {stage0_4[39]},
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage1_7[39],stage1_6[39],stage1_5[56],stage1_4[168],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage0_4[40]},
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage1_7[40],stage1_6[40],stage1_5[57],stage1_4[169],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361]},
      {stage0_4[41]},
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage1_7[41],stage1_6[41],stage1_5[58],stage1_4[170],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366]},
      {stage0_4[42]},
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage1_7[42],stage1_6[42],stage1_5[59],stage1_4[171],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370], stage0_3[371]},
      {stage0_4[43]},
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage1_7[43],stage1_6[43],stage1_5[60],stage1_4[172],stage1_3[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[44],stage1_6[44],stage1_5[61],stage1_4[173]}
   );
   gpc606_5 gpc183 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[45],stage1_6[45],stage1_5[62],stage1_4[174]}
   );
   gpc606_5 gpc184 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[46],stage1_6[46],stage1_5[63],stage1_4[175]}
   );
   gpc606_5 gpc185 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[47],stage1_6[47],stage1_5[64],stage1_4[176]}
   );
   gpc606_5 gpc186 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[48],stage1_6[48],stage1_5[65],stage1_4[177]}
   );
   gpc606_5 gpc187 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[49],stage1_6[49],stage1_5[66],stage1_4[178]}
   );
   gpc606_5 gpc188 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[50],stage1_6[50],stage1_5[67],stage1_4[179]}
   );
   gpc606_5 gpc189 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[51],stage1_6[51],stage1_5[68],stage1_4[180]}
   );
   gpc606_5 gpc190 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[52],stage1_6[52],stage1_5[69],stage1_4[181]}
   );
   gpc606_5 gpc191 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[53],stage1_6[53],stage1_5[70],stage1_4[182]}
   );
   gpc606_5 gpc192 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[54],stage1_6[54],stage1_5[71],stage1_4[183]}
   );
   gpc606_5 gpc193 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[55],stage1_6[55],stage1_5[72],stage1_4[184]}
   );
   gpc606_5 gpc194 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[56],stage1_6[56],stage1_5[73],stage1_4[185]}
   );
   gpc606_5 gpc195 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[57],stage1_6[57],stage1_5[74],stage1_4[186]}
   );
   gpc606_5 gpc196 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[58],stage1_6[58],stage1_5[75],stage1_4[187]}
   );
   gpc606_5 gpc197 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[59],stage1_6[59],stage1_5[76],stage1_4[188]}
   );
   gpc606_5 gpc198 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[60],stage1_6[60],stage1_5[77],stage1_4[189]}
   );
   gpc606_5 gpc199 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[61],stage1_6[61],stage1_5[78],stage1_4[190]}
   );
   gpc606_5 gpc200 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[62],stage1_6[62],stage1_5[79],stage1_4[191]}
   );
   gpc606_5 gpc201 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[63],stage1_6[63],stage1_5[80],stage1_4[192]}
   );
   gpc606_5 gpc202 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[64],stage1_6[64],stage1_5[81],stage1_4[193]}
   );
   gpc606_5 gpc203 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[65],stage1_6[65],stage1_5[82],stage1_4[194]}
   );
   gpc606_5 gpc204 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[66],stage1_6[66],stage1_5[83],stage1_4[195]}
   );
   gpc606_5 gpc205 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[67],stage1_6[67],stage1_5[84],stage1_4[196]}
   );
   gpc606_5 gpc206 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[68],stage1_6[68],stage1_5[85],stage1_4[197]}
   );
   gpc606_5 gpc207 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[69],stage1_6[69],stage1_5[86],stage1_4[198]}
   );
   gpc606_5 gpc208 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[70],stage1_6[70],stage1_5[87],stage1_4[199]}
   );
   gpc606_5 gpc209 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[71],stage1_6[71],stage1_5[88],stage1_4[200]}
   );
   gpc606_5 gpc210 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[72],stage1_6[72],stage1_5[89],stage1_4[201]}
   );
   gpc606_5 gpc211 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[73],stage1_6[73],stage1_5[90],stage1_4[202]}
   );
   gpc606_5 gpc212 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[74],stage1_6[74],stage1_5[91],stage1_4[203]}
   );
   gpc606_5 gpc213 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[75],stage1_6[75],stage1_5[92],stage1_4[204]}
   );
   gpc606_5 gpc214 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[76],stage1_6[76],stage1_5[93],stage1_4[205]}
   );
   gpc606_5 gpc215 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[77],stage1_6[77],stage1_5[94],stage1_4[206]}
   );
   gpc606_5 gpc216 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[78],stage1_6[78],stage1_5[95],stage1_4[207]}
   );
   gpc606_5 gpc217 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[79],stage1_6[79],stage1_5[96],stage1_4[208]}
   );
   gpc606_5 gpc218 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[80],stage1_6[80],stage1_5[97],stage1_4[209]}
   );
   gpc606_5 gpc219 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[81],stage1_6[81],stage1_5[98],stage1_4[210]}
   );
   gpc606_5 gpc220 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[82],stage1_6[82],stage1_5[99],stage1_4[211]}
   );
   gpc606_5 gpc221 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[83],stage1_6[83],stage1_5[100],stage1_4[212]}
   );
   gpc606_5 gpc222 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[84],stage1_6[84],stage1_5[101],stage1_4[213]}
   );
   gpc606_5 gpc223 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[85],stage1_6[85],stage1_5[102],stage1_4[214]}
   );
   gpc606_5 gpc224 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[86],stage1_6[86],stage1_5[103],stage1_4[215]}
   );
   gpc606_5 gpc225 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[87],stage1_6[87],stage1_5[104],stage1_4[216]}
   );
   gpc606_5 gpc226 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[88],stage1_6[88],stage1_5[105],stage1_4[217]}
   );
   gpc606_5 gpc227 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[89],stage1_6[89],stage1_5[106],stage1_4[218]}
   );
   gpc606_5 gpc228 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[90],stage1_6[90],stage1_5[107],stage1_4[219]}
   );
   gpc606_5 gpc229 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[91],stage1_6[91],stage1_5[108],stage1_4[220]}
   );
   gpc606_5 gpc230 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[92],stage1_6[92],stage1_5[109],stage1_4[221]}
   );
   gpc606_5 gpc231 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[93],stage1_6[93],stage1_5[110],stage1_4[222]}
   );
   gpc606_5 gpc232 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[94],stage1_6[94],stage1_5[111],stage1_4[223]}
   );
   gpc606_5 gpc233 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[95],stage1_6[95],stage1_5[112],stage1_4[224]}
   );
   gpc606_5 gpc234 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[96],stage1_6[96],stage1_5[113],stage1_4[225]}
   );
   gpc606_5 gpc235 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[97],stage1_6[97],stage1_5[114],stage1_4[226]}
   );
   gpc606_5 gpc236 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[98],stage1_6[98],stage1_5[115],stage1_4[227]}
   );
   gpc606_5 gpc237 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[99],stage1_6[99],stage1_5[116],stage1_4[228]}
   );
   gpc606_5 gpc238 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[100],stage1_6[100],stage1_5[117],stage1_4[229]}
   );
   gpc606_5 gpc239 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[101],stage1_6[101],stage1_5[118],stage1_4[230]}
   );
   gpc606_5 gpc240 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[102],stage1_6[102],stage1_5[119],stage1_4[231]}
   );
   gpc606_5 gpc241 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[103],stage1_6[103],stage1_5[120],stage1_4[232]}
   );
   gpc606_5 gpc242 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[104],stage1_6[104],stage1_5[121],stage1_4[233]}
   );
   gpc606_5 gpc243 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[105],stage1_6[105],stage1_5[122],stage1_4[234]}
   );
   gpc606_5 gpc244 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[106],stage1_6[106],stage1_5[123],stage1_4[235]}
   );
   gpc606_5 gpc245 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[107],stage1_6[107],stage1_5[124],stage1_4[236]}
   );
   gpc606_5 gpc246 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[108],stage1_6[108],stage1_5[125],stage1_4[237]}
   );
   gpc606_5 gpc247 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[109],stage1_6[109],stage1_5[126],stage1_4[238]}
   );
   gpc606_5 gpc248 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[110],stage1_6[110],stage1_5[127],stage1_4[239]}
   );
   gpc606_5 gpc249 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[111],stage1_6[111],stage1_5[128],stage1_4[240]}
   );
   gpc606_5 gpc250 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[112],stage1_6[112],stage1_5[129],stage1_4[241]}
   );
   gpc606_5 gpc251 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[113],stage1_6[113],stage1_5[130],stage1_4[242]}
   );
   gpc606_5 gpc252 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[114],stage1_6[114],stage1_5[131],stage1_4[243]}
   );
   gpc606_5 gpc253 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[115],stage1_6[115],stage1_5[132],stage1_4[244]}
   );
   gpc606_5 gpc254 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[116],stage1_6[116],stage1_5[133],stage1_4[245]}
   );
   gpc606_5 gpc255 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486], stage0_4[487]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[117],stage1_6[117],stage1_5[134],stage1_4[246]}
   );
   gpc606_5 gpc256 (
      {stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491], stage0_4[492], stage0_4[493]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[118],stage1_6[118],stage1_5[135],stage1_4[247]}
   );
   gpc606_5 gpc257 (
      {stage0_4[494], stage0_4[495], stage0_4[496], stage0_4[497], stage0_4[498], stage0_4[499]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[119],stage1_6[119],stage1_5[136],stage1_4[248]}
   );
   gpc606_5 gpc258 (
      {stage0_4[500], stage0_4[501], stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[120],stage1_6[120],stage1_5[137],stage1_4[249]}
   );
   gpc606_5 gpc259 (
      {stage0_4[506], stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage1_8[77],stage1_7[121],stage1_6[121],stage1_5[138],stage1_4[250]}
   );
   gpc606_5 gpc260 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[78],stage1_7[122],stage1_6[122],stage1_5[139]}
   );
   gpc606_5 gpc261 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[79],stage1_7[123],stage1_6[123],stage1_5[140]}
   );
   gpc606_5 gpc262 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[80],stage1_7[124],stage1_6[124],stage1_5[141]}
   );
   gpc606_5 gpc263 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[81],stage1_7[125],stage1_6[125],stage1_5[142]}
   );
   gpc606_5 gpc264 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[82],stage1_7[126],stage1_6[126],stage1_5[143]}
   );
   gpc606_5 gpc265 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[83],stage1_7[127],stage1_6[127],stage1_5[144]}
   );
   gpc606_5 gpc266 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[84],stage1_7[128],stage1_6[128],stage1_5[145]}
   );
   gpc606_5 gpc267 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[85],stage1_7[129],stage1_6[129],stage1_5[146]}
   );
   gpc606_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[86],stage1_7[130],stage1_6[130],stage1_5[147]}
   );
   gpc606_5 gpc269 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[87],stage1_7[131],stage1_6[131],stage1_5[148]}
   );
   gpc606_5 gpc270 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[88],stage1_7[132],stage1_6[132],stage1_5[149]}
   );
   gpc606_5 gpc271 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[89],stage1_7[133],stage1_6[133],stage1_5[150]}
   );
   gpc606_5 gpc272 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[90],stage1_7[134],stage1_6[134],stage1_5[151]}
   );
   gpc606_5 gpc273 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[91],stage1_7[135],stage1_6[135],stage1_5[152]}
   );
   gpc606_5 gpc274 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[92],stage1_7[136],stage1_6[136],stage1_5[153]}
   );
   gpc606_5 gpc275 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[93],stage1_7[137],stage1_6[137],stage1_5[154]}
   );
   gpc606_5 gpc276 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[94],stage1_7[138],stage1_6[138],stage1_5[155]}
   );
   gpc606_5 gpc277 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[95],stage1_7[139],stage1_6[139],stage1_5[156]}
   );
   gpc606_5 gpc278 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[96],stage1_7[140],stage1_6[140],stage1_5[157]}
   );
   gpc606_5 gpc279 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[97],stage1_7[141],stage1_6[141],stage1_5[158]}
   );
   gpc606_5 gpc280 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[98],stage1_7[142],stage1_6[142],stage1_5[159]}
   );
   gpc606_5 gpc281 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[99],stage1_7[143],stage1_6[143],stage1_5[160]}
   );
   gpc606_5 gpc282 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[100],stage1_7[144],stage1_6[144],stage1_5[161]}
   );
   gpc606_5 gpc283 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[101],stage1_7[145],stage1_6[145],stage1_5[162]}
   );
   gpc606_5 gpc284 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[102],stage1_7[146],stage1_6[146],stage1_5[163]}
   );
   gpc606_5 gpc285 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[103],stage1_7[147],stage1_6[147],stage1_5[164]}
   );
   gpc606_5 gpc286 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[104],stage1_7[148],stage1_6[148],stage1_5[165]}
   );
   gpc606_5 gpc287 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[105],stage1_7[149],stage1_6[149],stage1_5[166]}
   );
   gpc606_5 gpc288 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[106],stage1_7[150],stage1_6[150],stage1_5[167]}
   );
   gpc606_5 gpc289 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[107],stage1_7[151],stage1_6[151],stage1_5[168]}
   );
   gpc606_5 gpc290 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[108],stage1_7[152],stage1_6[152],stage1_5[169]}
   );
   gpc606_5 gpc291 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[109],stage1_7[153],stage1_6[153],stage1_5[170]}
   );
   gpc606_5 gpc292 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[110],stage1_7[154],stage1_6[154],stage1_5[171]}
   );
   gpc606_5 gpc293 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[111],stage1_7[155],stage1_6[155],stage1_5[172]}
   );
   gpc615_5 gpc294 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472]},
      {stage0_7[204]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[34],stage1_8[112],stage1_7[156],stage1_6[156]}
   );
   gpc615_5 gpc295 (
      {stage0_6[473], stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477]},
      {stage0_7[205]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[35],stage1_8[113],stage1_7[157],stage1_6[157]}
   );
   gpc615_5 gpc296 (
      {stage0_6[478], stage0_6[479], stage0_6[480], stage0_6[481], stage0_6[482]},
      {stage0_7[206]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[36],stage1_8[114],stage1_7[158],stage1_6[158]}
   );
   gpc615_5 gpc297 (
      {stage0_6[483], stage0_6[484], stage0_6[485], stage0_6[486], stage0_6[487]},
      {stage0_7[207]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[37],stage1_8[115],stage1_7[159],stage1_6[159]}
   );
   gpc615_5 gpc298 (
      {stage0_6[488], stage0_6[489], stage0_6[490], stage0_6[491], stage0_6[492]},
      {stage0_7[208]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[38],stage1_8[116],stage1_7[160],stage1_6[160]}
   );
   gpc615_5 gpc299 (
      {stage0_7[209], stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[39],stage1_8[117],stage1_7[161]}
   );
   gpc615_5 gpc300 (
      {stage0_7[214], stage0_7[215], stage0_7[216], stage0_7[217], stage0_7[218]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[40],stage1_8[118],stage1_7[162]}
   );
   gpc615_5 gpc301 (
      {stage0_7[219], stage0_7[220], stage0_7[221], stage0_7[222], stage0_7[223]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[41],stage1_8[119],stage1_7[163]}
   );
   gpc615_5 gpc302 (
      {stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227], stage0_7[228]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[42],stage1_8[120],stage1_7[164]}
   );
   gpc615_5 gpc303 (
      {stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[43],stage1_8[121],stage1_7[165]}
   );
   gpc615_5 gpc304 (
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[44],stage1_8[122],stage1_7[166]}
   );
   gpc615_5 gpc305 (
      {stage0_7[239], stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[45],stage1_8[123],stage1_7[167]}
   );
   gpc615_5 gpc306 (
      {stage0_7[244], stage0_7[245], stage0_7[246], stage0_7[247], stage0_7[248]},
      {stage0_8[37]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[12],stage1_9[46],stage1_8[124],stage1_7[168]}
   );
   gpc615_5 gpc307 (
      {stage0_7[249], stage0_7[250], stage0_7[251], stage0_7[252], stage0_7[253]},
      {stage0_8[38]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[13],stage1_9[47],stage1_8[125],stage1_7[169]}
   );
   gpc615_5 gpc308 (
      {stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257], stage0_7[258]},
      {stage0_8[39]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[14],stage1_9[48],stage1_8[126],stage1_7[170]}
   );
   gpc615_5 gpc309 (
      {stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage0_8[40]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[15],stage1_9[49],stage1_8[127],stage1_7[171]}
   );
   gpc615_5 gpc310 (
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268]},
      {stage0_8[41]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[16],stage1_9[50],stage1_8[128],stage1_7[172]}
   );
   gpc615_5 gpc311 (
      {stage0_7[269], stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273]},
      {stage0_8[42]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[17],stage1_9[51],stage1_8[129],stage1_7[173]}
   );
   gpc615_5 gpc312 (
      {stage0_7[274], stage0_7[275], stage0_7[276], stage0_7[277], stage0_7[278]},
      {stage0_8[43]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[18],stage1_9[52],stage1_8[130],stage1_7[174]}
   );
   gpc615_5 gpc313 (
      {stage0_7[279], stage0_7[280], stage0_7[281], stage0_7[282], stage0_7[283]},
      {stage0_8[44]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[19],stage1_9[53],stage1_8[131],stage1_7[175]}
   );
   gpc615_5 gpc314 (
      {stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287], stage0_7[288]},
      {stage0_8[45]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[20],stage1_9[54],stage1_8[132],stage1_7[176]}
   );
   gpc615_5 gpc315 (
      {stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage0_8[46]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[21],stage1_9[55],stage1_8[133],stage1_7[177]}
   );
   gpc615_5 gpc316 (
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298]},
      {stage0_8[47]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[22],stage1_9[56],stage1_8[134],stage1_7[178]}
   );
   gpc615_5 gpc317 (
      {stage0_7[299], stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303]},
      {stage0_8[48]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[23],stage1_9[57],stage1_8[135],stage1_7[179]}
   );
   gpc615_5 gpc318 (
      {stage0_7[304], stage0_7[305], stage0_7[306], stage0_7[307], stage0_7[308]},
      {stage0_8[49]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[24],stage1_9[58],stage1_8[136],stage1_7[180]}
   );
   gpc615_5 gpc319 (
      {stage0_7[309], stage0_7[310], stage0_7[311], stage0_7[312], stage0_7[313]},
      {stage0_8[50]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[25],stage1_9[59],stage1_8[137],stage1_7[181]}
   );
   gpc615_5 gpc320 (
      {stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317], stage0_7[318]},
      {stage0_8[51]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[26],stage1_9[60],stage1_8[138],stage1_7[182]}
   );
   gpc615_5 gpc321 (
      {stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage0_8[52]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[27],stage1_9[61],stage1_8[139],stage1_7[183]}
   );
   gpc615_5 gpc322 (
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328]},
      {stage0_8[53]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[28],stage1_9[62],stage1_8[140],stage1_7[184]}
   );
   gpc615_5 gpc323 (
      {stage0_7[329], stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333]},
      {stage0_8[54]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[29],stage1_9[63],stage1_8[141],stage1_7[185]}
   );
   gpc615_5 gpc324 (
      {stage0_7[334], stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338]},
      {stage0_8[55]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[30],stage1_9[64],stage1_8[142],stage1_7[186]}
   );
   gpc615_5 gpc325 (
      {stage0_7[339], stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343]},
      {stage0_8[56]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[31],stage1_9[65],stage1_8[143],stage1_7[187]}
   );
   gpc615_5 gpc326 (
      {stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348]},
      {stage0_8[57]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[32],stage1_9[66],stage1_8[144],stage1_7[188]}
   );
   gpc615_5 gpc327 (
      {stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage0_8[58]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[33],stage1_9[67],stage1_8[145],stage1_7[189]}
   );
   gpc615_5 gpc328 (
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358]},
      {stage0_8[59]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[34],stage1_9[68],stage1_8[146],stage1_7[190]}
   );
   gpc615_5 gpc329 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363]},
      {stage0_8[60]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[35],stage1_9[69],stage1_8[147],stage1_7[191]}
   );
   gpc606_5 gpc330 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[31],stage1_10[36],stage1_9[70],stage1_8[148]}
   );
   gpc606_5 gpc331 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[32],stage1_10[37],stage1_9[71],stage1_8[149]}
   );
   gpc606_5 gpc332 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[33],stage1_10[38],stage1_9[72],stage1_8[150]}
   );
   gpc606_5 gpc333 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[34],stage1_10[39],stage1_9[73],stage1_8[151]}
   );
   gpc606_5 gpc334 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[35],stage1_10[40],stage1_9[74],stage1_8[152]}
   );
   gpc606_5 gpc335 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[36],stage1_10[41],stage1_9[75],stage1_8[153]}
   );
   gpc606_5 gpc336 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[37],stage1_10[42],stage1_9[76],stage1_8[154]}
   );
   gpc606_5 gpc337 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[38],stage1_10[43],stage1_9[77],stage1_8[155]}
   );
   gpc606_5 gpc338 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[39],stage1_10[44],stage1_9[78],stage1_8[156]}
   );
   gpc606_5 gpc339 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[40],stage1_10[45],stage1_9[79],stage1_8[157]}
   );
   gpc606_5 gpc340 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[41],stage1_10[46],stage1_9[80],stage1_8[158]}
   );
   gpc606_5 gpc341 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[42],stage1_10[47],stage1_9[81],stage1_8[159]}
   );
   gpc606_5 gpc342 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[43],stage1_10[48],stage1_9[82],stage1_8[160]}
   );
   gpc606_5 gpc343 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[44],stage1_10[49],stage1_9[83],stage1_8[161]}
   );
   gpc606_5 gpc344 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[45],stage1_10[50],stage1_9[84],stage1_8[162]}
   );
   gpc606_5 gpc345 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[46],stage1_10[51],stage1_9[85],stage1_8[163]}
   );
   gpc606_5 gpc346 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[47],stage1_10[52],stage1_9[86],stage1_8[164]}
   );
   gpc606_5 gpc347 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[48],stage1_10[53],stage1_9[87],stage1_8[165]}
   );
   gpc606_5 gpc348 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[49],stage1_10[54],stage1_9[88],stage1_8[166]}
   );
   gpc606_5 gpc349 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[50],stage1_10[55],stage1_9[89],stage1_8[167]}
   );
   gpc606_5 gpc350 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[51],stage1_10[56],stage1_9[90],stage1_8[168]}
   );
   gpc606_5 gpc351 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[52],stage1_10[57],stage1_9[91],stage1_8[169]}
   );
   gpc606_5 gpc352 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[53],stage1_10[58],stage1_9[92],stage1_8[170]}
   );
   gpc606_5 gpc353 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[54],stage1_10[59],stage1_9[93],stage1_8[171]}
   );
   gpc606_5 gpc354 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[55],stage1_10[60],stage1_9[94],stage1_8[172]}
   );
   gpc606_5 gpc355 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[56],stage1_10[61],stage1_9[95],stage1_8[173]}
   );
   gpc606_5 gpc356 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[57],stage1_10[62],stage1_9[96],stage1_8[174]}
   );
   gpc606_5 gpc357 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[58],stage1_10[63],stage1_9[97],stage1_8[175]}
   );
   gpc606_5 gpc358 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[59],stage1_10[64],stage1_9[98],stage1_8[176]}
   );
   gpc606_5 gpc359 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[60],stage1_10[65],stage1_9[99],stage1_8[177]}
   );
   gpc606_5 gpc360 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[61],stage1_10[66],stage1_9[100],stage1_8[178]}
   );
   gpc606_5 gpc361 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[62],stage1_10[67],stage1_9[101],stage1_8[179]}
   );
   gpc606_5 gpc362 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[63],stage1_10[68],stage1_9[102],stage1_8[180]}
   );
   gpc606_5 gpc363 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[64],stage1_10[69],stage1_9[103],stage1_8[181]}
   );
   gpc606_5 gpc364 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[65],stage1_10[70],stage1_9[104],stage1_8[182]}
   );
   gpc606_5 gpc365 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[66],stage1_10[71],stage1_9[105],stage1_8[183]}
   );
   gpc606_5 gpc366 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[67],stage1_10[72],stage1_9[106],stage1_8[184]}
   );
   gpc606_5 gpc367 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[68],stage1_10[73],stage1_9[107],stage1_8[185]}
   );
   gpc606_5 gpc368 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[69],stage1_10[74],stage1_9[108],stage1_8[186]}
   );
   gpc606_5 gpc369 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[70],stage1_10[75],stage1_9[109],stage1_8[187]}
   );
   gpc606_5 gpc370 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[71],stage1_10[76],stage1_9[110],stage1_8[188]}
   );
   gpc606_5 gpc371 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[72],stage1_10[77],stage1_9[111],stage1_8[189]}
   );
   gpc606_5 gpc372 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[73],stage1_10[78],stage1_9[112],stage1_8[190]}
   );
   gpc606_5 gpc373 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[74],stage1_10[79],stage1_9[113],stage1_8[191]}
   );
   gpc606_5 gpc374 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[75],stage1_10[80],stage1_9[114],stage1_8[192]}
   );
   gpc606_5 gpc375 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[76],stage1_10[81],stage1_9[115],stage1_8[193]}
   );
   gpc606_5 gpc376 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[77],stage1_10[82],stage1_9[116],stage1_8[194]}
   );
   gpc606_5 gpc377 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[78],stage1_10[83],stage1_9[117],stage1_8[195]}
   );
   gpc606_5 gpc378 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[79],stage1_10[84],stage1_9[118],stage1_8[196]}
   );
   gpc606_5 gpc379 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[80],stage1_10[85],stage1_9[119],stage1_8[197]}
   );
   gpc606_5 gpc380 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[81],stage1_10[86],stage1_9[120],stage1_8[198]}
   );
   gpc606_5 gpc381 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[82],stage1_10[87],stage1_9[121],stage1_8[199]}
   );
   gpc606_5 gpc382 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[83],stage1_10[88],stage1_9[122],stage1_8[200]}
   );
   gpc606_5 gpc383 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[84],stage1_10[89],stage1_9[123],stage1_8[201]}
   );
   gpc606_5 gpc384 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[85],stage1_10[90],stage1_9[124],stage1_8[202]}
   );
   gpc606_5 gpc385 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[86],stage1_10[91],stage1_9[125],stage1_8[203]}
   );
   gpc606_5 gpc386 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[87],stage1_10[92],stage1_9[126],stage1_8[204]}
   );
   gpc606_5 gpc387 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[88],stage1_10[93],stage1_9[127],stage1_8[205]}
   );
   gpc606_5 gpc388 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[89],stage1_10[94],stage1_9[128],stage1_8[206]}
   );
   gpc606_5 gpc389 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[90],stage1_10[95],stage1_9[129],stage1_8[207]}
   );
   gpc606_5 gpc390 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[91],stage1_10[96],stage1_9[130],stage1_8[208]}
   );
   gpc606_5 gpc391 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[92],stage1_10[97],stage1_9[131],stage1_8[209]}
   );
   gpc606_5 gpc392 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[93],stage1_10[98],stage1_9[132],stage1_8[210]}
   );
   gpc606_5 gpc393 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[94],stage1_10[99],stage1_9[133],stage1_8[211]}
   );
   gpc606_5 gpc394 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[95],stage1_10[100],stage1_9[134],stage1_8[212]}
   );
   gpc606_5 gpc395 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[96],stage1_10[101],stage1_9[135],stage1_8[213]}
   );
   gpc606_5 gpc396 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[97],stage1_10[102],stage1_9[136],stage1_8[214]}
   );
   gpc606_5 gpc397 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[98],stage1_10[103],stage1_9[137],stage1_8[215]}
   );
   gpc606_5 gpc398 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[99],stage1_10[104],stage1_9[138],stage1_8[216]}
   );
   gpc606_5 gpc399 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[100],stage1_10[105],stage1_9[139],stage1_8[217]}
   );
   gpc606_5 gpc400 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[101],stage1_10[106],stage1_9[140],stage1_8[218]}
   );
   gpc606_5 gpc401 (
      {stage0_8[487], stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[102],stage1_10[107],stage1_9[141],stage1_8[219]}
   );
   gpc606_5 gpc402 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[72],stage1_11[103],stage1_10[108],stage1_9[142]}
   );
   gpc606_5 gpc403 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[73],stage1_11[104],stage1_10[109],stage1_9[143]}
   );
   gpc606_5 gpc404 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[74],stage1_11[105],stage1_10[110],stage1_9[144]}
   );
   gpc606_5 gpc405 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[75],stage1_11[106],stage1_10[111],stage1_9[145]}
   );
   gpc606_5 gpc406 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[76],stage1_11[107],stage1_10[112],stage1_9[146]}
   );
   gpc606_5 gpc407 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[77],stage1_11[108],stage1_10[113],stage1_9[147]}
   );
   gpc606_5 gpc408 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[78],stage1_11[109],stage1_10[114],stage1_9[148]}
   );
   gpc606_5 gpc409 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[79],stage1_11[110],stage1_10[115],stage1_9[149]}
   );
   gpc606_5 gpc410 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[80],stage1_11[111],stage1_10[116],stage1_9[150]}
   );
   gpc606_5 gpc411 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[81],stage1_11[112],stage1_10[117],stage1_9[151]}
   );
   gpc606_5 gpc412 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[82],stage1_11[113],stage1_10[118],stage1_9[152]}
   );
   gpc606_5 gpc413 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[83],stage1_11[114],stage1_10[119],stage1_9[153]}
   );
   gpc606_5 gpc414 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[84],stage1_11[115],stage1_10[120],stage1_9[154]}
   );
   gpc606_5 gpc415 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[85],stage1_11[116],stage1_10[121],stage1_9[155]}
   );
   gpc606_5 gpc416 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[86],stage1_11[117],stage1_10[122],stage1_9[156]}
   );
   gpc606_5 gpc417 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[87],stage1_11[118],stage1_10[123],stage1_9[157]}
   );
   gpc606_5 gpc418 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[88],stage1_11[119],stage1_10[124],stage1_9[158]}
   );
   gpc606_5 gpc419 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[89],stage1_11[120],stage1_10[125],stage1_9[159]}
   );
   gpc606_5 gpc420 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[90],stage1_11[121],stage1_10[126],stage1_9[160]}
   );
   gpc606_5 gpc421 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[91],stage1_11[122],stage1_10[127],stage1_9[161]}
   );
   gpc606_5 gpc422 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[92],stage1_11[123],stage1_10[128],stage1_9[162]}
   );
   gpc615_5 gpc423 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[126]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[21],stage1_12[93],stage1_11[124],stage1_10[129]}
   );
   gpc615_5 gpc424 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[127]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[22],stage1_12[94],stage1_11[125],stage1_10[130]}
   );
   gpc615_5 gpc425 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[128]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[23],stage1_12[95],stage1_11[126],stage1_10[131]}
   );
   gpc615_5 gpc426 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[129]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[24],stage1_12[96],stage1_11[127],stage1_10[132]}
   );
   gpc615_5 gpc427 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[130]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[25],stage1_12[97],stage1_11[128],stage1_10[133]}
   );
   gpc615_5 gpc428 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[131]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[26],stage1_12[98],stage1_11[129],stage1_10[134]}
   );
   gpc615_5 gpc429 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[132]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[27],stage1_12[99],stage1_11[130],stage1_10[135]}
   );
   gpc615_5 gpc430 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[133]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[28],stage1_12[100],stage1_11[131],stage1_10[136]}
   );
   gpc615_5 gpc431 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[134]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[29],stage1_12[101],stage1_11[132],stage1_10[137]}
   );
   gpc615_5 gpc432 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[135]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[30],stage1_12[102],stage1_11[133],stage1_10[138]}
   );
   gpc615_5 gpc433 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[136]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[31],stage1_12[103],stage1_11[134],stage1_10[139]}
   );
   gpc615_5 gpc434 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[137]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[32],stage1_12[104],stage1_11[135],stage1_10[140]}
   );
   gpc615_5 gpc435 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[138]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[33],stage1_12[105],stage1_11[136],stage1_10[141]}
   );
   gpc615_5 gpc436 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[139]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[34],stage1_12[106],stage1_11[137],stage1_10[142]}
   );
   gpc615_5 gpc437 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[84]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[14],stage1_13[35],stage1_12[107],stage1_11[138]}
   );
   gpc615_5 gpc438 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[85]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[15],stage1_13[36],stage1_12[108],stage1_11[139]}
   );
   gpc615_5 gpc439 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[86]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[16],stage1_13[37],stage1_12[109],stage1_11[140]}
   );
   gpc615_5 gpc440 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[87]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[17],stage1_13[38],stage1_12[110],stage1_11[141]}
   );
   gpc615_5 gpc441 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[88]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[18],stage1_13[39],stage1_12[111],stage1_11[142]}
   );
   gpc615_5 gpc442 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[89]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[19],stage1_13[40],stage1_12[112],stage1_11[143]}
   );
   gpc615_5 gpc443 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[90]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[20],stage1_13[41],stage1_12[113],stage1_11[144]}
   );
   gpc615_5 gpc444 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[91]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[21],stage1_13[42],stage1_12[114],stage1_11[145]}
   );
   gpc615_5 gpc445 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[92]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[22],stage1_13[43],stage1_12[115],stage1_11[146]}
   );
   gpc615_5 gpc446 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[93]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[23],stage1_13[44],stage1_12[116],stage1_11[147]}
   );
   gpc615_5 gpc447 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[94]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[24],stage1_13[45],stage1_12[117],stage1_11[148]}
   );
   gpc615_5 gpc448 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[95]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[25],stage1_13[46],stage1_12[118],stage1_11[149]}
   );
   gpc615_5 gpc449 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[96]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[26],stage1_13[47],stage1_12[119],stage1_11[150]}
   );
   gpc615_5 gpc450 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[97]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[27],stage1_13[48],stage1_12[120],stage1_11[151]}
   );
   gpc615_5 gpc451 (
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214]},
      {stage0_12[98]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[28],stage1_13[49],stage1_12[121],stage1_11[152]}
   );
   gpc615_5 gpc452 (
      {stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage0_12[99]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[29],stage1_13[50],stage1_12[122],stage1_11[153]}
   );
   gpc615_5 gpc453 (
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224]},
      {stage0_12[100]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[30],stage1_13[51],stage1_12[123],stage1_11[154]}
   );
   gpc615_5 gpc454 (
      {stage0_11[225], stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229]},
      {stage0_12[101]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[31],stage1_13[52],stage1_12[124],stage1_11[155]}
   );
   gpc615_5 gpc455 (
      {stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233], stage0_11[234]},
      {stage0_12[102]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[32],stage1_13[53],stage1_12[125],stage1_11[156]}
   );
   gpc615_5 gpc456 (
      {stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage0_12[103]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[33],stage1_13[54],stage1_12[126],stage1_11[157]}
   );
   gpc615_5 gpc457 (
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244]},
      {stage0_12[104]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[34],stage1_13[55],stage1_12[127],stage1_11[158]}
   );
   gpc615_5 gpc458 (
      {stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage0_12[105]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[35],stage1_13[56],stage1_12[128],stage1_11[159]}
   );
   gpc615_5 gpc459 (
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254]},
      {stage0_12[106]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[36],stage1_13[57],stage1_12[129],stage1_11[160]}
   );
   gpc615_5 gpc460 (
      {stage0_11[255], stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259]},
      {stage0_12[107]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[37],stage1_13[58],stage1_12[130],stage1_11[161]}
   );
   gpc615_5 gpc461 (
      {stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263], stage0_11[264]},
      {stage0_12[108]},
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage1_15[24],stage1_14[38],stage1_13[59],stage1_12[131],stage1_11[162]}
   );
   gpc615_5 gpc462 (
      {stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage0_12[109]},
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage1_15[25],stage1_14[39],stage1_13[60],stage1_12[132],stage1_11[163]}
   );
   gpc615_5 gpc463 (
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274]},
      {stage0_12[110]},
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage1_15[26],stage1_14[40],stage1_13[61],stage1_12[133],stage1_11[164]}
   );
   gpc615_5 gpc464 (
      {stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage0_12[111]},
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage1_15[27],stage1_14[41],stage1_13[62],stage1_12[134],stage1_11[165]}
   );
   gpc615_5 gpc465 (
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[112]},
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage1_15[28],stage1_14[42],stage1_13[63],stage1_12[135],stage1_11[166]}
   );
   gpc615_5 gpc466 (
      {stage0_11[285], stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289]},
      {stage0_12[113]},
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage1_15[29],stage1_14[43],stage1_13[64],stage1_12[136],stage1_11[167]}
   );
   gpc615_5 gpc467 (
      {stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293], stage0_11[294]},
      {stage0_12[114]},
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage1_15[30],stage1_14[44],stage1_13[65],stage1_12[137],stage1_11[168]}
   );
   gpc615_5 gpc468 (
      {stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage0_12[115]},
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage1_15[31],stage1_14[45],stage1_13[66],stage1_12[138],stage1_11[169]}
   );
   gpc615_5 gpc469 (
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304]},
      {stage0_12[116]},
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage1_15[32],stage1_14[46],stage1_13[67],stage1_12[139],stage1_11[170]}
   );
   gpc615_5 gpc470 (
      {stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage0_12[117]},
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage1_15[33],stage1_14[47],stage1_13[68],stage1_12[140],stage1_11[171]}
   );
   gpc615_5 gpc471 (
      {stage0_11[310], stage0_11[311], stage0_11[312], stage0_11[313], stage0_11[314]},
      {stage0_12[118]},
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage1_15[34],stage1_14[48],stage1_13[69],stage1_12[141],stage1_11[172]}
   );
   gpc615_5 gpc472 (
      {stage0_11[315], stage0_11[316], stage0_11[317], stage0_11[318], stage0_11[319]},
      {stage0_12[119]},
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage1_15[35],stage1_14[49],stage1_13[70],stage1_12[142],stage1_11[173]}
   );
   gpc615_5 gpc473 (
      {stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323], stage0_11[324]},
      {stage0_12[120]},
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage1_15[36],stage1_14[50],stage1_13[71],stage1_12[143],stage1_11[174]}
   );
   gpc615_5 gpc474 (
      {stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage0_12[121]},
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage1_15[37],stage1_14[51],stage1_13[72],stage1_12[144],stage1_11[175]}
   );
   gpc615_5 gpc475 (
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334]},
      {stage0_12[122]},
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage1_15[38],stage1_14[52],stage1_13[73],stage1_12[145],stage1_11[176]}
   );
   gpc615_5 gpc476 (
      {stage0_11[335], stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339]},
      {stage0_12[123]},
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage1_15[39],stage1_14[53],stage1_13[74],stage1_12[146],stage1_11[177]}
   );
   gpc615_5 gpc477 (
      {stage0_11[340], stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344]},
      {stage0_12[124]},
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage1_15[40],stage1_14[54],stage1_13[75],stage1_12[147],stage1_11[178]}
   );
   gpc615_5 gpc478 (
      {stage0_11[345], stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349]},
      {stage0_12[125]},
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage1_15[41],stage1_14[55],stage1_13[76],stage1_12[148],stage1_11[179]}
   );
   gpc615_5 gpc479 (
      {stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354]},
      {stage0_12[126]},
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage1_15[42],stage1_14[56],stage1_13[77],stage1_12[149],stage1_11[180]}
   );
   gpc615_5 gpc480 (
      {stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage0_12[127]},
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage1_15[43],stage1_14[57],stage1_13[78],stage1_12[150],stage1_11[181]}
   );
   gpc615_5 gpc481 (
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364]},
      {stage0_12[128]},
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage1_15[44],stage1_14[58],stage1_13[79],stage1_12[151],stage1_11[182]}
   );
   gpc615_5 gpc482 (
      {stage0_11[365], stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369]},
      {stage0_12[129]},
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage1_15[45],stage1_14[59],stage1_13[80],stage1_12[152],stage1_11[183]}
   );
   gpc615_5 gpc483 (
      {stage0_11[370], stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374]},
      {stage0_12[130]},
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage1_15[46],stage1_14[60],stage1_13[81],stage1_12[153],stage1_11[184]}
   );
   gpc615_5 gpc484 (
      {stage0_11[375], stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379]},
      {stage0_12[131]},
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage1_15[47],stage1_14[61],stage1_13[82],stage1_12[154],stage1_11[185]}
   );
   gpc606_5 gpc485 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[48],stage1_14[62],stage1_13[83],stage1_12[155]}
   );
   gpc606_5 gpc486 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[49],stage1_14[63],stage1_13[84],stage1_12[156]}
   );
   gpc606_5 gpc487 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[50],stage1_14[64],stage1_13[85],stage1_12[157]}
   );
   gpc606_5 gpc488 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[51],stage1_14[65],stage1_13[86],stage1_12[158]}
   );
   gpc606_5 gpc489 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[52],stage1_14[66],stage1_13[87],stage1_12[159]}
   );
   gpc606_5 gpc490 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[53],stage1_14[67],stage1_13[88],stage1_12[160]}
   );
   gpc606_5 gpc491 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[54],stage1_14[68],stage1_13[89],stage1_12[161]}
   );
   gpc606_5 gpc492 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[55],stage1_14[69],stage1_13[90],stage1_12[162]}
   );
   gpc606_5 gpc493 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[56],stage1_14[70],stage1_13[91],stage1_12[163]}
   );
   gpc606_5 gpc494 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[57],stage1_14[71],stage1_13[92],stage1_12[164]}
   );
   gpc606_5 gpc495 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[58],stage1_14[72],stage1_13[93],stage1_12[165]}
   );
   gpc606_5 gpc496 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[59],stage1_14[73],stage1_13[94],stage1_12[166]}
   );
   gpc606_5 gpc497 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[60],stage1_14[74],stage1_13[95],stage1_12[167]}
   );
   gpc606_5 gpc498 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[61],stage1_14[75],stage1_13[96],stage1_12[168]}
   );
   gpc606_5 gpc499 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[62],stage1_14[76],stage1_13[97],stage1_12[169]}
   );
   gpc606_5 gpc500 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[63],stage1_14[77],stage1_13[98],stage1_12[170]}
   );
   gpc606_5 gpc501 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[64],stage1_14[78],stage1_13[99],stage1_12[171]}
   );
   gpc606_5 gpc502 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[65],stage1_14[79],stage1_13[100],stage1_12[172]}
   );
   gpc606_5 gpc503 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[66],stage1_14[80],stage1_13[101],stage1_12[173]}
   );
   gpc606_5 gpc504 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[67],stage1_14[81],stage1_13[102],stage1_12[174]}
   );
   gpc606_5 gpc505 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[68],stage1_14[82],stage1_13[103],stage1_12[175]}
   );
   gpc606_5 gpc506 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[69],stage1_14[83],stage1_13[104],stage1_12[176]}
   );
   gpc606_5 gpc507 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[70],stage1_14[84],stage1_13[105],stage1_12[177]}
   );
   gpc606_5 gpc508 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[71],stage1_14[85],stage1_13[106],stage1_12[178]}
   );
   gpc606_5 gpc509 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[72],stage1_14[86],stage1_13[107],stage1_12[179]}
   );
   gpc606_5 gpc510 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[73],stage1_14[87],stage1_13[108],stage1_12[180]}
   );
   gpc606_5 gpc511 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[74],stage1_14[88],stage1_13[109],stage1_12[181]}
   );
   gpc606_5 gpc512 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[75],stage1_14[89],stage1_13[110],stage1_12[182]}
   );
   gpc606_5 gpc513 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[76],stage1_14[90],stage1_13[111],stage1_12[183]}
   );
   gpc606_5 gpc514 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[77],stage1_14[91],stage1_13[112],stage1_12[184]}
   );
   gpc606_5 gpc515 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[78],stage1_14[92],stage1_13[113],stage1_12[185]}
   );
   gpc606_5 gpc516 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[79],stage1_14[93],stage1_13[114],stage1_12[186]}
   );
   gpc606_5 gpc517 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[80],stage1_14[94],stage1_13[115],stage1_12[187]}
   );
   gpc606_5 gpc518 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[81],stage1_14[95],stage1_13[116],stage1_12[188]}
   );
   gpc606_5 gpc519 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[82],stage1_14[96],stage1_13[117],stage1_12[189]}
   );
   gpc606_5 gpc520 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[83],stage1_14[97],stage1_13[118],stage1_12[190]}
   );
   gpc606_5 gpc521 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[84],stage1_14[98],stage1_13[119],stage1_12[191]}
   );
   gpc606_5 gpc522 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[85],stage1_14[99],stage1_13[120],stage1_12[192]}
   );
   gpc606_5 gpc523 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[86],stage1_14[100],stage1_13[121],stage1_12[193]}
   );
   gpc606_5 gpc524 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[87],stage1_14[101],stage1_13[122],stage1_12[194]}
   );
   gpc606_5 gpc525 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[88],stage1_14[102],stage1_13[123],stage1_12[195]}
   );
   gpc606_5 gpc526 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[89],stage1_14[103],stage1_13[124],stage1_12[196]}
   );
   gpc606_5 gpc527 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[90],stage1_14[104],stage1_13[125],stage1_12[197]}
   );
   gpc606_5 gpc528 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[91],stage1_14[105],stage1_13[126],stage1_12[198]}
   );
   gpc606_5 gpc529 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[92],stage1_14[106],stage1_13[127],stage1_12[199]}
   );
   gpc606_5 gpc530 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[93],stage1_14[107],stage1_13[128],stage1_12[200]}
   );
   gpc606_5 gpc531 (
      {stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[94],stage1_14[108],stage1_13[129],stage1_12[201]}
   );
   gpc606_5 gpc532 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[95],stage1_14[109],stage1_13[130],stage1_12[202]}
   );
   gpc606_5 gpc533 (
      {stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[96],stage1_14[110],stage1_13[131],stage1_12[203]}
   );
   gpc606_5 gpc534 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[97],stage1_14[111],stage1_13[132],stage1_12[204]}
   );
   gpc606_5 gpc535 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[98],stage1_14[112],stage1_13[133],stage1_12[205]}
   );
   gpc606_5 gpc536 (
      {stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[99],stage1_14[113],stage1_13[134],stage1_12[206]}
   );
   gpc606_5 gpc537 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[100],stage1_14[114],stage1_13[135],stage1_12[207]}
   );
   gpc606_5 gpc538 (
      {stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[101],stage1_14[115],stage1_13[136],stage1_12[208]}
   );
   gpc606_5 gpc539 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[102],stage1_14[116],stage1_13[137],stage1_12[209]}
   );
   gpc606_5 gpc540 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[103],stage1_14[117],stage1_13[138],stage1_12[210]}
   );
   gpc606_5 gpc541 (
      {stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[104],stage1_14[118],stage1_13[139],stage1_12[211]}
   );
   gpc606_5 gpc542 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[105],stage1_14[119],stage1_13[140],stage1_12[212]}
   );
   gpc606_5 gpc543 (
      {stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[106],stage1_14[120],stage1_13[141],stage1_12[213]}
   );
   gpc606_5 gpc544 (
      {stage0_12[486], stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[107],stage1_14[121],stage1_13[142],stage1_12[214]}
   );
   gpc606_5 gpc545 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496], stage0_12[497]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[108],stage1_14[122],stage1_13[143],stage1_12[215]}
   );
   gpc606_5 gpc546 (
      {stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501], stage0_12[502], stage0_12[503]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[109],stage1_14[123],stage1_13[144],stage1_12[216]}
   );
   gpc606_5 gpc547 (
      {stage0_12[504], stage0_12[505], stage0_12[506], stage0_12[507], stage0_12[508], stage0_12[509]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[110],stage1_14[124],stage1_13[145],stage1_12[217]}
   );
   gpc606_5 gpc548 (
      {stage0_12[510], stage0_12[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage1_16[63],stage1_15[111],stage1_14[125],stage1_13[146],stage1_12[218]}
   );
   gpc606_5 gpc549 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[64],stage1_15[112],stage1_14[126],stage1_13[147]}
   );
   gpc606_5 gpc550 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[65],stage1_15[113],stage1_14[127],stage1_13[148]}
   );
   gpc606_5 gpc551 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[66],stage1_15[114],stage1_14[128],stage1_13[149]}
   );
   gpc606_5 gpc552 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[67],stage1_15[115],stage1_14[129],stage1_13[150]}
   );
   gpc606_5 gpc553 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[68],stage1_15[116],stage1_14[130],stage1_13[151]}
   );
   gpc606_5 gpc554 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[69],stage1_15[117],stage1_14[131],stage1_13[152]}
   );
   gpc606_5 gpc555 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[70],stage1_15[118],stage1_14[132],stage1_13[153]}
   );
   gpc606_5 gpc556 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[71],stage1_15[119],stage1_14[133],stage1_13[154]}
   );
   gpc606_5 gpc557 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[72],stage1_15[120],stage1_14[134],stage1_13[155]}
   );
   gpc606_5 gpc558 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[73],stage1_15[121],stage1_14[135],stage1_13[156]}
   );
   gpc606_5 gpc559 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[74],stage1_15[122],stage1_14[136],stage1_13[157]}
   );
   gpc606_5 gpc560 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[75],stage1_15[123],stage1_14[137],stage1_13[158]}
   );
   gpc606_5 gpc561 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[76],stage1_15[124],stage1_14[138],stage1_13[159]}
   );
   gpc606_5 gpc562 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[77],stage1_15[125],stage1_14[139],stage1_13[160]}
   );
   gpc606_5 gpc563 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[78],stage1_15[126],stage1_14[140],stage1_13[161]}
   );
   gpc606_5 gpc564 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[79],stage1_15[127],stage1_14[141],stage1_13[162]}
   );
   gpc606_5 gpc565 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[80],stage1_15[128],stage1_14[142],stage1_13[163]}
   );
   gpc606_5 gpc566 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[81],stage1_15[129],stage1_14[143],stage1_13[164]}
   );
   gpc606_5 gpc567 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[82],stage1_15[130],stage1_14[144],stage1_13[165]}
   );
   gpc606_5 gpc568 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[83],stage1_15[131],stage1_14[145],stage1_13[166]}
   );
   gpc606_5 gpc569 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[84],stage1_15[132],stage1_14[146],stage1_13[167]}
   );
   gpc606_5 gpc570 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[85],stage1_15[133],stage1_14[147],stage1_13[168]}
   );
   gpc606_5 gpc571 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[86],stage1_15[134],stage1_14[148],stage1_13[169]}
   );
   gpc606_5 gpc572 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[87],stage1_15[135],stage1_14[149],stage1_13[170]}
   );
   gpc606_5 gpc573 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[88],stage1_15[136],stage1_14[150],stage1_13[171]}
   );
   gpc606_5 gpc574 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[89],stage1_15[137],stage1_14[151],stage1_13[172]}
   );
   gpc606_5 gpc575 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[90],stage1_15[138],stage1_14[152],stage1_13[173]}
   );
   gpc606_5 gpc576 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[91],stage1_15[139],stage1_14[153],stage1_13[174]}
   );
   gpc606_5 gpc577 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[92],stage1_15[140],stage1_14[154],stage1_13[175]}
   );
   gpc606_5 gpc578 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466], stage0_13[467]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[93],stage1_15[141],stage1_14[155],stage1_13[176]}
   );
   gpc606_5 gpc579 (
      {stage0_13[468], stage0_13[469], stage0_13[470], stage0_13[471], stage0_13[472], stage0_13[473]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[94],stage1_15[142],stage1_14[156],stage1_13[177]}
   );
   gpc606_5 gpc580 (
      {stage0_13[474], stage0_13[475], stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[95],stage1_15[143],stage1_14[157],stage1_13[178]}
   );
   gpc606_5 gpc581 (
      {stage0_13[480], stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[96],stage1_15[144],stage1_14[158],stage1_13[179]}
   );
   gpc606_5 gpc582 (
      {stage0_13[486], stage0_13[487], stage0_13[488], stage0_13[489], stage0_13[490], stage0_13[491]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[97],stage1_15[145],stage1_14[159],stage1_13[180]}
   );
   gpc606_5 gpc583 (
      {stage0_13[492], stage0_13[493], stage0_13[494], stage0_13[495], stage0_13[496], stage0_13[497]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[98],stage1_15[146],stage1_14[160],stage1_13[181]}
   );
   gpc606_5 gpc584 (
      {stage0_13[498], stage0_13[499], stage0_13[500], stage0_13[501], stage0_13[502], stage0_13[503]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[99],stage1_15[147],stage1_14[161],stage1_13[182]}
   );
   gpc606_5 gpc585 (
      {stage0_13[504], stage0_13[505], stage0_13[506], stage0_13[507], stage0_13[508], stage0_13[509]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[100],stage1_15[148],stage1_14[162],stage1_13[183]}
   );
   gpc606_5 gpc586 (
      {stage0_13[510], stage0_13[511], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[101],stage1_15[149],stage1_14[163],stage1_13[184]}
   );
   gpc615_5 gpc587 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388]},
      {stage0_15[228]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[38],stage1_16[102],stage1_15[150],stage1_14[164]}
   );
   gpc615_5 gpc588 (
      {stage0_14[389], stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393]},
      {stage0_15[229]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[39],stage1_16[103],stage1_15[151],stage1_14[165]}
   );
   gpc615_5 gpc589 (
      {stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397], stage0_14[398]},
      {stage0_15[230]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[40],stage1_16[104],stage1_15[152],stage1_14[166]}
   );
   gpc615_5 gpc590 (
      {stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage0_15[231]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[41],stage1_16[105],stage1_15[153],stage1_14[167]}
   );
   gpc615_5 gpc591 (
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408]},
      {stage0_15[232]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[42],stage1_16[106],stage1_15[154],stage1_14[168]}
   );
   gpc615_5 gpc592 (
      {stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_15[233]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[43],stage1_16[107],stage1_15[155],stage1_14[169]}
   );
   gpc615_5 gpc593 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_15[234]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[44],stage1_16[108],stage1_15[156],stage1_14[170]}
   );
   gpc615_5 gpc594 (
      {stage0_14[419], stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423]},
      {stage0_15[235]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[45],stage1_16[109],stage1_15[157],stage1_14[171]}
   );
   gpc615_5 gpc595 (
      {stage0_14[424], stage0_14[425], stage0_14[426], stage0_14[427], stage0_14[428]},
      {stage0_15[236]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[46],stage1_16[110],stage1_15[158],stage1_14[172]}
   );
   gpc615_5 gpc596 (
      {stage0_15[237], stage0_15[238], stage0_15[239], stage0_15[240], stage0_15[241]},
      {stage0_16[54]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[9],stage1_17[47],stage1_16[111],stage1_15[159]}
   );
   gpc615_5 gpc597 (
      {stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245], stage0_15[246]},
      {stage0_16[55]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[10],stage1_17[48],stage1_16[112],stage1_15[160]}
   );
   gpc615_5 gpc598 (
      {stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage0_16[56]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[11],stage1_17[49],stage1_16[113],stage1_15[161]}
   );
   gpc615_5 gpc599 (
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256]},
      {stage0_16[57]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[12],stage1_17[50],stage1_16[114],stage1_15[162]}
   );
   gpc615_5 gpc600 (
      {stage0_15[257], stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261]},
      {stage0_16[58]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[13],stage1_17[51],stage1_16[115],stage1_15[163]}
   );
   gpc615_5 gpc601 (
      {stage0_15[262], stage0_15[263], stage0_15[264], stage0_15[265], stage0_15[266]},
      {stage0_16[59]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[14],stage1_17[52],stage1_16[116],stage1_15[164]}
   );
   gpc615_5 gpc602 (
      {stage0_15[267], stage0_15[268], stage0_15[269], stage0_15[270], stage0_15[271]},
      {stage0_16[60]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[15],stage1_17[53],stage1_16[117],stage1_15[165]}
   );
   gpc615_5 gpc603 (
      {stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275], stage0_15[276]},
      {stage0_16[61]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[16],stage1_17[54],stage1_16[118],stage1_15[166]}
   );
   gpc615_5 gpc604 (
      {stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage0_16[62]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[17],stage1_17[55],stage1_16[119],stage1_15[167]}
   );
   gpc615_5 gpc605 (
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286]},
      {stage0_16[63]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[18],stage1_17[56],stage1_16[120],stage1_15[168]}
   );
   gpc615_5 gpc606 (
      {stage0_15[287], stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291]},
      {stage0_16[64]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[19],stage1_17[57],stage1_16[121],stage1_15[169]}
   );
   gpc615_5 gpc607 (
      {stage0_15[292], stage0_15[293], stage0_15[294], stage0_15[295], stage0_15[296]},
      {stage0_16[65]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[20],stage1_17[58],stage1_16[122],stage1_15[170]}
   );
   gpc615_5 gpc608 (
      {stage0_15[297], stage0_15[298], stage0_15[299], stage0_15[300], stage0_15[301]},
      {stage0_16[66]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[21],stage1_17[59],stage1_16[123],stage1_15[171]}
   );
   gpc615_5 gpc609 (
      {stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305], stage0_15[306]},
      {stage0_16[67]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[22],stage1_17[60],stage1_16[124],stage1_15[172]}
   );
   gpc615_5 gpc610 (
      {stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage0_16[68]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[23],stage1_17[61],stage1_16[125],stage1_15[173]}
   );
   gpc615_5 gpc611 (
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316]},
      {stage0_16[69]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[24],stage1_17[62],stage1_16[126],stage1_15[174]}
   );
   gpc615_5 gpc612 (
      {stage0_15[317], stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321]},
      {stage0_16[70]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[25],stage1_17[63],stage1_16[127],stage1_15[175]}
   );
   gpc615_5 gpc613 (
      {stage0_15[322], stage0_15[323], stage0_15[324], stage0_15[325], stage0_15[326]},
      {stage0_16[71]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[26],stage1_17[64],stage1_16[128],stage1_15[176]}
   );
   gpc615_5 gpc614 (
      {stage0_15[327], stage0_15[328], stage0_15[329], stage0_15[330], stage0_15[331]},
      {stage0_16[72]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[27],stage1_17[65],stage1_16[129],stage1_15[177]}
   );
   gpc615_5 gpc615 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336]},
      {stage0_16[73]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[28],stage1_17[66],stage1_16[130],stage1_15[178]}
   );
   gpc615_5 gpc616 (
      {stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage0_16[74]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[29],stage1_17[67],stage1_16[131],stage1_15[179]}
   );
   gpc615_5 gpc617 (
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346]},
      {stage0_16[75]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[30],stage1_17[68],stage1_16[132],stage1_15[180]}
   );
   gpc615_5 gpc618 (
      {stage0_15[347], stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351]},
      {stage0_16[76]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[31],stage1_17[69],stage1_16[133],stage1_15[181]}
   );
   gpc615_5 gpc619 (
      {stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355], stage0_15[356]},
      {stage0_16[77]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[32],stage1_17[70],stage1_16[134],stage1_15[182]}
   );
   gpc615_5 gpc620 (
      {stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360], stage0_15[361]},
      {stage0_16[78]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[33],stage1_17[71],stage1_16[135],stage1_15[183]}
   );
   gpc615_5 gpc621 (
      {stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365], stage0_15[366]},
      {stage0_16[79]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[34],stage1_17[72],stage1_16[136],stage1_15[184]}
   );
   gpc615_5 gpc622 (
      {stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage0_16[80]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[35],stage1_17[73],stage1_16[137],stage1_15[185]}
   );
   gpc615_5 gpc623 (
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376]},
      {stage0_16[81]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[36],stage1_17[74],stage1_16[138],stage1_15[186]}
   );
   gpc615_5 gpc624 (
      {stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381]},
      {stage0_16[82]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[37],stage1_17[75],stage1_16[139],stage1_15[187]}
   );
   gpc615_5 gpc625 (
      {stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385], stage0_15[386]},
      {stage0_16[83]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[38],stage1_17[76],stage1_16[140],stage1_15[188]}
   );
   gpc615_5 gpc626 (
      {stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390], stage0_15[391]},
      {stage0_16[84]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[39],stage1_17[77],stage1_16[141],stage1_15[189]}
   );
   gpc615_5 gpc627 (
      {stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395], stage0_15[396]},
      {stage0_16[85]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[40],stage1_17[78],stage1_16[142],stage1_15[190]}
   );
   gpc615_5 gpc628 (
      {stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage0_16[86]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[41],stage1_17[79],stage1_16[143],stage1_15[191]}
   );
   gpc615_5 gpc629 (
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406]},
      {stage0_16[87]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[42],stage1_17[80],stage1_16[144],stage1_15[192]}
   );
   gpc615_5 gpc630 (
      {stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411]},
      {stage0_16[88]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[43],stage1_17[81],stage1_16[145],stage1_15[193]}
   );
   gpc615_5 gpc631 (
      {stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415], stage0_15[416]},
      {stage0_16[89]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[44],stage1_17[82],stage1_16[146],stage1_15[194]}
   );
   gpc615_5 gpc632 (
      {stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420], stage0_15[421]},
      {stage0_16[90]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[45],stage1_17[83],stage1_16[147],stage1_15[195]}
   );
   gpc615_5 gpc633 (
      {stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425], stage0_15[426]},
      {stage0_16[91]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[46],stage1_17[84],stage1_16[148],stage1_15[196]}
   );
   gpc615_5 gpc634 (
      {stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage0_16[92]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[47],stage1_17[85],stage1_16[149],stage1_15[197]}
   );
   gpc615_5 gpc635 (
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436]},
      {stage0_16[93]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[48],stage1_17[86],stage1_16[150],stage1_15[198]}
   );
   gpc615_5 gpc636 (
      {stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441]},
      {stage0_16[94]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[49],stage1_17[87],stage1_16[151],stage1_15[199]}
   );
   gpc615_5 gpc637 (
      {stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445], stage0_15[446]},
      {stage0_16[95]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[50],stage1_17[88],stage1_16[152],stage1_15[200]}
   );
   gpc615_5 gpc638 (
      {stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450], stage0_15[451]},
      {stage0_16[96]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[51],stage1_17[89],stage1_16[153],stage1_15[201]}
   );
   gpc615_5 gpc639 (
      {stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455], stage0_15[456]},
      {stage0_16[97]},
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage1_19[43],stage1_18[52],stage1_17[90],stage1_16[154],stage1_15[202]}
   );
   gpc606_5 gpc640 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[44],stage1_18[53],stage1_17[91],stage1_16[155]}
   );
   gpc606_5 gpc641 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[45],stage1_18[54],stage1_17[92],stage1_16[156]}
   );
   gpc606_5 gpc642 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[46],stage1_18[55],stage1_17[93],stage1_16[157]}
   );
   gpc606_5 gpc643 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[47],stage1_18[56],stage1_17[94],stage1_16[158]}
   );
   gpc606_5 gpc644 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[48],stage1_18[57],stage1_17[95],stage1_16[159]}
   );
   gpc606_5 gpc645 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[49],stage1_18[58],stage1_17[96],stage1_16[160]}
   );
   gpc606_5 gpc646 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[50],stage1_18[59],stage1_17[97],stage1_16[161]}
   );
   gpc606_5 gpc647 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[51],stage1_18[60],stage1_17[98],stage1_16[162]}
   );
   gpc606_5 gpc648 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[52],stage1_18[61],stage1_17[99],stage1_16[163]}
   );
   gpc606_5 gpc649 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[53],stage1_18[62],stage1_17[100],stage1_16[164]}
   );
   gpc606_5 gpc650 (
      {stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[54],stage1_18[63],stage1_17[101],stage1_16[165]}
   );
   gpc606_5 gpc651 (
      {stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[55],stage1_18[64],stage1_17[102],stage1_16[166]}
   );
   gpc606_5 gpc652 (
      {stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[56],stage1_18[65],stage1_17[103],stage1_16[167]}
   );
   gpc606_5 gpc653 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[57],stage1_18[66],stage1_17[104],stage1_16[168]}
   );
   gpc606_5 gpc654 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[58],stage1_18[67],stage1_17[105],stage1_16[169]}
   );
   gpc606_5 gpc655 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[59],stage1_18[68],stage1_17[106],stage1_16[170]}
   );
   gpc606_5 gpc656 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[60],stage1_18[69],stage1_17[107],stage1_16[171]}
   );
   gpc606_5 gpc657 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[61],stage1_18[70],stage1_17[108],stage1_16[172]}
   );
   gpc606_5 gpc658 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[62],stage1_18[71],stage1_17[109],stage1_16[173]}
   );
   gpc606_5 gpc659 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[63],stage1_18[72],stage1_17[110],stage1_16[174]}
   );
   gpc606_5 gpc660 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[64],stage1_18[73],stage1_17[111],stage1_16[175]}
   );
   gpc606_5 gpc661 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[65],stage1_18[74],stage1_17[112],stage1_16[176]}
   );
   gpc606_5 gpc662 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[66],stage1_18[75],stage1_17[113],stage1_16[177]}
   );
   gpc606_5 gpc663 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[67],stage1_18[76],stage1_17[114],stage1_16[178]}
   );
   gpc606_5 gpc664 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[68],stage1_18[77],stage1_17[115],stage1_16[179]}
   );
   gpc606_5 gpc665 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[69],stage1_18[78],stage1_17[116],stage1_16[180]}
   );
   gpc606_5 gpc666 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[70],stage1_18[79],stage1_17[117],stage1_16[181]}
   );
   gpc606_5 gpc667 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[71],stage1_18[80],stage1_17[118],stage1_16[182]}
   );
   gpc606_5 gpc668 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[72],stage1_18[81],stage1_17[119],stage1_16[183]}
   );
   gpc606_5 gpc669 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[73],stage1_18[82],stage1_17[120],stage1_16[184]}
   );
   gpc606_5 gpc670 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[74],stage1_18[83],stage1_17[121],stage1_16[185]}
   );
   gpc606_5 gpc671 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[75],stage1_18[84],stage1_17[122],stage1_16[186]}
   );
   gpc606_5 gpc672 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[76],stage1_18[85],stage1_17[123],stage1_16[187]}
   );
   gpc606_5 gpc673 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[77],stage1_18[86],stage1_17[124],stage1_16[188]}
   );
   gpc606_5 gpc674 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[78],stage1_18[87],stage1_17[125],stage1_16[189]}
   );
   gpc606_5 gpc675 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[79],stage1_18[88],stage1_17[126],stage1_16[190]}
   );
   gpc606_5 gpc676 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[80],stage1_18[89],stage1_17[127],stage1_16[191]}
   );
   gpc606_5 gpc677 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[81],stage1_18[90],stage1_17[128],stage1_16[192]}
   );
   gpc606_5 gpc678 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[82],stage1_18[91],stage1_17[129],stage1_16[193]}
   );
   gpc606_5 gpc679 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[83],stage1_18[92],stage1_17[130],stage1_16[194]}
   );
   gpc606_5 gpc680 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[84],stage1_18[93],stage1_17[131],stage1_16[195]}
   );
   gpc606_5 gpc681 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[85],stage1_18[94],stage1_17[132],stage1_16[196]}
   );
   gpc606_5 gpc682 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[86],stage1_18[95],stage1_17[133],stage1_16[197]}
   );
   gpc606_5 gpc683 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[87],stage1_18[96],stage1_17[134],stage1_16[198]}
   );
   gpc606_5 gpc684 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[88],stage1_18[97],stage1_17[135],stage1_16[199]}
   );
   gpc606_5 gpc685 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[89],stage1_18[98],stage1_17[136],stage1_16[200]}
   );
   gpc606_5 gpc686 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[90],stage1_18[99],stage1_17[137],stage1_16[201]}
   );
   gpc606_5 gpc687 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[91],stage1_18[100],stage1_17[138],stage1_16[202]}
   );
   gpc606_5 gpc688 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[92],stage1_18[101],stage1_17[139],stage1_16[203]}
   );
   gpc606_5 gpc689 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[93],stage1_18[102],stage1_17[140],stage1_16[204]}
   );
   gpc606_5 gpc690 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[94],stage1_18[103],stage1_17[141],stage1_16[205]}
   );
   gpc606_5 gpc691 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[95],stage1_18[104],stage1_17[142],stage1_16[206]}
   );
   gpc606_5 gpc692 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[96],stage1_18[105],stage1_17[143],stage1_16[207]}
   );
   gpc606_5 gpc693 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[97],stage1_18[106],stage1_17[144],stage1_16[208]}
   );
   gpc606_5 gpc694 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[98],stage1_18[107],stage1_17[145],stage1_16[209]}
   );
   gpc606_5 gpc695 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[99],stage1_18[108],stage1_17[146],stage1_16[210]}
   );
   gpc606_5 gpc696 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[100],stage1_18[109],stage1_17[147],stage1_16[211]}
   );
   gpc606_5 gpc697 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[101],stage1_18[110],stage1_17[148],stage1_16[212]}
   );
   gpc606_5 gpc698 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[102],stage1_18[111],stage1_17[149],stage1_16[213]}
   );
   gpc606_5 gpc699 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[103],stage1_18[112],stage1_17[150],stage1_16[214]}
   );
   gpc606_5 gpc700 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[104],stage1_18[113],stage1_17[151],stage1_16[215]}
   );
   gpc606_5 gpc701 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[105],stage1_18[114],stage1_17[152],stage1_16[216]}
   );
   gpc606_5 gpc702 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[106],stage1_18[115],stage1_17[153],stage1_16[217]}
   );
   gpc606_5 gpc703 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[107],stage1_18[116],stage1_17[154],stage1_16[218]}
   );
   gpc606_5 gpc704 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[108],stage1_18[117],stage1_17[155],stage1_16[219]}
   );
   gpc606_5 gpc705 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[109],stage1_18[118],stage1_17[156],stage1_16[220]}
   );
   gpc606_5 gpc706 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[110],stage1_18[119],stage1_17[157],stage1_16[221]}
   );
   gpc606_5 gpc707 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[111],stage1_18[120],stage1_17[158],stage1_16[222]}
   );
   gpc606_5 gpc708 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[112],stage1_18[121],stage1_17[159],stage1_16[223]}
   );
   gpc606_5 gpc709 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[69],stage1_19[113],stage1_18[122],stage1_17[160]}
   );
   gpc606_5 gpc710 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[70],stage1_19[114],stage1_18[123],stage1_17[161]}
   );
   gpc606_5 gpc711 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[71],stage1_19[115],stage1_18[124],stage1_17[162]}
   );
   gpc606_5 gpc712 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[72],stage1_19[116],stage1_18[125],stage1_17[163]}
   );
   gpc606_5 gpc713 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[73],stage1_19[117],stage1_18[126],stage1_17[164]}
   );
   gpc606_5 gpc714 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[74],stage1_19[118],stage1_18[127],stage1_17[165]}
   );
   gpc606_5 gpc715 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[75],stage1_19[119],stage1_18[128],stage1_17[166]}
   );
   gpc606_5 gpc716 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[76],stage1_19[120],stage1_18[129],stage1_17[167]}
   );
   gpc606_5 gpc717 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[77],stage1_19[121],stage1_18[130],stage1_17[168]}
   );
   gpc606_5 gpc718 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[78],stage1_19[122],stage1_18[131],stage1_17[169]}
   );
   gpc606_5 gpc719 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[79],stage1_19[123],stage1_18[132],stage1_17[170]}
   );
   gpc606_5 gpc720 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[80],stage1_19[124],stage1_18[133],stage1_17[171]}
   );
   gpc606_5 gpc721 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[81],stage1_19[125],stage1_18[134],stage1_17[172]}
   );
   gpc606_5 gpc722 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[82],stage1_19[126],stage1_18[135],stage1_17[173]}
   );
   gpc606_5 gpc723 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[83],stage1_19[127],stage1_18[136],stage1_17[174]}
   );
   gpc606_5 gpc724 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[84],stage1_19[128],stage1_18[137],stage1_17[175]}
   );
   gpc606_5 gpc725 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[85],stage1_19[129],stage1_18[138],stage1_17[176]}
   );
   gpc606_5 gpc726 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[86],stage1_19[130],stage1_18[139],stage1_17[177]}
   );
   gpc606_5 gpc727 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[87],stage1_19[131],stage1_18[140],stage1_17[178]}
   );
   gpc606_5 gpc728 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[88],stage1_19[132],stage1_18[141],stage1_17[179]}
   );
   gpc606_5 gpc729 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[89],stage1_19[133],stage1_18[142],stage1_17[180]}
   );
   gpc606_5 gpc730 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[90],stage1_19[134],stage1_18[143],stage1_17[181]}
   );
   gpc606_5 gpc731 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[91],stage1_19[135],stage1_18[144],stage1_17[182]}
   );
   gpc606_5 gpc732 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[92],stage1_19[136],stage1_18[145],stage1_17[183]}
   );
   gpc606_5 gpc733 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[93],stage1_19[137],stage1_18[146],stage1_17[184]}
   );
   gpc606_5 gpc734 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[94],stage1_19[138],stage1_18[147],stage1_17[185]}
   );
   gpc606_5 gpc735 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[95],stage1_19[139],stage1_18[148],stage1_17[186]}
   );
   gpc606_5 gpc736 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[96],stage1_19[140],stage1_18[149],stage1_17[187]}
   );
   gpc606_5 gpc737 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[97],stage1_19[141],stage1_18[150],stage1_17[188]}
   );
   gpc606_5 gpc738 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[98],stage1_19[142],stage1_18[151],stage1_17[189]}
   );
   gpc606_5 gpc739 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[99],stage1_19[143],stage1_18[152],stage1_17[190]}
   );
   gpc606_5 gpc740 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[100],stage1_19[144],stage1_18[153],stage1_17[191]}
   );
   gpc606_5 gpc741 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[101],stage1_19[145],stage1_18[154],stage1_17[192]}
   );
   gpc606_5 gpc742 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[102],stage1_19[146],stage1_18[155],stage1_17[193]}
   );
   gpc606_5 gpc743 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[103],stage1_19[147],stage1_18[156],stage1_17[194]}
   );
   gpc606_5 gpc744 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[104],stage1_19[148],stage1_18[157],stage1_17[195]}
   );
   gpc606_5 gpc745 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[105],stage1_19[149],stage1_18[158],stage1_17[196]}
   );
   gpc606_5 gpc746 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[106],stage1_19[150],stage1_18[159],stage1_17[197]}
   );
   gpc615_5 gpc747 (
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418]},
      {stage0_19[228]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[107],stage1_19[151],stage1_18[160]}
   );
   gpc615_5 gpc748 (
      {stage0_18[419], stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423]},
      {stage0_19[229]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[108],stage1_19[152],stage1_18[161]}
   );
   gpc615_5 gpc749 (
      {stage0_18[424], stage0_18[425], stage0_18[426], stage0_18[427], stage0_18[428]},
      {stage0_19[230]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[109],stage1_19[153],stage1_18[162]}
   );
   gpc615_5 gpc750 (
      {stage0_18[429], stage0_18[430], stage0_18[431], stage0_18[432], stage0_18[433]},
      {stage0_19[231]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[110],stage1_19[154],stage1_18[163]}
   );
   gpc615_5 gpc751 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[24]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[42],stage1_20[111],stage1_19[155]}
   );
   gpc615_5 gpc752 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[25]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[43],stage1_20[112],stage1_19[156]}
   );
   gpc615_5 gpc753 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[26]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[44],stage1_20[113],stage1_19[157]}
   );
   gpc615_5 gpc754 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[27]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[7],stage1_21[45],stage1_20[114],stage1_19[158]}
   );
   gpc615_5 gpc755 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[28]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[8],stage1_21[46],stage1_20[115],stage1_19[159]}
   );
   gpc615_5 gpc756 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[29]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[9],stage1_21[47],stage1_20[116],stage1_19[160]}
   );
   gpc615_5 gpc757 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[30]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[10],stage1_21[48],stage1_20[117],stage1_19[161]}
   );
   gpc615_5 gpc758 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[31]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[11],stage1_21[49],stage1_20[118],stage1_19[162]}
   );
   gpc615_5 gpc759 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[32]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[12],stage1_21[50],stage1_20[119],stage1_19[163]}
   );
   gpc615_5 gpc760 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[33]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[13],stage1_21[51],stage1_20[120],stage1_19[164]}
   );
   gpc615_5 gpc761 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[34]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[14],stage1_21[52],stage1_20[121],stage1_19[165]}
   );
   gpc615_5 gpc762 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[35]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[15],stage1_21[53],stage1_20[122],stage1_19[166]}
   );
   gpc615_5 gpc763 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[36]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[16],stage1_21[54],stage1_20[123],stage1_19[167]}
   );
   gpc615_5 gpc764 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[37]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[17],stage1_21[55],stage1_20[124],stage1_19[168]}
   );
   gpc615_5 gpc765 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[38]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[18],stage1_21[56],stage1_20[125],stage1_19[169]}
   );
   gpc615_5 gpc766 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[39]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[19],stage1_21[57],stage1_20[126],stage1_19[170]}
   );
   gpc615_5 gpc767 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[40]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[20],stage1_21[58],stage1_20[127],stage1_19[171]}
   );
   gpc615_5 gpc768 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[41]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[21],stage1_21[59],stage1_20[128],stage1_19[172]}
   );
   gpc615_5 gpc769 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[42]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[22],stage1_21[60],stage1_20[129],stage1_19[173]}
   );
   gpc615_5 gpc770 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[43]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[23],stage1_21[61],stage1_20[130],stage1_19[174]}
   );
   gpc615_5 gpc771 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[44]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[24],stage1_21[62],stage1_20[131],stage1_19[175]}
   );
   gpc615_5 gpc772 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[45]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[25],stage1_21[63],stage1_20[132],stage1_19[176]}
   );
   gpc615_5 gpc773 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[46]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[26],stage1_21[64],stage1_20[133],stage1_19[177]}
   );
   gpc615_5 gpc774 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[47]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[27],stage1_21[65],stage1_20[134],stage1_19[178]}
   );
   gpc615_5 gpc775 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[48]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[28],stage1_21[66],stage1_20[135],stage1_19[179]}
   );
   gpc615_5 gpc776 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[49]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[29],stage1_21[67],stage1_20[136],stage1_19[180]}
   );
   gpc615_5 gpc777 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[50]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[30],stage1_21[68],stage1_20[137],stage1_19[181]}
   );
   gpc615_5 gpc778 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[51]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[31],stage1_21[69],stage1_20[138],stage1_19[182]}
   );
   gpc615_5 gpc779 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[52]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[32],stage1_21[70],stage1_20[139],stage1_19[183]}
   );
   gpc615_5 gpc780 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[53]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[33],stage1_21[71],stage1_20[140],stage1_19[184]}
   );
   gpc615_5 gpc781 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[54]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[34],stage1_21[72],stage1_20[141],stage1_19[185]}
   );
   gpc615_5 gpc782 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[55]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[35],stage1_21[73],stage1_20[142],stage1_19[186]}
   );
   gpc615_5 gpc783 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[56]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[36],stage1_21[74],stage1_20[143],stage1_19[187]}
   );
   gpc615_5 gpc784 (
      {stage0_19[397], stage0_19[398], stage0_19[399], stage0_19[400], stage0_19[401]},
      {stage0_20[57]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[37],stage1_21[75],stage1_20[144],stage1_19[188]}
   );
   gpc615_5 gpc785 (
      {stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405], stage0_19[406]},
      {stage0_20[58]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[38],stage1_21[76],stage1_20[145],stage1_19[189]}
   );
   gpc615_5 gpc786 (
      {stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410], stage0_19[411]},
      {stage0_20[59]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[39],stage1_21[77],stage1_20[146],stage1_19[190]}
   );
   gpc615_5 gpc787 (
      {stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415], stage0_19[416]},
      {stage0_20[60]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[40],stage1_21[78],stage1_20[147],stage1_19[191]}
   );
   gpc615_5 gpc788 (
      {stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420], stage0_19[421]},
      {stage0_20[61]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[41],stage1_21[79],stage1_20[148],stage1_19[192]}
   );
   gpc615_5 gpc789 (
      {stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425], stage0_19[426]},
      {stage0_20[62]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[42],stage1_21[80],stage1_20[149],stage1_19[193]}
   );
   gpc615_5 gpc790 (
      {stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430], stage0_19[431]},
      {stage0_20[63]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[43],stage1_21[81],stage1_20[150],stage1_19[194]}
   );
   gpc615_5 gpc791 (
      {stage0_19[432], stage0_19[433], stage0_19[434], stage0_19[435], stage0_19[436]},
      {stage0_20[64]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[44],stage1_21[82],stage1_20[151],stage1_19[195]}
   );
   gpc615_5 gpc792 (
      {stage0_19[437], stage0_19[438], stage0_19[439], stage0_19[440], stage0_19[441]},
      {stage0_20[65]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage1_23[41],stage1_22[45],stage1_21[83],stage1_20[152],stage1_19[196]}
   );
   gpc615_5 gpc793 (
      {stage0_19[442], stage0_19[443], stage0_19[444], stage0_19[445], stage0_19[446]},
      {stage0_20[66]},
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage1_23[42],stage1_22[46],stage1_21[84],stage1_20[153],stage1_19[197]}
   );
   gpc615_5 gpc794 (
      {stage0_19[447], stage0_19[448], stage0_19[449], stage0_19[450], stage0_19[451]},
      {stage0_20[67]},
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage1_23[43],stage1_22[47],stage1_21[85],stage1_20[154],stage1_19[198]}
   );
   gpc615_5 gpc795 (
      {stage0_19[452], stage0_19[453], stage0_19[454], stage0_19[455], stage0_19[456]},
      {stage0_20[68]},
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage1_23[44],stage1_22[48],stage1_21[86],stage1_20[155],stage1_19[199]}
   );
   gpc615_5 gpc796 (
      {stage0_19[457], stage0_19[458], stage0_19[459], stage0_19[460], stage0_19[461]},
      {stage0_20[69]},
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage1_23[45],stage1_22[49],stage1_21[87],stage1_20[156],stage1_19[200]}
   );
   gpc615_5 gpc797 (
      {stage0_19[462], stage0_19[463], stage0_19[464], stage0_19[465], stage0_19[466]},
      {stage0_20[70]},
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage1_23[46],stage1_22[50],stage1_21[88],stage1_20[157],stage1_19[201]}
   );
   gpc615_5 gpc798 (
      {stage0_19[467], stage0_19[468], stage0_19[469], stage0_19[470], stage0_19[471]},
      {stage0_20[71]},
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage1_23[47],stage1_22[51],stage1_21[89],stage1_20[158],stage1_19[202]}
   );
   gpc615_5 gpc799 (
      {stage0_19[472], stage0_19[473], stage0_19[474], stage0_19[475], stage0_19[476]},
      {stage0_20[72]},
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage1_23[48],stage1_22[52],stage1_21[90],stage1_20[159],stage1_19[203]}
   );
   gpc615_5 gpc800 (
      {stage0_19[477], stage0_19[478], stage0_19[479], stage0_19[480], stage0_19[481]},
      {stage0_20[73]},
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage1_23[49],stage1_22[53],stage1_21[91],stage1_20[160],stage1_19[204]}
   );
   gpc615_5 gpc801 (
      {stage0_19[482], stage0_19[483], stage0_19[484], stage0_19[485], stage0_19[486]},
      {stage0_20[74]},
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage1_23[50],stage1_22[54],stage1_21[92],stage1_20[161],stage1_19[205]}
   );
   gpc615_5 gpc802 (
      {stage0_19[487], stage0_19[488], stage0_19[489], stage0_19[490], stage0_19[491]},
      {stage0_20[75]},
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage1_23[51],stage1_22[55],stage1_21[93],stage1_20[162],stage1_19[206]}
   );
   gpc615_5 gpc803 (
      {stage0_19[492], stage0_19[493], stage0_19[494], stage0_19[495], stage0_19[496]},
      {stage0_20[76]},
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage1_23[52],stage1_22[56],stage1_21[94],stage1_20[163],stage1_19[207]}
   );
   gpc615_5 gpc804 (
      {stage0_19[497], stage0_19[498], stage0_19[499], stage0_19[500], stage0_19[501]},
      {stage0_20[77]},
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage1_23[53],stage1_22[57],stage1_21[95],stage1_20[164],stage1_19[208]}
   );
   gpc606_5 gpc805 (
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[54],stage1_22[58],stage1_21[96],stage1_20[165]}
   );
   gpc606_5 gpc806 (
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[55],stage1_22[59],stage1_21[97],stage1_20[166]}
   );
   gpc606_5 gpc807 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[56],stage1_22[60],stage1_21[98],stage1_20[167]}
   );
   gpc606_5 gpc808 (
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[57],stage1_22[61],stage1_21[99],stage1_20[168]}
   );
   gpc606_5 gpc809 (
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[58],stage1_22[62],stage1_21[100],stage1_20[169]}
   );
   gpc606_5 gpc810 (
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[59],stage1_22[63],stage1_21[101],stage1_20[170]}
   );
   gpc606_5 gpc811 (
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[60],stage1_22[64],stage1_21[102],stage1_20[171]}
   );
   gpc606_5 gpc812 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[61],stage1_22[65],stage1_21[103],stage1_20[172]}
   );
   gpc606_5 gpc813 (
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[62],stage1_22[66],stage1_21[104],stage1_20[173]}
   );
   gpc606_5 gpc814 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[63],stage1_22[67],stage1_21[105],stage1_20[174]}
   );
   gpc606_5 gpc815 (
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[64],stage1_22[68],stage1_21[106],stage1_20[175]}
   );
   gpc606_5 gpc816 (
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[65],stage1_22[69],stage1_21[107],stage1_20[176]}
   );
   gpc606_5 gpc817 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[66],stage1_22[70],stage1_21[108],stage1_20[177]}
   );
   gpc606_5 gpc818 (
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[67],stage1_22[71],stage1_21[109],stage1_20[178]}
   );
   gpc606_5 gpc819 (
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[68],stage1_22[72],stage1_21[110],stage1_20[179]}
   );
   gpc606_5 gpc820 (
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[69],stage1_22[73],stage1_21[111],stage1_20[180]}
   );
   gpc606_5 gpc821 (
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[70],stage1_22[74],stage1_21[112],stage1_20[181]}
   );
   gpc606_5 gpc822 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[71],stage1_22[75],stage1_21[113],stage1_20[182]}
   );
   gpc606_5 gpc823 (
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[72],stage1_22[76],stage1_21[114],stage1_20[183]}
   );
   gpc606_5 gpc824 (
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[73],stage1_22[77],stage1_21[115],stage1_20[184]}
   );
   gpc606_5 gpc825 (
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[74],stage1_22[78],stage1_21[116],stage1_20[185]}
   );
   gpc606_5 gpc826 (
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[75],stage1_22[79],stage1_21[117],stage1_20[186]}
   );
   gpc606_5 gpc827 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[76],stage1_22[80],stage1_21[118],stage1_20[187]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[77],stage1_22[81],stage1_21[119],stage1_20[188]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[78],stage1_22[82],stage1_21[120],stage1_20[189]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[79],stage1_22[83],stage1_21[121],stage1_20[190]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[80],stage1_22[84],stage1_21[122],stage1_20[191]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[81],stage1_22[85],stage1_21[123],stage1_20[192]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[82],stage1_22[86],stage1_21[124],stage1_20[193]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[83],stage1_22[87],stage1_21[125],stage1_20[194]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[84],stage1_22[88],stage1_21[126],stage1_20[195]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[85],stage1_22[89],stage1_21[127],stage1_20[196]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[86],stage1_22[90],stage1_21[128],stage1_20[197]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[87],stage1_22[91],stage1_21[129],stage1_20[198]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[88],stage1_22[92],stage1_21[130],stage1_20[199]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[89],stage1_22[93],stage1_21[131],stage1_20[200]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[90],stage1_22[94],stage1_21[132],stage1_20[201]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[91],stage1_22[95],stage1_21[133],stage1_20[202]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[92],stage1_22[96],stage1_21[134],stage1_20[203]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[93],stage1_22[97],stage1_21[135],stage1_20[204]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[94],stage1_22[98],stage1_21[136],stage1_20[205]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[95],stage1_22[99],stage1_21[137],stage1_20[206]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[96],stage1_22[100],stage1_21[138],stage1_20[207]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[97],stage1_22[101],stage1_21[139],stage1_20[208]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[98],stage1_22[102],stage1_21[140],stage1_20[209]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[99],stage1_22[103],stage1_21[141],stage1_20[210]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[100],stage1_22[104],stage1_21[142],stage1_20[211]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[101],stage1_22[105],stage1_21[143],stage1_20[212]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291], stage0_22[292], stage0_22[293]},
      {stage1_24[48],stage1_23[102],stage1_22[106],stage1_21[144],stage1_20[213]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[294], stage0_22[295], stage0_22[296], stage0_22[297], stage0_22[298], stage0_22[299]},
      {stage1_24[49],stage1_23[103],stage1_22[107],stage1_21[145],stage1_20[214]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[300], stage0_22[301], stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305]},
      {stage1_24[50],stage1_23[104],stage1_22[108],stage1_21[146],stage1_20[215]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[306], stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage1_24[51],stage1_23[105],stage1_22[109],stage1_21[147],stage1_20[216]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316], stage0_22[317]},
      {stage1_24[52],stage1_23[106],stage1_22[110],stage1_21[148],stage1_20[217]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321], stage0_22[322], stage0_22[323]},
      {stage1_24[53],stage1_23[107],stage1_22[111],stage1_21[149],stage1_20[218]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[324], stage0_22[325], stage0_22[326], stage0_22[327], stage0_22[328], stage0_22[329]},
      {stage1_24[54],stage1_23[108],stage1_22[112],stage1_21[150],stage1_20[219]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[330], stage0_22[331], stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335]},
      {stage1_24[55],stage1_23[109],stage1_22[113],stage1_21[151],stage1_20[220]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[336], stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage1_24[56],stage1_23[110],stage1_22[114],stage1_21[152],stage1_20[221]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346], stage0_22[347]},
      {stage1_24[57],stage1_23[111],stage1_22[115],stage1_21[153],stage1_20[222]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351], stage0_22[352], stage0_22[353]},
      {stage1_24[58],stage1_23[112],stage1_22[116],stage1_21[154],stage1_20[223]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[354], stage0_22[355], stage0_22[356], stage0_22[357], stage0_22[358], stage0_22[359]},
      {stage1_24[59],stage1_23[113],stage1_22[117],stage1_21[155],stage1_20[224]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[360], stage0_22[361], stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365]},
      {stage1_24[60],stage1_23[114],stage1_22[118],stage1_21[156],stage1_20[225]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[366], stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage1_24[61],stage1_23[115],stage1_22[119],stage1_21[157],stage1_20[226]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376], stage0_22[377]},
      {stage1_24[62],stage1_23[116],stage1_22[120],stage1_21[158],stage1_20[227]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381], stage0_22[382], stage0_22[383]},
      {stage1_24[63],stage1_23[117],stage1_22[121],stage1_21[159],stage1_20[228]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[384], stage0_22[385], stage0_22[386], stage0_22[387], stage0_22[388], stage0_22[389]},
      {stage1_24[64],stage1_23[118],stage1_22[122],stage1_21[160],stage1_20[229]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[390], stage0_22[391], stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395]},
      {stage1_24[65],stage1_23[119],stage1_22[123],stage1_21[161],stage1_20[230]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[396], stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage1_24[66],stage1_23[120],stage1_22[124],stage1_21[162],stage1_20[231]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage1_24[67],stage1_23[121],stage1_22[125],stage1_21[163],stage1_20[232]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412], stage0_22[413]},
      {stage1_24[68],stage1_23[122],stage1_22[126],stage1_21[164],stage1_20[233]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417], stage0_22[418], stage0_22[419]},
      {stage1_24[69],stage1_23[123],stage1_22[127],stage1_21[165],stage1_20[234]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[420], stage0_22[421], stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425]},
      {stage1_24[70],stage1_23[124],stage1_22[128],stage1_21[166],stage1_20[235]}
   );
   gpc606_5 gpc876 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[71],stage1_23[125],stage1_22[129],stage1_21[167]}
   );
   gpc606_5 gpc877 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[72],stage1_23[126],stage1_22[130],stage1_21[168]}
   );
   gpc606_5 gpc878 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[73],stage1_23[127],stage1_22[131],stage1_21[169]}
   );
   gpc606_5 gpc879 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[74],stage1_23[128],stage1_22[132],stage1_21[170]}
   );
   gpc606_5 gpc880 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[75],stage1_23[129],stage1_22[133],stage1_21[171]}
   );
   gpc606_5 gpc881 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[76],stage1_23[130],stage1_22[134],stage1_21[172]}
   );
   gpc606_5 gpc882 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[77],stage1_23[131],stage1_22[135],stage1_21[173]}
   );
   gpc606_5 gpc883 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[78],stage1_23[132],stage1_22[136],stage1_21[174]}
   );
   gpc606_5 gpc884 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[79],stage1_23[133],stage1_22[137],stage1_21[175]}
   );
   gpc606_5 gpc885 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[80],stage1_23[134],stage1_22[138],stage1_21[176]}
   );
   gpc606_5 gpc886 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[81],stage1_23[135],stage1_22[139],stage1_21[177]}
   );
   gpc606_5 gpc887 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[82],stage1_23[136],stage1_22[140],stage1_21[178]}
   );
   gpc606_5 gpc888 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[83],stage1_23[137],stage1_22[141],stage1_21[179]}
   );
   gpc606_5 gpc889 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[84],stage1_23[138],stage1_22[142],stage1_21[180]}
   );
   gpc606_5 gpc890 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[85],stage1_23[139],stage1_22[143],stage1_21[181]}
   );
   gpc606_5 gpc891 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[86],stage1_23[140],stage1_22[144],stage1_21[182]}
   );
   gpc606_5 gpc892 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[87],stage1_23[141],stage1_22[145],stage1_21[183]}
   );
   gpc606_5 gpc893 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[88],stage1_23[142],stage1_22[146],stage1_21[184]}
   );
   gpc606_5 gpc894 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[89],stage1_23[143],stage1_22[147],stage1_21[185]}
   );
   gpc606_5 gpc895 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[90],stage1_23[144],stage1_22[148],stage1_21[186]}
   );
   gpc606_5 gpc896 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[91],stage1_23[145],stage1_22[149],stage1_21[187]}
   );
   gpc606_5 gpc897 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[92],stage1_23[146],stage1_22[150],stage1_21[188]}
   );
   gpc606_5 gpc898 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[93],stage1_23[147],stage1_22[151],stage1_21[189]}
   );
   gpc606_5 gpc899 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[94],stage1_23[148],stage1_22[152],stage1_21[190]}
   );
   gpc606_5 gpc900 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[95],stage1_23[149],stage1_22[153],stage1_21[191]}
   );
   gpc606_5 gpc901 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[96],stage1_23[150],stage1_22[154],stage1_21[192]}
   );
   gpc606_5 gpc902 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[97],stage1_23[151],stage1_22[155],stage1_21[193]}
   );
   gpc606_5 gpc903 (
      {stage0_21[486], stage0_21[487], stage0_21[488], stage0_21[489], stage0_21[490], stage0_21[491]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[98],stage1_23[152],stage1_22[156],stage1_21[194]}
   );
   gpc606_5 gpc904 (
      {stage0_21[492], stage0_21[493], stage0_21[494], stage0_21[495], stage0_21[496], stage0_21[497]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[99],stage1_23[153],stage1_22[157],stage1_21[195]}
   );
   gpc606_5 gpc905 (
      {stage0_21[498], stage0_21[499], stage0_21[500], stage0_21[501], stage0_21[502], stage0_21[503]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[100],stage1_23[154],stage1_22[158],stage1_21[196]}
   );
   gpc615_5 gpc906 (
      {stage0_22[426], stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430]},
      {stage0_23[180]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[30],stage1_24[101],stage1_23[155],stage1_22[159]}
   );
   gpc615_5 gpc907 (
      {stage0_22[431], stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435]},
      {stage0_23[181]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[31],stage1_24[102],stage1_23[156],stage1_22[160]}
   );
   gpc615_5 gpc908 (
      {stage0_22[436], stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440]},
      {stage0_23[182]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[32],stage1_24[103],stage1_23[157],stage1_22[161]}
   );
   gpc615_5 gpc909 (
      {stage0_22[441], stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445]},
      {stage0_23[183]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[33],stage1_24[104],stage1_23[158],stage1_22[162]}
   );
   gpc615_5 gpc910 (
      {stage0_22[446], stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450]},
      {stage0_23[184]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[34],stage1_24[105],stage1_23[159],stage1_22[163]}
   );
   gpc615_5 gpc911 (
      {stage0_22[451], stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455]},
      {stage0_23[185]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[35],stage1_24[106],stage1_23[160],stage1_22[164]}
   );
   gpc615_5 gpc912 (
      {stage0_22[456], stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460]},
      {stage0_23[186]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[36],stage1_24[107],stage1_23[161],stage1_22[165]}
   );
   gpc615_5 gpc913 (
      {stage0_22[461], stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465]},
      {stage0_23[187]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[37],stage1_24[108],stage1_23[162],stage1_22[166]}
   );
   gpc615_5 gpc914 (
      {stage0_22[466], stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470]},
      {stage0_23[188]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[38],stage1_24[109],stage1_23[163],stage1_22[167]}
   );
   gpc615_5 gpc915 (
      {stage0_22[471], stage0_22[472], stage0_22[473], stage0_22[474], stage0_22[475]},
      {stage0_23[189]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[39],stage1_24[110],stage1_23[164],stage1_22[168]}
   );
   gpc615_5 gpc916 (
      {stage0_22[476], stage0_22[477], stage0_22[478], stage0_22[479], stage0_22[480]},
      {stage0_23[190]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[40],stage1_24[111],stage1_23[165],stage1_22[169]}
   );
   gpc606_5 gpc917 (
      {stage0_23[191], stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[11],stage1_25[41],stage1_24[112],stage1_23[166]}
   );
   gpc606_5 gpc918 (
      {stage0_23[197], stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[12],stage1_25[42],stage1_24[113],stage1_23[167]}
   );
   gpc606_5 gpc919 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[13],stage1_25[43],stage1_24[114],stage1_23[168]}
   );
   gpc606_5 gpc920 (
      {stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[14],stage1_25[44],stage1_24[115],stage1_23[169]}
   );
   gpc606_5 gpc921 (
      {stage0_23[215], stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[15],stage1_25[45],stage1_24[116],stage1_23[170]}
   );
   gpc606_5 gpc922 (
      {stage0_23[221], stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[16],stage1_25[46],stage1_24[117],stage1_23[171]}
   );
   gpc606_5 gpc923 (
      {stage0_23[227], stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[17],stage1_25[47],stage1_24[118],stage1_23[172]}
   );
   gpc606_5 gpc924 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[18],stage1_25[48],stage1_24[119],stage1_23[173]}
   );
   gpc606_5 gpc925 (
      {stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[19],stage1_25[49],stage1_24[120],stage1_23[174]}
   );
   gpc606_5 gpc926 (
      {stage0_23[245], stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[20],stage1_25[50],stage1_24[121],stage1_23[175]}
   );
   gpc606_5 gpc927 (
      {stage0_23[251], stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[21],stage1_25[51],stage1_24[122],stage1_23[176]}
   );
   gpc606_5 gpc928 (
      {stage0_23[257], stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[22],stage1_25[52],stage1_24[123],stage1_23[177]}
   );
   gpc606_5 gpc929 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[23],stage1_25[53],stage1_24[124],stage1_23[178]}
   );
   gpc606_5 gpc930 (
      {stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[24],stage1_25[54],stage1_24[125],stage1_23[179]}
   );
   gpc606_5 gpc931 (
      {stage0_23[275], stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[25],stage1_25[55],stage1_24[126],stage1_23[180]}
   );
   gpc606_5 gpc932 (
      {stage0_23[281], stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[26],stage1_25[56],stage1_24[127],stage1_23[181]}
   );
   gpc606_5 gpc933 (
      {stage0_23[287], stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[27],stage1_25[57],stage1_24[128],stage1_23[182]}
   );
   gpc606_5 gpc934 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[28],stage1_25[58],stage1_24[129],stage1_23[183]}
   );
   gpc606_5 gpc935 (
      {stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[29],stage1_25[59],stage1_24[130],stage1_23[184]}
   );
   gpc606_5 gpc936 (
      {stage0_23[305], stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[30],stage1_25[60],stage1_24[131],stage1_23[185]}
   );
   gpc606_5 gpc937 (
      {stage0_23[311], stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[31],stage1_25[61],stage1_24[132],stage1_23[186]}
   );
   gpc606_5 gpc938 (
      {stage0_23[317], stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[32],stage1_25[62],stage1_24[133],stage1_23[187]}
   );
   gpc606_5 gpc939 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[33],stage1_25[63],stage1_24[134],stage1_23[188]}
   );
   gpc606_5 gpc940 (
      {stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[34],stage1_25[64],stage1_24[135],stage1_23[189]}
   );
   gpc606_5 gpc941 (
      {stage0_23[335], stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[35],stage1_25[65],stage1_24[136],stage1_23[190]}
   );
   gpc606_5 gpc942 (
      {stage0_23[341], stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[36],stage1_25[66],stage1_24[137],stage1_23[191]}
   );
   gpc606_5 gpc943 (
      {stage0_23[347], stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[37],stage1_25[67],stage1_24[138],stage1_23[192]}
   );
   gpc606_5 gpc944 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[38],stage1_25[68],stage1_24[139],stage1_23[193]}
   );
   gpc606_5 gpc945 (
      {stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[39],stage1_25[69],stage1_24[140],stage1_23[194]}
   );
   gpc606_5 gpc946 (
      {stage0_23[365], stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[40],stage1_25[70],stage1_24[141],stage1_23[195]}
   );
   gpc606_5 gpc947 (
      {stage0_23[371], stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[41],stage1_25[71],stage1_24[142],stage1_23[196]}
   );
   gpc606_5 gpc948 (
      {stage0_23[377], stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[42],stage1_25[72],stage1_24[143],stage1_23[197]}
   );
   gpc615_5 gpc949 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[66]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[43],stage1_25[73],stage1_24[144],stage1_23[198]}
   );
   gpc615_5 gpc950 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[67]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[44],stage1_25[74],stage1_24[145],stage1_23[199]}
   );
   gpc615_5 gpc951 (
      {stage0_23[393], stage0_23[394], stage0_23[395], stage0_23[396], stage0_23[397]},
      {stage0_24[68]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[45],stage1_25[75],stage1_24[146],stage1_23[200]}
   );
   gpc615_5 gpc952 (
      {stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401], stage0_23[402]},
      {stage0_24[69]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[46],stage1_25[76],stage1_24[147],stage1_23[201]}
   );
   gpc615_5 gpc953 (
      {stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage0_24[70]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[47],stage1_25[77],stage1_24[148],stage1_23[202]}
   );
   gpc615_5 gpc954 (
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412]},
      {stage0_24[71]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[48],stage1_25[78],stage1_24[149],stage1_23[203]}
   );
   gpc615_5 gpc955 (
      {stage0_23[413], stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417]},
      {stage0_24[72]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[49],stage1_25[79],stage1_24[150],stage1_23[204]}
   );
   gpc606_5 gpc956 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[39],stage1_26[50],stage1_25[80],stage1_24[151]}
   );
   gpc606_5 gpc957 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[40],stage1_26[51],stage1_25[81],stage1_24[152]}
   );
   gpc606_5 gpc958 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[41],stage1_26[52],stage1_25[82],stage1_24[153]}
   );
   gpc606_5 gpc959 (
      {stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[42],stage1_26[53],stage1_25[83],stage1_24[154]}
   );
   gpc606_5 gpc960 (
      {stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[43],stage1_26[54],stage1_25[84],stage1_24[155]}
   );
   gpc606_5 gpc961 (
      {stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[44],stage1_26[55],stage1_25[85],stage1_24[156]}
   );
   gpc606_5 gpc962 (
      {stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113], stage0_24[114]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[45],stage1_26[56],stage1_25[86],stage1_24[157]}
   );
   gpc606_5 gpc963 (
      {stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119], stage0_24[120]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[46],stage1_26[57],stage1_25[87],stage1_24[158]}
   );
   gpc606_5 gpc964 (
      {stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125], stage0_24[126]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[47],stage1_26[58],stage1_25[88],stage1_24[159]}
   );
   gpc606_5 gpc965 (
      {stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131], stage0_24[132]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[48],stage1_26[59],stage1_25[89],stage1_24[160]}
   );
   gpc606_5 gpc966 (
      {stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137], stage0_24[138]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[49],stage1_26[60],stage1_25[90],stage1_24[161]}
   );
   gpc606_5 gpc967 (
      {stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143], stage0_24[144]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[50],stage1_26[61],stage1_25[91],stage1_24[162]}
   );
   gpc606_5 gpc968 (
      {stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149], stage0_24[150]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[51],stage1_26[62],stage1_25[92],stage1_24[163]}
   );
   gpc606_5 gpc969 (
      {stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155], stage0_24[156]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[52],stage1_26[63],stage1_25[93],stage1_24[164]}
   );
   gpc606_5 gpc970 (
      {stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161], stage0_24[162]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[53],stage1_26[64],stage1_25[94],stage1_24[165]}
   );
   gpc606_5 gpc971 (
      {stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167], stage0_24[168]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[54],stage1_26[65],stage1_25[95],stage1_24[166]}
   );
   gpc606_5 gpc972 (
      {stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172], stage0_24[173], stage0_24[174]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[55],stage1_26[66],stage1_25[96],stage1_24[167]}
   );
   gpc606_5 gpc973 (
      {stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178], stage0_24[179], stage0_24[180]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[56],stage1_26[67],stage1_25[97],stage1_24[168]}
   );
   gpc606_5 gpc974 (
      {stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184], stage0_24[185], stage0_24[186]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[57],stage1_26[68],stage1_25[98],stage1_24[169]}
   );
   gpc606_5 gpc975 (
      {stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190], stage0_24[191], stage0_24[192]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[58],stage1_26[69],stage1_25[99],stage1_24[170]}
   );
   gpc606_5 gpc976 (
      {stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196], stage0_24[197], stage0_24[198]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[59],stage1_26[70],stage1_25[100],stage1_24[171]}
   );
   gpc606_5 gpc977 (
      {stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[60],stage1_26[71],stage1_25[101],stage1_24[172]}
   );
   gpc606_5 gpc978 (
      {stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[61],stage1_26[72],stage1_25[102],stage1_24[173]}
   );
   gpc606_5 gpc979 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215], stage0_24[216]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[62],stage1_26[73],stage1_25[103],stage1_24[174]}
   );
   gpc606_5 gpc980 (
      {stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220], stage0_24[221], stage0_24[222]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[63],stage1_26[74],stage1_25[104],stage1_24[175]}
   );
   gpc606_5 gpc981 (
      {stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226], stage0_24[227], stage0_24[228]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[64],stage1_26[75],stage1_25[105],stage1_24[176]}
   );
   gpc606_5 gpc982 (
      {stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[65],stage1_26[76],stage1_25[106],stage1_24[177]}
   );
   gpc606_5 gpc983 (
      {stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[66],stage1_26[77],stage1_25[107],stage1_24[178]}
   );
   gpc606_5 gpc984 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245], stage0_24[246]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[67],stage1_26[78],stage1_25[108],stage1_24[179]}
   );
   gpc606_5 gpc985 (
      {stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250], stage0_24[251], stage0_24[252]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[68],stage1_26[79],stage1_25[109],stage1_24[180]}
   );
   gpc606_5 gpc986 (
      {stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256], stage0_24[257], stage0_24[258]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[69],stage1_26[80],stage1_25[110],stage1_24[181]}
   );
   gpc606_5 gpc987 (
      {stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[70],stage1_26[81],stage1_25[111],stage1_24[182]}
   );
   gpc606_5 gpc988 (
      {stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[71],stage1_26[82],stage1_25[112],stage1_24[183]}
   );
   gpc606_5 gpc989 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275], stage0_24[276]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[72],stage1_26[83],stage1_25[113],stage1_24[184]}
   );
   gpc606_5 gpc990 (
      {stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280], stage0_24[281], stage0_24[282]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[73],stage1_26[84],stage1_25[114],stage1_24[185]}
   );
   gpc606_5 gpc991 (
      {stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286], stage0_24[287], stage0_24[288]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[74],stage1_26[85],stage1_25[115],stage1_24[186]}
   );
   gpc606_5 gpc992 (
      {stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[75],stage1_26[86],stage1_25[116],stage1_24[187]}
   );
   gpc606_5 gpc993 (
      {stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[76],stage1_26[87],stage1_25[117],stage1_24[188]}
   );
   gpc606_5 gpc994 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305], stage0_24[306]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[77],stage1_26[88],stage1_25[118],stage1_24[189]}
   );
   gpc606_5 gpc995 (
      {stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310], stage0_24[311], stage0_24[312]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[78],stage1_26[89],stage1_25[119],stage1_24[190]}
   );
   gpc606_5 gpc996 (
      {stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316], stage0_24[317], stage0_24[318]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[79],stage1_26[90],stage1_25[120],stage1_24[191]}
   );
   gpc606_5 gpc997 (
      {stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[80],stage1_26[91],stage1_25[121],stage1_24[192]}
   );
   gpc606_5 gpc998 (
      {stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[81],stage1_26[92],stage1_25[122],stage1_24[193]}
   );
   gpc606_5 gpc999 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335], stage0_24[336]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[82],stage1_26[93],stage1_25[123],stage1_24[194]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340], stage0_24[341], stage0_24[342]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[83],stage1_26[94],stage1_25[124],stage1_24[195]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346], stage0_24[347], stage0_24[348]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[84],stage1_26[95],stage1_25[125],stage1_24[196]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[85],stage1_26[96],stage1_25[126],stage1_24[197]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[86],stage1_26[97],stage1_25[127],stage1_24[198]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[87],stage1_26[98],stage1_25[128],stage1_24[199]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371], stage0_24[372]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[88],stage1_26[99],stage1_25[129],stage1_24[200]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376], stage0_24[377], stage0_24[378]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[89],stage1_26[100],stage1_25[130],stage1_24[201]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[90],stage1_26[101],stage1_25[131],stage1_24[202]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[91],stage1_26[102],stage1_25[132],stage1_24[203]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[92],stage1_26[103],stage1_25[133],stage1_24[204]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401], stage0_24[402]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[93],stage1_26[104],stage1_25[134],stage1_24[205]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406], stage0_24[407], stage0_24[408]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[94],stage1_26[105],stage1_25[135],stage1_24[206]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[95],stage1_26[106],stage1_25[136],stage1_24[207]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[96],stage1_26[107],stage1_25[137],stage1_24[208]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[97],stage1_26[108],stage1_25[138],stage1_24[209]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431], stage0_24[432]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[98],stage1_26[109],stage1_25[139],stage1_24[210]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436], stage0_24[437], stage0_24[438]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[99],stage1_26[110],stage1_25[140],stage1_24[211]}
   );
   gpc606_5 gpc1017 (
      {stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[100],stage1_26[111],stage1_25[141],stage1_24[212]}
   );
   gpc606_5 gpc1018 (
      {stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[101],stage1_26[112],stage1_25[142],stage1_24[213]}
   );
   gpc606_5 gpc1019 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[102],stage1_26[113],stage1_25[143],stage1_24[214]}
   );
   gpc606_5 gpc1020 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461], stage0_24[462]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[103],stage1_26[114],stage1_25[144],stage1_24[215]}
   );
   gpc606_5 gpc1021 (
      {stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466], stage0_24[467], stage0_24[468]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[104],stage1_26[115],stage1_25[145],stage1_24[216]}
   );
   gpc606_5 gpc1022 (
      {stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[105],stage1_26[116],stage1_25[146],stage1_24[217]}
   );
   gpc606_5 gpc1023 (
      {stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[106],stage1_26[117],stage1_25[147],stage1_24[218]}
   );
   gpc606_5 gpc1024 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[107],stage1_26[118],stage1_25[148],stage1_24[219]}
   );
   gpc606_5 gpc1025 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491], stage0_24[492]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[108],stage1_26[119],stage1_25[149],stage1_24[220]}
   );
   gpc606_5 gpc1026 (
      {stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496], stage0_24[497], stage0_24[498]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[109],stage1_26[120],stage1_25[150],stage1_24[221]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[71],stage1_27[110],stage1_26[121],stage1_25[151]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[72],stage1_27[111],stage1_26[122],stage1_25[152]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[426]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[73],stage1_27[112],stage1_26[123],stage1_25[153]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[427]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[74],stage1_27[113],stage1_26[124],stage1_25[154]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[428]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[75],stage1_27[114],stage1_26[125],stage1_25[155]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[429]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[76],stage1_27[115],stage1_26[126],stage1_25[156]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[430]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[77],stage1_27[116],stage1_26[127],stage1_25[157]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[431]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[78],stage1_27[117],stage1_26[128],stage1_25[158]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[432]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[79],stage1_27[118],stage1_26[129],stage1_25[159]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[433]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[80],stage1_27[119],stage1_26[130],stage1_25[160]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[434]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[81],stage1_27[120],stage1_26[131],stage1_25[161]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[435]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[82],stage1_27[121],stage1_26[132],stage1_25[162]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[436]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[83],stage1_27[122],stage1_26[133],stage1_25[163]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[437]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[84],stage1_27[123],stage1_26[134],stage1_25[164]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[438]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[85],stage1_27[124],stage1_26[135],stage1_25[165]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[439]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[86],stage1_27[125],stage1_26[136],stage1_25[166]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[440]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[87],stage1_27[126],stage1_26[137],stage1_25[167]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[441]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[88],stage1_27[127],stage1_26[138],stage1_25[168]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[442]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[89],stage1_27[128],stage1_26[139],stage1_25[169]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[443]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[90],stage1_27[129],stage1_26[140],stage1_25[170]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[444]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[91],stage1_27[130],stage1_26[141],stage1_25[171]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[445]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[92],stage1_27[131],stage1_26[142],stage1_25[172]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[446]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[93],stage1_27[132],stage1_26[143],stage1_25[173]}
   );
   gpc615_5 gpc1050 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[447]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[94],stage1_27[133],stage1_26[144],stage1_25[174]}
   );
   gpc615_5 gpc1051 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[448]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[95],stage1_27[134],stage1_26[145],stage1_25[175]}
   );
   gpc615_5 gpc1052 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[449]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[96],stage1_27[135],stage1_26[146],stage1_25[176]}
   );
   gpc615_5 gpc1053 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[450]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[97],stage1_27[136],stage1_26[147],stage1_25[177]}
   );
   gpc615_5 gpc1054 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[451]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[98],stage1_27[137],stage1_26[148],stage1_25[178]}
   );
   gpc615_5 gpc1055 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[452]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[99],stage1_27[138],stage1_26[149],stage1_25[179]}
   );
   gpc615_5 gpc1056 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[453]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[100],stage1_27[139],stage1_26[150],stage1_25[180]}
   );
   gpc615_5 gpc1057 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[454]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[101],stage1_27[140],stage1_26[151],stage1_25[181]}
   );
   gpc615_5 gpc1058 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[455]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[102],stage1_27[141],stage1_26[152],stage1_25[182]}
   );
   gpc615_5 gpc1059 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[456]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[103],stage1_27[142],stage1_26[153],stage1_25[183]}
   );
   gpc615_5 gpc1060 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[457]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[104],stage1_27[143],stage1_26[154],stage1_25[184]}
   );
   gpc615_5 gpc1061 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[458]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[105],stage1_27[144],stage1_26[155],stage1_25[185]}
   );
   gpc615_5 gpc1062 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[459]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[106],stage1_27[145],stage1_26[156],stage1_25[186]}
   );
   gpc615_5 gpc1063 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[460]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[107],stage1_27[146],stage1_26[157],stage1_25[187]}
   );
   gpc615_5 gpc1064 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[461]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[108],stage1_27[147],stage1_26[158],stage1_25[188]}
   );
   gpc615_5 gpc1065 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[462]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[109],stage1_27[148],stage1_26[159],stage1_25[189]}
   );
   gpc615_5 gpc1066 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[463]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[110],stage1_27[149],stage1_26[160],stage1_25[190]}
   );
   gpc615_5 gpc1067 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[464]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[111],stage1_27[150],stage1_26[161],stage1_25[191]}
   );
   gpc615_5 gpc1068 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[465]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[112],stage1_27[151],stage1_26[162],stage1_25[192]}
   );
   gpc615_5 gpc1069 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[466]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[113],stage1_27[152],stage1_26[163],stage1_25[193]}
   );
   gpc615_5 gpc1070 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[467]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[114],stage1_27[153],stage1_26[164],stage1_25[194]}
   );
   gpc615_5 gpc1071 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[468]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[115],stage1_27[154],stage1_26[165],stage1_25[195]}
   );
   gpc615_5 gpc1072 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[469]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[116],stage1_27[155],stage1_26[166],stage1_25[196]}
   );
   gpc615_5 gpc1073 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[470]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[117],stage1_27[156],stage1_26[167],stage1_25[197]}
   );
   gpc615_5 gpc1074 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[471]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[118],stage1_27[157],stage1_26[168],stage1_25[198]}
   );
   gpc615_5 gpc1075 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[472]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[119],stage1_27[158],stage1_26[169],stage1_25[199]}
   );
   gpc615_5 gpc1076 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[473]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[120],stage1_27[159],stage1_26[170],stage1_25[200]}
   );
   gpc615_5 gpc1077 (
      {stage0_25[486], stage0_25[487], stage0_25[488], stage0_25[489], stage0_25[490]},
      {stage0_26[474]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[121],stage1_27[160],stage1_26[171],stage1_25[201]}
   );
   gpc615_5 gpc1078 (
      {stage0_25[491], stage0_25[492], stage0_25[493], stage0_25[494], stage0_25[495]},
      {stage0_26[475]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[122],stage1_27[161],stage1_26[172],stage1_25[202]}
   );
   gpc615_5 gpc1079 (
      {stage0_25[496], stage0_25[497], stage0_25[498], stage0_25[499], stage0_25[500]},
      {stage0_26[476]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[123],stage1_27[162],stage1_26[173],stage1_25[203]}
   );
   gpc615_5 gpc1080 (
      {stage0_25[501], stage0_25[502], stage0_25[503], stage0_25[504], stage0_25[505]},
      {stage0_26[477]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[124],stage1_27[163],stage1_26[174],stage1_25[204]}
   );
   gpc615_5 gpc1081 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[324]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[54],stage1_28[125],stage1_27[164],stage1_26[175]}
   );
   gpc615_5 gpc1082 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[325]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[55],stage1_28[126],stage1_27[165],stage1_26[176]}
   );
   gpc615_5 gpc1083 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[326]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[56],stage1_28[127],stage1_27[166],stage1_26[177]}
   );
   gpc615_5 gpc1084 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[327]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[57],stage1_28[128],stage1_27[167],stage1_26[178]}
   );
   gpc615_5 gpc1085 (
      {stage0_26[498], stage0_26[499], stage0_26[500], stage0_26[501], stage0_26[502]},
      {stage0_27[328]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[58],stage1_28[129],stage1_27[168],stage1_26[179]}
   );
   gpc7_3 gpc1086 (
      {stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[59],stage1_28[130],stage1_27[169]}
   );
   gpc7_3 gpc1087 (
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage1_29[60],stage1_28[131],stage1_27[170]}
   );
   gpc615_5 gpc1088 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[30]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[61],stage1_28[132],stage1_27[171]}
   );
   gpc615_5 gpc1089 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[31]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[62],stage1_28[133],stage1_27[172]}
   );
   gpc615_5 gpc1090 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[32]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[63],stage1_28[134],stage1_27[173]}
   );
   gpc615_5 gpc1091 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[33]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[64],stage1_28[135],stage1_27[174]}
   );
   gpc615_5 gpc1092 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[34]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[65],stage1_28[136],stage1_27[175]}
   );
   gpc615_5 gpc1093 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[35]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[66],stage1_28[137],stage1_27[176]}
   );
   gpc615_5 gpc1094 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[36]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[67],stage1_28[138],stage1_27[177]}
   );
   gpc615_5 gpc1095 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[37]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[68],stage1_28[139],stage1_27[178]}
   );
   gpc615_5 gpc1096 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[38]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[69],stage1_28[140],stage1_27[179]}
   );
   gpc615_5 gpc1097 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[39]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[70],stage1_28[141],stage1_27[180]}
   );
   gpc615_5 gpc1098 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[40]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[15],stage1_29[71],stage1_28[142],stage1_27[181]}
   );
   gpc615_5 gpc1099 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[41]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[16],stage1_29[72],stage1_28[143],stage1_27[182]}
   );
   gpc615_5 gpc1100 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[42]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[17],stage1_29[73],stage1_28[144],stage1_27[183]}
   );
   gpc615_5 gpc1101 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[43]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[18],stage1_29[74],stage1_28[145],stage1_27[184]}
   );
   gpc615_5 gpc1102 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[44]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[19],stage1_29[75],stage1_28[146],stage1_27[185]}
   );
   gpc615_5 gpc1103 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[45]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[20],stage1_29[76],stage1_28[147],stage1_27[186]}
   );
   gpc615_5 gpc1104 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[46]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[21],stage1_29[77],stage1_28[148],stage1_27[187]}
   );
   gpc615_5 gpc1105 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[47]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[22],stage1_29[78],stage1_28[149],stage1_27[188]}
   );
   gpc615_5 gpc1106 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[48]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[23],stage1_29[79],stage1_28[150],stage1_27[189]}
   );
   gpc615_5 gpc1107 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[49]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[24],stage1_29[80],stage1_28[151],stage1_27[190]}
   );
   gpc615_5 gpc1108 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[50]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[25],stage1_29[81],stage1_28[152],stage1_27[191]}
   );
   gpc615_5 gpc1109 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[51]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[26],stage1_29[82],stage1_28[153],stage1_27[192]}
   );
   gpc615_5 gpc1110 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[52]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[27],stage1_29[83],stage1_28[154],stage1_27[193]}
   );
   gpc615_5 gpc1111 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[53]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[28],stage1_29[84],stage1_28[155],stage1_27[194]}
   );
   gpc615_5 gpc1112 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[54]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[29],stage1_29[85],stage1_28[156],stage1_27[195]}
   );
   gpc615_5 gpc1113 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[55]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[30],stage1_29[86],stage1_28[157],stage1_27[196]}
   );
   gpc615_5 gpc1114 (
      {stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477]},
      {stage0_28[56]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[31],stage1_29[87],stage1_28[158],stage1_27[197]}
   );
   gpc615_5 gpc1115 (
      {stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_28[57]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[32],stage1_29[88],stage1_28[159],stage1_27[198]}
   );
   gpc615_5 gpc1116 (
      {stage0_27[483], stage0_27[484], stage0_27[485], stage0_27[486], stage0_27[487]},
      {stage0_28[58]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[33],stage1_29[89],stage1_28[160],stage1_27[199]}
   );
   gpc615_5 gpc1117 (
      {stage0_27[488], stage0_27[489], stage0_27[490], stage0_27[491], stage0_27[492]},
      {stage0_28[59]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[34],stage1_29[90],stage1_28[161],stage1_27[200]}
   );
   gpc615_5 gpc1118 (
      {stage0_27[493], stage0_27[494], stage0_27[495], stage0_27[496], stage0_27[497]},
      {stage0_28[60]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[35],stage1_29[91],stage1_28[162],stage1_27[201]}
   );
   gpc615_5 gpc1119 (
      {stage0_27[498], stage0_27[499], stage0_27[500], stage0_27[501], stage0_27[502]},
      {stage0_28[61]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[36],stage1_29[92],stage1_28[163],stage1_27[202]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65], stage0_28[66], stage0_28[67]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[32],stage1_30[37],stage1_29[93],stage1_28[164]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71], stage0_28[72], stage0_28[73]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[33],stage1_30[38],stage1_29[94],stage1_28[165]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78], stage0_28[79]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[34],stage1_30[39],stage1_29[95],stage1_28[166]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84], stage0_28[85]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[35],stage1_30[40],stage1_29[96],stage1_28[167]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90], stage0_28[91]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[36],stage1_30[41],stage1_29[97],stage1_28[168]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[37],stage1_30[42],stage1_29[98],stage1_28[169]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[38],stage1_30[43],stage1_29[99],stage1_28[170]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[39],stage1_30[44],stage1_29[100],stage1_28[171]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[40],stage1_30[45],stage1_29[101],stage1_28[172]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[41],stage1_30[46],stage1_29[102],stage1_28[173]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[42],stage1_30[47],stage1_29[103],stage1_28[174]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[43],stage1_30[48],stage1_29[104],stage1_28[175]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[44],stage1_30[49],stage1_29[105],stage1_28[176]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144], stage0_28[145]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[45],stage1_30[50],stage1_29[106],stage1_28[177]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150], stage0_28[151]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[46],stage1_30[51],stage1_29[107],stage1_28[178]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156], stage0_28[157]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[47],stage1_30[52],stage1_29[108],stage1_28[179]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162], stage0_28[163]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[48],stage1_30[53],stage1_29[109],stage1_28[180]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168], stage0_28[169]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[49],stage1_30[54],stage1_29[110],stage1_28[181]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174], stage0_28[175]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[50],stage1_30[55],stage1_29[111],stage1_28[182]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180], stage0_28[181]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[51],stage1_30[56],stage1_29[112],stage1_28[183]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186], stage0_28[187]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[52],stage1_30[57],stage1_29[113],stage1_28[184]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192], stage0_28[193]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[53],stage1_30[58],stage1_29[114],stage1_28[185]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198], stage0_28[199]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[54],stage1_30[59],stage1_29[115],stage1_28[186]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204], stage0_28[205]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[55],stage1_30[60],stage1_29[116],stage1_28[187]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210], stage0_28[211]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[56],stage1_30[61],stage1_29[117],stage1_28[188]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216], stage0_28[217]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[57],stage1_30[62],stage1_29[118],stage1_28[189]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222], stage0_28[223]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[58],stage1_30[63],stage1_29[119],stage1_28[190]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228], stage0_28[229]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[59],stage1_30[64],stage1_29[120],stage1_28[191]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234], stage0_28[235]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[60],stage1_30[65],stage1_29[121],stage1_28[192]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240], stage0_28[241]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[61],stage1_30[66],stage1_29[122],stage1_28[193]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246], stage0_28[247]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[62],stage1_30[67],stage1_29[123],stage1_28[194]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252], stage0_28[253]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[63],stage1_30[68],stage1_29[124],stage1_28[195]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258], stage0_28[259]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[64],stage1_30[69],stage1_29[125],stage1_28[196]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264], stage0_28[265]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[65],stage1_30[70],stage1_29[126],stage1_28[197]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270], stage0_28[271]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[66],stage1_30[71],stage1_29[127],stage1_28[198]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276], stage0_28[277]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[67],stage1_30[72],stage1_29[128],stage1_28[199]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282], stage0_28[283]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[68],stage1_30[73],stage1_29[129],stage1_28[200]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288], stage0_28[289]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[69],stage1_30[74],stage1_29[130],stage1_28[201]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294], stage0_28[295]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[70],stage1_30[75],stage1_29[131],stage1_28[202]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300], stage0_28[301]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[71],stage1_30[76],stage1_29[132],stage1_28[203]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306], stage0_28[307]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[72],stage1_30[77],stage1_29[133],stage1_28[204]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312], stage0_28[313]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[73],stage1_30[78],stage1_29[134],stage1_28[205]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[74],stage1_30[79],stage1_29[135],stage1_28[206]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[75],stage1_30[80],stage1_29[136],stage1_28[207]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330], stage0_28[331]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[76],stage1_30[81],stage1_29[137],stage1_28[208]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336], stage0_28[337]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[77],stage1_30[82],stage1_29[138],stage1_28[209]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342], stage0_28[343]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[78],stage1_30[83],stage1_29[139],stage1_28[210]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[79],stage1_30[84],stage1_29[140],stage1_28[211]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[80],stage1_30[85],stage1_29[141],stage1_28[212]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360], stage0_28[361]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[81],stage1_30[86],stage1_29[142],stage1_28[213]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366], stage0_28[367]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[82],stage1_30[87],stage1_29[143],stage1_28[214]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372], stage0_28[373]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[83],stage1_30[88],stage1_29[144],stage1_28[215]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[84],stage1_30[89],stage1_29[145],stage1_28[216]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[85],stage1_30[90],stage1_29[146],stage1_28[217]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390], stage0_28[391]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[86],stage1_30[91],stage1_29[147],stage1_28[218]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396], stage0_28[397]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[87],stage1_30[92],stage1_29[148],stage1_28[219]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402], stage0_28[403]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[88],stage1_30[93],stage1_29[149],stage1_28[220]}
   );
   gpc606_5 gpc1177 (
      {stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[89],stage1_30[94],stage1_29[150],stage1_28[221]}
   );
   gpc606_5 gpc1178 (
      {stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[90],stage1_30[95],stage1_29[151],stage1_28[222]}
   );
   gpc606_5 gpc1179 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420], stage0_28[421]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[91],stage1_30[96],stage1_29[152],stage1_28[223]}
   );
   gpc606_5 gpc1180 (
      {stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426], stage0_28[427]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[92],stage1_30[97],stage1_29[153],stage1_28[224]}
   );
   gpc606_5 gpc1181 (
      {stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432], stage0_28[433]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[93],stage1_30[98],stage1_29[154],stage1_28[225]}
   );
   gpc606_5 gpc1182 (
      {stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[94],stage1_30[99],stage1_29[155],stage1_28[226]}
   );
   gpc606_5 gpc1183 (
      {stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[95],stage1_30[100],stage1_29[156],stage1_28[227]}
   );
   gpc606_5 gpc1184 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450], stage0_28[451]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[96],stage1_30[101],stage1_29[157],stage1_28[228]}
   );
   gpc606_5 gpc1185 (
      {stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456], stage0_28[457]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[97],stage1_30[102],stage1_29[158],stage1_28[229]}
   );
   gpc606_5 gpc1186 (
      {stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462], stage0_28[463]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[98],stage1_30[103],stage1_29[159],stage1_28[230]}
   );
   gpc606_5 gpc1187 (
      {stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[99],stage1_30[104],stage1_29[160],stage1_28[231]}
   );
   gpc606_5 gpc1188 (
      {stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[100],stage1_30[105],stage1_29[161],stage1_28[232]}
   );
   gpc606_5 gpc1189 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480], stage0_28[481]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[101],stage1_30[106],stage1_29[162],stage1_28[233]}
   );
   gpc606_5 gpc1190 (
      {stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485], stage0_28[486], stage0_28[487]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[102],stage1_30[107],stage1_29[163],stage1_28[234]}
   );
   gpc606_5 gpc1191 (
      {stage0_28[488], stage0_28[489], stage0_28[490], stage0_28[491], stage0_28[492], stage0_28[493]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[103],stage1_30[108],stage1_29[164],stage1_28[235]}
   );
   gpc606_5 gpc1192 (
      {stage0_28[494], stage0_28[495], stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[104],stage1_30[109],stage1_29[165],stage1_28[236]}
   );
   gpc606_5 gpc1193 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[73],stage1_31[105],stage1_30[110],stage1_29[166]}
   );
   gpc606_5 gpc1194 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[74],stage1_31[106],stage1_30[111],stage1_29[167]}
   );
   gpc606_5 gpc1195 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[75],stage1_31[107],stage1_30[112],stage1_29[168]}
   );
   gpc606_5 gpc1196 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[76],stage1_31[108],stage1_30[113],stage1_29[169]}
   );
   gpc606_5 gpc1197 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[77],stage1_31[109],stage1_30[114],stage1_29[170]}
   );
   gpc606_5 gpc1198 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[78],stage1_31[110],stage1_30[115],stage1_29[171]}
   );
   gpc606_5 gpc1199 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[79],stage1_31[111],stage1_30[116],stage1_29[172]}
   );
   gpc606_5 gpc1200 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[80],stage1_31[112],stage1_30[117],stage1_29[173]}
   );
   gpc606_5 gpc1201 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[81],stage1_31[113],stage1_30[118],stage1_29[174]}
   );
   gpc606_5 gpc1202 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[82],stage1_31[114],stage1_30[119],stage1_29[175]}
   );
   gpc606_5 gpc1203 (
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[83],stage1_31[115],stage1_30[120],stage1_29[176]}
   );
   gpc606_5 gpc1204 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[84],stage1_31[116],stage1_30[121],stage1_29[177]}
   );
   gpc606_5 gpc1205 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[85],stage1_31[117],stage1_30[122],stage1_29[178]}
   );
   gpc606_5 gpc1206 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[86],stage1_31[118],stage1_30[123],stage1_29[179]}
   );
   gpc606_5 gpc1207 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[87],stage1_31[119],stage1_30[124],stage1_29[180]}
   );
   gpc606_5 gpc1208 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[88],stage1_31[120],stage1_30[125],stage1_29[181]}
   );
   gpc606_5 gpc1209 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[89],stage1_31[121],stage1_30[126],stage1_29[182]}
   );
   gpc606_5 gpc1210 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[90],stage1_31[122],stage1_30[127],stage1_29[183]}
   );
   gpc606_5 gpc1211 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[91],stage1_31[123],stage1_30[128],stage1_29[184]}
   );
   gpc606_5 gpc1212 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[92],stage1_31[124],stage1_30[129],stage1_29[185]}
   );
   gpc606_5 gpc1213 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[93],stage1_31[125],stage1_30[130],stage1_29[186]}
   );
   gpc606_5 gpc1214 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[94],stage1_31[126],stage1_30[131],stage1_29[187]}
   );
   gpc606_5 gpc1215 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[95],stage1_31[127],stage1_30[132],stage1_29[188]}
   );
   gpc606_5 gpc1216 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[96],stage1_31[128],stage1_30[133],stage1_29[189]}
   );
   gpc606_5 gpc1217 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[97],stage1_31[129],stage1_30[134],stage1_29[190]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[98],stage1_31[130],stage1_30[135],stage1_29[191]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[99],stage1_31[131],stage1_30[136],stage1_29[192]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[100],stage1_31[132],stage1_30[137],stage1_29[193]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[101],stage1_31[133],stage1_30[138],stage1_29[194]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[102],stage1_31[134],stage1_30[139],stage1_29[195]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[103],stage1_31[135],stage1_30[140],stage1_29[196]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[104],stage1_31[136],stage1_30[141],stage1_29[197]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[105],stage1_31[137],stage1_30[142],stage1_29[198]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[106],stage1_31[138],stage1_30[143],stage1_29[199]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[107],stage1_31[139],stage1_30[144],stage1_29[200]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[108],stage1_31[140],stage1_30[145],stage1_29[201]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[109],stage1_31[141],stage1_30[146],stage1_29[202]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[110],stage1_31[142],stage1_30[147],stage1_29[203]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[111],stage1_31[143],stage1_30[148],stage1_29[204]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[112],stage1_31[144],stage1_30[149],stage1_29[205]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[113],stage1_31[145],stage1_30[150],stage1_29[206]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[114],stage1_31[146],stage1_30[151],stage1_29[207]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[115],stage1_31[147],stage1_30[152],stage1_29[208]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[116],stage1_31[148],stage1_30[153],stage1_29[209]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460], stage0_29[461]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[117],stage1_31[149],stage1_30[154],stage1_29[210]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466], stage0_29[467]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[118],stage1_31[150],stage1_30[155],stage1_29[211]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472], stage0_29[473]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[119],stage1_31[151],stage1_30[156],stage1_29[212]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[120],stage1_31[152],stage1_30[157],stage1_29[213]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[121],stage1_31[153],stage1_30[158],stage1_29[214]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490], stage0_29[491]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[122],stage1_31[154],stage1_30[159],stage1_29[215]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496], stage0_29[497]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[123],stage1_31[155],stage1_30[160],stage1_29[216]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502], stage0_29[503]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[124],stage1_31[156],stage1_30[161],stage1_29[217]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508], stage0_29[509]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[125],stage1_31[157],stage1_30[162],stage1_29[218]}
   );
   gpc1415_5 gpc1246 (
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442]},
      {stage0_31[318]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[53],stage1_32[126],stage1_31[158],stage1_30[163]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage0_32[4]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[1],stage1_33[54],stage1_32[127],stage1_31[159]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328]},
      {stage0_32[5]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[2],stage1_33[55],stage1_32[128],stage1_31[160]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[329], stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333]},
      {stage0_32[6]},
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage1_35[2],stage1_34[3],stage1_33[56],stage1_32[129],stage1_31[161]}
   );
   gpc615_5 gpc1250 (
      {stage0_31[334], stage0_31[335], stage0_31[336], stage0_31[337], stage0_31[338]},
      {stage0_32[7]},
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage1_35[3],stage1_34[4],stage1_33[57],stage1_32[130],stage1_31[162]}
   );
   gpc615_5 gpc1251 (
      {stage0_31[339], stage0_31[340], stage0_31[341], stage0_31[342], stage0_31[343]},
      {stage0_32[8]},
      {stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29], stage0_33[30]},
      {stage1_35[4],stage1_34[5],stage1_33[58],stage1_32[131],stage1_31[163]}
   );
   gpc615_5 gpc1252 (
      {stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347], stage0_31[348]},
      {stage0_32[9]},
      {stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35], stage0_33[36]},
      {stage1_35[5],stage1_34[6],stage1_33[59],stage1_32[132],stage1_31[164]}
   );
   gpc615_5 gpc1253 (
      {stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage0_32[10]},
      {stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41], stage0_33[42]},
      {stage1_35[6],stage1_34[7],stage1_33[60],stage1_32[133],stage1_31[165]}
   );
   gpc615_5 gpc1254 (
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358]},
      {stage0_32[11]},
      {stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47], stage0_33[48]},
      {stage1_35[7],stage1_34[8],stage1_33[61],stage1_32[134],stage1_31[166]}
   );
   gpc615_5 gpc1255 (
      {stage0_31[359], stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363]},
      {stage0_32[12]},
      {stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53], stage0_33[54]},
      {stage1_35[8],stage1_34[9],stage1_33[62],stage1_32[135],stage1_31[167]}
   );
   gpc615_5 gpc1256 (
      {stage0_31[364], stage0_31[365], stage0_31[366], stage0_31[367], stage0_31[368]},
      {stage0_32[13]},
      {stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59], stage0_33[60]},
      {stage1_35[9],stage1_34[10],stage1_33[63],stage1_32[136],stage1_31[168]}
   );
   gpc615_5 gpc1257 (
      {stage0_31[369], stage0_31[370], stage0_31[371], stage0_31[372], stage0_31[373]},
      {stage0_32[14]},
      {stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65], stage0_33[66]},
      {stage1_35[10],stage1_34[11],stage1_33[64],stage1_32[137],stage1_31[169]}
   );
   gpc615_5 gpc1258 (
      {stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377], stage0_31[378]},
      {stage0_32[15]},
      {stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71], stage0_33[72]},
      {stage1_35[11],stage1_34[12],stage1_33[65],stage1_32[138],stage1_31[170]}
   );
   gpc615_5 gpc1259 (
      {stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage0_32[16]},
      {stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77], stage0_33[78]},
      {stage1_35[12],stage1_34[13],stage1_33[66],stage1_32[139],stage1_31[171]}
   );
   gpc615_5 gpc1260 (
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388]},
      {stage0_32[17]},
      {stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83], stage0_33[84]},
      {stage1_35[13],stage1_34[14],stage1_33[67],stage1_32[140],stage1_31[172]}
   );
   gpc615_5 gpc1261 (
      {stage0_31[389], stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393]},
      {stage0_32[18]},
      {stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89], stage0_33[90]},
      {stage1_35[14],stage1_34[15],stage1_33[68],stage1_32[141],stage1_31[173]}
   );
   gpc615_5 gpc1262 (
      {stage0_31[394], stage0_31[395], stage0_31[396], stage0_31[397], stage0_31[398]},
      {stage0_32[19]},
      {stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95], stage0_33[96]},
      {stage1_35[15],stage1_34[16],stage1_33[69],stage1_32[142],stage1_31[174]}
   );
   gpc615_5 gpc1263 (
      {stage0_31[399], stage0_31[400], stage0_31[401], stage0_31[402], stage0_31[403]},
      {stage0_32[20]},
      {stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101], stage0_33[102]},
      {stage1_35[16],stage1_34[17],stage1_33[70],stage1_32[143],stage1_31[175]}
   );
   gpc615_5 gpc1264 (
      {stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407], stage0_31[408]},
      {stage0_32[21]},
      {stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107], stage0_33[108]},
      {stage1_35[17],stage1_34[18],stage1_33[71],stage1_32[144],stage1_31[176]}
   );
   gpc615_5 gpc1265 (
      {stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage0_32[22]},
      {stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113], stage0_33[114]},
      {stage1_35[18],stage1_34[19],stage1_33[72],stage1_32[145],stage1_31[177]}
   );
   gpc615_5 gpc1266 (
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418]},
      {stage0_32[23]},
      {stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119], stage0_33[120]},
      {stage1_35[19],stage1_34[20],stage1_33[73],stage1_32[146],stage1_31[178]}
   );
   gpc615_5 gpc1267 (
      {stage0_31[419], stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423]},
      {stage0_32[24]},
      {stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125], stage0_33[126]},
      {stage1_35[20],stage1_34[21],stage1_33[74],stage1_32[147],stage1_31[179]}
   );
   gpc615_5 gpc1268 (
      {stage0_31[424], stage0_31[425], stage0_31[426], stage0_31[427], stage0_31[428]},
      {stage0_32[25]},
      {stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131], stage0_33[132]},
      {stage1_35[21],stage1_34[22],stage1_33[75],stage1_32[148],stage1_31[180]}
   );
   gpc615_5 gpc1269 (
      {stage0_31[429], stage0_31[430], stage0_31[431], stage0_31[432], stage0_31[433]},
      {stage0_32[26]},
      {stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137], stage0_33[138]},
      {stage1_35[22],stage1_34[23],stage1_33[76],stage1_32[149],stage1_31[181]}
   );
   gpc615_5 gpc1270 (
      {stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437], stage0_31[438]},
      {stage0_32[27]},
      {stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143], stage0_33[144]},
      {stage1_35[23],stage1_34[24],stage1_33[77],stage1_32[150],stage1_31[182]}
   );
   gpc615_5 gpc1271 (
      {stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage0_32[28]},
      {stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149], stage0_33[150]},
      {stage1_35[24],stage1_34[25],stage1_33[78],stage1_32[151],stage1_31[183]}
   );
   gpc615_5 gpc1272 (
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448]},
      {stage0_32[29]},
      {stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155], stage0_33[156]},
      {stage1_35[25],stage1_34[26],stage1_33[79],stage1_32[152],stage1_31[184]}
   );
   gpc615_5 gpc1273 (
      {stage0_31[449], stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453]},
      {stage0_32[30]},
      {stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161], stage0_33[162]},
      {stage1_35[26],stage1_34[27],stage1_33[80],stage1_32[153],stage1_31[185]}
   );
   gpc615_5 gpc1274 (
      {stage0_31[454], stage0_31[455], stage0_31[456], stage0_31[457], stage0_31[458]},
      {stage0_32[31]},
      {stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167], stage0_33[168]},
      {stage1_35[27],stage1_34[28],stage1_33[81],stage1_32[154],stage1_31[186]}
   );
   gpc615_5 gpc1275 (
      {stage0_31[459], stage0_31[460], stage0_31[461], stage0_31[462], stage0_31[463]},
      {stage0_32[32]},
      {stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173], stage0_33[174]},
      {stage1_35[28],stage1_34[29],stage1_33[82],stage1_32[155],stage1_31[187]}
   );
   gpc615_5 gpc1276 (
      {stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467], stage0_31[468]},
      {stage0_32[33]},
      {stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179], stage0_33[180]},
      {stage1_35[29],stage1_34[30],stage1_33[83],stage1_32[156],stage1_31[188]}
   );
   gpc615_5 gpc1277 (
      {stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage0_32[34]},
      {stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185], stage0_33[186]},
      {stage1_35[30],stage1_34[31],stage1_33[84],stage1_32[157],stage1_31[189]}
   );
   gpc615_5 gpc1278 (
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478]},
      {stage0_32[35]},
      {stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191], stage0_33[192]},
      {stage1_35[31],stage1_34[32],stage1_33[85],stage1_32[158],stage1_31[190]}
   );
   gpc615_5 gpc1279 (
      {stage0_31[479], stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483]},
      {stage0_32[36]},
      {stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197], stage0_33[198]},
      {stage1_35[32],stage1_34[33],stage1_33[86],stage1_32[159],stage1_31[191]}
   );
   gpc615_5 gpc1280 (
      {stage0_31[484], stage0_31[485], stage0_31[486], stage0_31[487], stage0_31[488]},
      {stage0_32[37]},
      {stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203], stage0_33[204]},
      {stage1_35[33],stage1_34[34],stage1_33[87],stage1_32[160],stage1_31[192]}
   );
   gpc615_5 gpc1281 (
      {stage0_31[489], stage0_31[490], stage0_31[491], stage0_31[492], stage0_31[493]},
      {stage0_32[38]},
      {stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209], stage0_33[210]},
      {stage1_35[34],stage1_34[35],stage1_33[88],stage1_32[161],stage1_31[193]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[35],stage1_34[36],stage1_33[89],stage1_32[162]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[36],stage1_34[37],stage1_33[90],stage1_32[163]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[37],stage1_34[38],stage1_33[91],stage1_32[164]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[38],stage1_34[39],stage1_33[92],stage1_32[165]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[63], stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[39],stage1_34[40],stage1_33[93],stage1_32[166]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73], stage0_32[74]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[40],stage1_34[41],stage1_33[94],stage1_32[167]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78], stage0_32[79], stage0_32[80]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[41],stage1_34[42],stage1_33[95],stage1_32[168]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[81], stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[42],stage1_34[43],stage1_33[96],stage1_32[169]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[87], stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[43],stage1_34[44],stage1_33[97],stage1_32[170]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[93], stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[44],stage1_34[45],stage1_33[98],stage1_32[171]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103], stage0_32[104]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[45],stage1_34[46],stage1_33[99],stage1_32[172]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108], stage0_32[109], stage0_32[110]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[46],stage1_34[47],stage1_33[100],stage1_32[173]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[111], stage0_32[112], stage0_32[113], stage0_32[114], stage0_32[115], stage0_32[116]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[47],stage1_34[48],stage1_33[101],stage1_32[174]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[117], stage0_32[118], stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[48],stage1_34[49],stage1_33[102],stage1_32[175]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[123], stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[49],stage1_34[50],stage1_33[103],stage1_32[176]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[129], stage0_32[130], stage0_32[131], stage0_32[132], stage0_32[133], stage0_32[134]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[50],stage1_34[51],stage1_33[104],stage1_32[177]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[135], stage0_32[136], stage0_32[137], stage0_32[138], stage0_32[139], stage0_32[140]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[51],stage1_34[52],stage1_33[105],stage1_32[178]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[141], stage0_32[142], stage0_32[143], stage0_32[144], stage0_32[145], stage0_32[146]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[52],stage1_34[53],stage1_33[106],stage1_32[179]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[147], stage0_32[148], stage0_32[149], stage0_32[150], stage0_32[151], stage0_32[152]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[53],stage1_34[54],stage1_33[107],stage1_32[180]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[153], stage0_32[154], stage0_32[155], stage0_32[156], stage0_32[157], stage0_32[158]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[54],stage1_34[55],stage1_33[108],stage1_32[181]}
   );
   gpc606_5 gpc1302 (
      {stage0_32[159], stage0_32[160], stage0_32[161], stage0_32[162], stage0_32[163], stage0_32[164]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[55],stage1_34[56],stage1_33[109],stage1_32[182]}
   );
   gpc606_5 gpc1303 (
      {stage0_32[165], stage0_32[166], stage0_32[167], stage0_32[168], stage0_32[169], stage0_32[170]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[56],stage1_34[57],stage1_33[110],stage1_32[183]}
   );
   gpc606_5 gpc1304 (
      {stage0_32[171], stage0_32[172], stage0_32[173], stage0_32[174], stage0_32[175], stage0_32[176]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[57],stage1_34[58],stage1_33[111],stage1_32[184]}
   );
   gpc606_5 gpc1305 (
      {stage0_32[177], stage0_32[178], stage0_32[179], stage0_32[180], stage0_32[181], stage0_32[182]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[58],stage1_34[59],stage1_33[112],stage1_32[185]}
   );
   gpc606_5 gpc1306 (
      {stage0_32[183], stage0_32[184], stage0_32[185], stage0_32[186], stage0_32[187], stage0_32[188]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[59],stage1_34[60],stage1_33[113],stage1_32[186]}
   );
   gpc606_5 gpc1307 (
      {stage0_32[189], stage0_32[190], stage0_32[191], stage0_32[192], stage0_32[193], stage0_32[194]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[60],stage1_34[61],stage1_33[114],stage1_32[187]}
   );
   gpc606_5 gpc1308 (
      {stage0_32[195], stage0_32[196], stage0_32[197], stage0_32[198], stage0_32[199], stage0_32[200]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[61],stage1_34[62],stage1_33[115],stage1_32[188]}
   );
   gpc606_5 gpc1309 (
      {stage0_32[201], stage0_32[202], stage0_32[203], stage0_32[204], stage0_32[205], stage0_32[206]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[62],stage1_34[63],stage1_33[116],stage1_32[189]}
   );
   gpc606_5 gpc1310 (
      {stage0_32[207], stage0_32[208], stage0_32[209], stage0_32[210], stage0_32[211], stage0_32[212]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[63],stage1_34[64],stage1_33[117],stage1_32[190]}
   );
   gpc606_5 gpc1311 (
      {stage0_32[213], stage0_32[214], stage0_32[215], stage0_32[216], stage0_32[217], stage0_32[218]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[64],stage1_34[65],stage1_33[118],stage1_32[191]}
   );
   gpc606_5 gpc1312 (
      {stage0_32[219], stage0_32[220], stage0_32[221], stage0_32[222], stage0_32[223], stage0_32[224]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[65],stage1_34[66],stage1_33[119],stage1_32[192]}
   );
   gpc606_5 gpc1313 (
      {stage0_32[225], stage0_32[226], stage0_32[227], stage0_32[228], stage0_32[229], stage0_32[230]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[66],stage1_34[67],stage1_33[120],stage1_32[193]}
   );
   gpc606_5 gpc1314 (
      {stage0_32[231], stage0_32[232], stage0_32[233], stage0_32[234], stage0_32[235], stage0_32[236]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[67],stage1_34[68],stage1_33[121],stage1_32[194]}
   );
   gpc606_5 gpc1315 (
      {stage0_32[237], stage0_32[238], stage0_32[239], stage0_32[240], stage0_32[241], stage0_32[242]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[68],stage1_34[69],stage1_33[122],stage1_32[195]}
   );
   gpc606_5 gpc1316 (
      {stage0_32[243], stage0_32[244], stage0_32[245], stage0_32[246], stage0_32[247], stage0_32[248]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[69],stage1_34[70],stage1_33[123],stage1_32[196]}
   );
   gpc606_5 gpc1317 (
      {stage0_32[249], stage0_32[250], stage0_32[251], stage0_32[252], stage0_32[253], stage0_32[254]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[70],stage1_34[71],stage1_33[124],stage1_32[197]}
   );
   gpc606_5 gpc1318 (
      {stage0_32[255], stage0_32[256], stage0_32[257], stage0_32[258], stage0_32[259], stage0_32[260]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[71],stage1_34[72],stage1_33[125],stage1_32[198]}
   );
   gpc606_5 gpc1319 (
      {stage0_32[261], stage0_32[262], stage0_32[263], stage0_32[264], stage0_32[265], stage0_32[266]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[72],stage1_34[73],stage1_33[126],stage1_32[199]}
   );
   gpc606_5 gpc1320 (
      {stage0_32[267], stage0_32[268], stage0_32[269], stage0_32[270], stage0_32[271], stage0_32[272]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[73],stage1_34[74],stage1_33[127],stage1_32[200]}
   );
   gpc606_5 gpc1321 (
      {stage0_32[273], stage0_32[274], stage0_32[275], stage0_32[276], stage0_32[277], stage0_32[278]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[74],stage1_34[75],stage1_33[128],stage1_32[201]}
   );
   gpc606_5 gpc1322 (
      {stage0_32[279], stage0_32[280], stage0_32[281], stage0_32[282], stage0_32[283], stage0_32[284]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[75],stage1_34[76],stage1_33[129],stage1_32[202]}
   );
   gpc606_5 gpc1323 (
      {stage0_32[285], stage0_32[286], stage0_32[287], stage0_32[288], stage0_32[289], stage0_32[290]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[76],stage1_34[77],stage1_33[130],stage1_32[203]}
   );
   gpc606_5 gpc1324 (
      {stage0_32[291], stage0_32[292], stage0_32[293], stage0_32[294], stage0_32[295], stage0_32[296]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[77],stage1_34[78],stage1_33[131],stage1_32[204]}
   );
   gpc606_5 gpc1325 (
      {stage0_32[297], stage0_32[298], stage0_32[299], stage0_32[300], stage0_32[301], stage0_32[302]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[78],stage1_34[79],stage1_33[132],stage1_32[205]}
   );
   gpc615_5 gpc1326 (
      {stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage0_34[264]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[44],stage1_35[79],stage1_34[80],stage1_33[133]}
   );
   gpc615_5 gpc1327 (
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220]},
      {stage0_34[265]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[45],stage1_35[80],stage1_34[81],stage1_33[134]}
   );
   gpc615_5 gpc1328 (
      {stage0_33[221], stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225]},
      {stage0_34[266]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[46],stage1_35[81],stage1_34[82],stage1_33[135]}
   );
   gpc615_5 gpc1329 (
      {stage0_33[226], stage0_33[227], stage0_33[228], stage0_33[229], stage0_33[230]},
      {stage0_34[267]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[47],stage1_35[82],stage1_34[83],stage1_33[136]}
   );
   gpc615_5 gpc1330 (
      {stage0_33[231], stage0_33[232], stage0_33[233], stage0_33[234], stage0_33[235]},
      {stage0_34[268]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[48],stage1_35[83],stage1_34[84],stage1_33[137]}
   );
   gpc615_5 gpc1331 (
      {stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239], stage0_33[240]},
      {stage0_34[269]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[49],stage1_35[84],stage1_34[85],stage1_33[138]}
   );
   gpc615_5 gpc1332 (
      {stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage0_34[270]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[50],stage1_35[85],stage1_34[86],stage1_33[139]}
   );
   gpc615_5 gpc1333 (
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250]},
      {stage0_34[271]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[51],stage1_35[86],stage1_34[87],stage1_33[140]}
   );
   gpc615_5 gpc1334 (
      {stage0_33[251], stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255]},
      {stage0_34[272]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[52],stage1_35[87],stage1_34[88],stage1_33[141]}
   );
   gpc615_5 gpc1335 (
      {stage0_33[256], stage0_33[257], stage0_33[258], stage0_33[259], stage0_33[260]},
      {stage0_34[273]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[53],stage1_35[88],stage1_34[89],stage1_33[142]}
   );
   gpc615_5 gpc1336 (
      {stage0_33[261], stage0_33[262], stage0_33[263], stage0_33[264], stage0_33[265]},
      {stage0_34[274]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[54],stage1_35[89],stage1_34[90],stage1_33[143]}
   );
   gpc615_5 gpc1337 (
      {stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269], stage0_33[270]},
      {stage0_34[275]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[55],stage1_35[90],stage1_34[91],stage1_33[144]}
   );
   gpc615_5 gpc1338 (
      {stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage0_34[276]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[56],stage1_35[91],stage1_34[92],stage1_33[145]}
   );
   gpc615_5 gpc1339 (
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280]},
      {stage0_34[277]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[57],stage1_35[92],stage1_34[93],stage1_33[146]}
   );
   gpc615_5 gpc1340 (
      {stage0_33[281], stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285]},
      {stage0_34[278]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[58],stage1_35[93],stage1_34[94],stage1_33[147]}
   );
   gpc615_5 gpc1341 (
      {stage0_33[286], stage0_33[287], stage0_33[288], stage0_33[289], stage0_33[290]},
      {stage0_34[279]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[59],stage1_35[94],stage1_34[95],stage1_33[148]}
   );
   gpc615_5 gpc1342 (
      {stage0_33[291], stage0_33[292], stage0_33[293], stage0_33[294], stage0_33[295]},
      {stage0_34[280]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[60],stage1_35[95],stage1_34[96],stage1_33[149]}
   );
   gpc615_5 gpc1343 (
      {stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299], stage0_33[300]},
      {stage0_34[281]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[61],stage1_35[96],stage1_34[97],stage1_33[150]}
   );
   gpc615_5 gpc1344 (
      {stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage0_34[282]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage1_37[18],stage1_36[62],stage1_35[97],stage1_34[98],stage1_33[151]}
   );
   gpc615_5 gpc1345 (
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310]},
      {stage0_34[283]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage1_37[19],stage1_36[63],stage1_35[98],stage1_34[99],stage1_33[152]}
   );
   gpc615_5 gpc1346 (
      {stage0_33[311], stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315]},
      {stage0_34[284]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage1_37[20],stage1_36[64],stage1_35[99],stage1_34[100],stage1_33[153]}
   );
   gpc615_5 gpc1347 (
      {stage0_33[316], stage0_33[317], stage0_33[318], stage0_33[319], stage0_33[320]},
      {stage0_34[285]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage1_37[21],stage1_36[65],stage1_35[100],stage1_34[101],stage1_33[154]}
   );
   gpc615_5 gpc1348 (
      {stage0_33[321], stage0_33[322], stage0_33[323], stage0_33[324], stage0_33[325]},
      {stage0_34[286]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage1_37[22],stage1_36[66],stage1_35[101],stage1_34[102],stage1_33[155]}
   );
   gpc615_5 gpc1349 (
      {stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329], stage0_33[330]},
      {stage0_34[287]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage1_37[23],stage1_36[67],stage1_35[102],stage1_34[103],stage1_33[156]}
   );
   gpc615_5 gpc1350 (
      {stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_34[288]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage1_37[24],stage1_36[68],stage1_35[103],stage1_34[104],stage1_33[157]}
   );
   gpc615_5 gpc1351 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340]},
      {stage0_34[289]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage1_37[25],stage1_36[69],stage1_35[104],stage1_34[105],stage1_33[158]}
   );
   gpc615_5 gpc1352 (
      {stage0_33[341], stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345]},
      {stage0_34[290]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage1_37[26],stage1_36[70],stage1_35[105],stage1_34[106],stage1_33[159]}
   );
   gpc615_5 gpc1353 (
      {stage0_33[346], stage0_33[347], stage0_33[348], stage0_33[349], stage0_33[350]},
      {stage0_34[291]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage1_37[27],stage1_36[71],stage1_35[106],stage1_34[107],stage1_33[160]}
   );
   gpc615_5 gpc1354 (
      {stage0_33[351], stage0_33[352], stage0_33[353], stage0_33[354], stage0_33[355]},
      {stage0_34[292]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage1_37[28],stage1_36[72],stage1_35[107],stage1_34[108],stage1_33[161]}
   );
   gpc615_5 gpc1355 (
      {stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359], stage0_33[360]},
      {stage0_34[293]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage1_37[29],stage1_36[73],stage1_35[108],stage1_34[109],stage1_33[162]}
   );
   gpc615_5 gpc1356 (
      {stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_34[294]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage1_37[30],stage1_36[74],stage1_35[109],stage1_34[110],stage1_33[163]}
   );
   gpc615_5 gpc1357 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370]},
      {stage0_34[295]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage1_37[31],stage1_36[75],stage1_35[110],stage1_34[111],stage1_33[164]}
   );
   gpc615_5 gpc1358 (
      {stage0_33[371], stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375]},
      {stage0_34[296]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage1_37[32],stage1_36[76],stage1_35[111],stage1_34[112],stage1_33[165]}
   );
   gpc615_5 gpc1359 (
      {stage0_33[376], stage0_33[377], stage0_33[378], stage0_33[379], stage0_33[380]},
      {stage0_34[297]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage1_37[33],stage1_36[77],stage1_35[112],stage1_34[113],stage1_33[166]}
   );
   gpc615_5 gpc1360 (
      {stage0_33[381], stage0_33[382], stage0_33[383], stage0_33[384], stage0_33[385]},
      {stage0_34[298]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage1_37[34],stage1_36[78],stage1_35[113],stage1_34[114],stage1_33[167]}
   );
   gpc615_5 gpc1361 (
      {stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389], stage0_33[390]},
      {stage0_34[299]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage1_37[35],stage1_36[79],stage1_35[114],stage1_34[115],stage1_33[168]}
   );
   gpc615_5 gpc1362 (
      {stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_34[300]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage1_37[36],stage1_36[80],stage1_35[115],stage1_34[116],stage1_33[169]}
   );
   gpc615_5 gpc1363 (
      {stage0_33[396], stage0_33[397], stage0_33[398], stage0_33[399], stage0_33[400]},
      {stage0_34[301]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage1_37[37],stage1_36[81],stage1_35[116],stage1_34[117],stage1_33[170]}
   );
   gpc615_5 gpc1364 (
      {stage0_33[401], stage0_33[402], stage0_33[403], stage0_33[404], stage0_33[405]},
      {stage0_34[302]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage1_37[38],stage1_36[82],stage1_35[117],stage1_34[118],stage1_33[171]}
   );
   gpc615_5 gpc1365 (
      {stage0_33[406], stage0_33[407], stage0_33[408], stage0_33[409], stage0_33[410]},
      {stage0_34[303]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage1_37[39],stage1_36[83],stage1_35[118],stage1_34[119],stage1_33[172]}
   );
   gpc615_5 gpc1366 (
      {stage0_33[411], stage0_33[412], stage0_33[413], stage0_33[414], stage0_33[415]},
      {stage0_34[304]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage1_37[40],stage1_36[84],stage1_35[119],stage1_34[120],stage1_33[173]}
   );
   gpc615_5 gpc1367 (
      {stage0_33[416], stage0_33[417], stage0_33[418], stage0_33[419], stage0_33[420]},
      {stage0_34[305]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage1_37[41],stage1_36[85],stage1_35[120],stage1_34[121],stage1_33[174]}
   );
   gpc615_5 gpc1368 (
      {stage0_33[421], stage0_33[422], stage0_33[423], stage0_33[424], stage0_33[425]},
      {stage0_34[306]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage1_37[42],stage1_36[86],stage1_35[121],stage1_34[122],stage1_33[175]}
   );
   gpc615_5 gpc1369 (
      {stage0_33[426], stage0_33[427], stage0_33[428], stage0_33[429], stage0_33[430]},
      {stage0_34[307]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage1_37[43],stage1_36[87],stage1_35[122],stage1_34[123],stage1_33[176]}
   );
   gpc615_5 gpc1370 (
      {stage0_33[431], stage0_33[432], stage0_33[433], stage0_33[434], stage0_33[435]},
      {stage0_34[308]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage1_37[44],stage1_36[88],stage1_35[123],stage1_34[124],stage1_33[177]}
   );
   gpc615_5 gpc1371 (
      {stage0_33[436], stage0_33[437], stage0_33[438], stage0_33[439], stage0_33[440]},
      {stage0_34[309]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage1_37[45],stage1_36[89],stage1_35[124],stage1_34[125],stage1_33[178]}
   );
   gpc615_5 gpc1372 (
      {stage0_33[441], stage0_33[442], stage0_33[443], stage0_33[444], stage0_33[445]},
      {stage0_34[310]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage1_37[46],stage1_36[90],stage1_35[125],stage1_34[126],stage1_33[179]}
   );
   gpc615_5 gpc1373 (
      {stage0_33[446], stage0_33[447], stage0_33[448], stage0_33[449], stage0_33[450]},
      {stage0_34[311]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage1_37[47],stage1_36[91],stage1_35[126],stage1_34[127],stage1_33[180]}
   );
   gpc615_5 gpc1374 (
      {stage0_33[451], stage0_33[452], stage0_33[453], stage0_33[454], stage0_33[455]},
      {stage0_34[312]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage1_37[48],stage1_36[92],stage1_35[127],stage1_34[128],stage1_33[181]}
   );
   gpc615_5 gpc1375 (
      {stage0_33[456], stage0_33[457], stage0_33[458], stage0_33[459], stage0_33[460]},
      {stage0_34[313]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage1_37[49],stage1_36[93],stage1_35[128],stage1_34[129],stage1_33[182]}
   );
   gpc615_5 gpc1376 (
      {stage0_33[461], stage0_33[462], stage0_33[463], stage0_33[464], stage0_33[465]},
      {stage0_34[314]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage1_37[50],stage1_36[94],stage1_35[129],stage1_34[130],stage1_33[183]}
   );
   gpc615_5 gpc1377 (
      {stage0_33[466], stage0_33[467], stage0_33[468], stage0_33[469], stage0_33[470]},
      {stage0_34[315]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage1_37[51],stage1_36[95],stage1_35[130],stage1_34[131],stage1_33[184]}
   );
   gpc615_5 gpc1378 (
      {stage0_33[471], stage0_33[472], stage0_33[473], stage0_33[474], stage0_33[475]},
      {stage0_34[316]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage1_37[52],stage1_36[96],stage1_35[131],stage1_34[132],stage1_33[185]}
   );
   gpc615_5 gpc1379 (
      {stage0_33[476], stage0_33[477], stage0_33[478], stage0_33[479], stage0_33[480]},
      {stage0_34[317]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage1_37[53],stage1_36[97],stage1_35[132],stage1_34[133],stage1_33[186]}
   );
   gpc615_5 gpc1380 (
      {stage0_33[481], stage0_33[482], stage0_33[483], stage0_33[484], stage0_33[485]},
      {stage0_34[318]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage1_37[54],stage1_36[98],stage1_35[133],stage1_34[134],stage1_33[187]}
   );
   gpc615_5 gpc1381 (
      {stage0_33[486], stage0_33[487], stage0_33[488], stage0_33[489], stage0_33[490]},
      {stage0_34[319]},
      {stage0_35[330], stage0_35[331], stage0_35[332], stage0_35[333], stage0_35[334], stage0_35[335]},
      {stage1_37[55],stage1_36[99],stage1_35[134],stage1_34[135],stage1_33[188]}
   );
   gpc1163_5 gpc1382 (
      {stage0_34[320], stage0_34[321], stage0_34[322]},
      {stage0_35[336], stage0_35[337], stage0_35[338], stage0_35[339], stage0_35[340], stage0_35[341]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[56],stage1_36[100],stage1_35[135],stage1_34[136]}
   );
   gpc1163_5 gpc1383 (
      {stage0_34[323], stage0_34[324], stage0_34[325]},
      {stage0_35[342], stage0_35[343], stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[57],stage1_36[101],stage1_35[136],stage1_34[137]}
   );
   gpc615_5 gpc1384 (
      {stage0_34[326], stage0_34[327], stage0_34[328], stage0_34[329], stage0_34[330]},
      {stage0_35[348]},
      {stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5], stage0_36[6], stage0_36[7]},
      {stage1_38[2],stage1_37[58],stage1_36[102],stage1_35[137],stage1_34[138]}
   );
   gpc615_5 gpc1385 (
      {stage0_34[331], stage0_34[332], stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[349]},
      {stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13]},
      {stage1_38[3],stage1_37[59],stage1_36[103],stage1_35[138],stage1_34[139]}
   );
   gpc615_5 gpc1386 (
      {stage0_34[336], stage0_34[337], stage0_34[338], stage0_34[339], stage0_34[340]},
      {stage0_35[350]},
      {stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19]},
      {stage1_38[4],stage1_37[60],stage1_36[104],stage1_35[139],stage1_34[140]}
   );
   gpc615_5 gpc1387 (
      {stage0_34[341], stage0_34[342], stage0_34[343], stage0_34[344], stage0_34[345]},
      {stage0_35[351]},
      {stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25]},
      {stage1_38[5],stage1_37[61],stage1_36[105],stage1_35[140],stage1_34[141]}
   );
   gpc615_5 gpc1388 (
      {stage0_34[346], stage0_34[347], stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[352]},
      {stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31]},
      {stage1_38[6],stage1_37[62],stage1_36[106],stage1_35[141],stage1_34[142]}
   );
   gpc615_5 gpc1389 (
      {stage0_34[351], stage0_34[352], stage0_34[353], stage0_34[354], stage0_34[355]},
      {stage0_35[353]},
      {stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37]},
      {stage1_38[7],stage1_37[63],stage1_36[107],stage1_35[142],stage1_34[143]}
   );
   gpc615_5 gpc1390 (
      {stage0_34[356], stage0_34[357], stage0_34[358], stage0_34[359], stage0_34[360]},
      {stage0_35[354]},
      {stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43]},
      {stage1_38[8],stage1_37[64],stage1_36[108],stage1_35[143],stage1_34[144]}
   );
   gpc615_5 gpc1391 (
      {stage0_34[361], stage0_34[362], stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[355]},
      {stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48], stage0_36[49]},
      {stage1_38[9],stage1_37[65],stage1_36[109],stage1_35[144],stage1_34[145]}
   );
   gpc615_5 gpc1392 (
      {stage0_34[366], stage0_34[367], stage0_34[368], stage0_34[369], stage0_34[370]},
      {stage0_35[356]},
      {stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54], stage0_36[55]},
      {stage1_38[10],stage1_37[66],stage1_36[110],stage1_35[145],stage1_34[146]}
   );
   gpc615_5 gpc1393 (
      {stage0_34[371], stage0_34[372], stage0_34[373], stage0_34[374], stage0_34[375]},
      {stage0_35[357]},
      {stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60], stage0_36[61]},
      {stage1_38[11],stage1_37[67],stage1_36[111],stage1_35[146],stage1_34[147]}
   );
   gpc615_5 gpc1394 (
      {stage0_34[376], stage0_34[377], stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[358]},
      {stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66], stage0_36[67]},
      {stage1_38[12],stage1_37[68],stage1_36[112],stage1_35[147],stage1_34[148]}
   );
   gpc615_5 gpc1395 (
      {stage0_34[381], stage0_34[382], stage0_34[383], stage0_34[384], stage0_34[385]},
      {stage0_35[359]},
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage1_38[13],stage1_37[69],stage1_36[113],stage1_35[148],stage1_34[149]}
   );
   gpc615_5 gpc1396 (
      {stage0_34[386], stage0_34[387], stage0_34[388], stage0_34[389], stage0_34[390]},
      {stage0_35[360]},
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage1_38[14],stage1_37[70],stage1_36[114],stage1_35[149],stage1_34[150]}
   );
   gpc615_5 gpc1397 (
      {stage0_34[391], stage0_34[392], stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[361]},
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage1_38[15],stage1_37[71],stage1_36[115],stage1_35[150],stage1_34[151]}
   );
   gpc606_5 gpc1398 (
      {stage0_35[362], stage0_35[363], stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367]},
      {stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5], stage0_37[6], stage0_37[7]},
      {stage1_39[0],stage1_38[16],stage1_37[72],stage1_36[116],stage1_35[151]}
   );
   gpc606_5 gpc1399 (
      {stage0_35[368], stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12], stage0_37[13]},
      {stage1_39[1],stage1_38[17],stage1_37[73],stage1_36[117],stage1_35[152]}
   );
   gpc606_5 gpc1400 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378], stage0_35[379]},
      {stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17], stage0_37[18], stage0_37[19]},
      {stage1_39[2],stage1_38[18],stage1_37[74],stage1_36[118],stage1_35[153]}
   );
   gpc606_5 gpc1401 (
      {stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383], stage0_35[384], stage0_35[385]},
      {stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23], stage0_37[24], stage0_37[25]},
      {stage1_39[3],stage1_38[19],stage1_37[75],stage1_36[119],stage1_35[154]}
   );
   gpc606_5 gpc1402 (
      {stage0_35[386], stage0_35[387], stage0_35[388], stage0_35[389], stage0_35[390], stage0_35[391]},
      {stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29], stage0_37[30], stage0_37[31]},
      {stage1_39[4],stage1_38[20],stage1_37[76],stage1_36[120],stage1_35[155]}
   );
   gpc606_5 gpc1403 (
      {stage0_35[392], stage0_35[393], stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397]},
      {stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35], stage0_37[36], stage0_37[37]},
      {stage1_39[5],stage1_38[21],stage1_37[77],stage1_36[121],stage1_35[156]}
   );
   gpc606_5 gpc1404 (
      {stage0_35[398], stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41], stage0_37[42], stage0_37[43]},
      {stage1_39[6],stage1_38[22],stage1_37[78],stage1_36[122],stage1_35[157]}
   );
   gpc606_5 gpc1405 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408], stage0_35[409]},
      {stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48], stage0_37[49]},
      {stage1_39[7],stage1_38[23],stage1_37[79],stage1_36[123],stage1_35[158]}
   );
   gpc606_5 gpc1406 (
      {stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413], stage0_35[414], stage0_35[415]},
      {stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54], stage0_37[55]},
      {stage1_39[8],stage1_38[24],stage1_37[80],stage1_36[124],stage1_35[159]}
   );
   gpc606_5 gpc1407 (
      {stage0_35[416], stage0_35[417], stage0_35[418], stage0_35[419], stage0_35[420], stage0_35[421]},
      {stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60], stage0_37[61]},
      {stage1_39[9],stage1_38[25],stage1_37[81],stage1_36[125],stage1_35[160]}
   );
   gpc606_5 gpc1408 (
      {stage0_35[422], stage0_35[423], stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427]},
      {stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66], stage0_37[67]},
      {stage1_39[10],stage1_38[26],stage1_37[82],stage1_36[126],stage1_35[161]}
   );
   gpc606_5 gpc1409 (
      {stage0_35[428], stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72], stage0_37[73]},
      {stage1_39[11],stage1_38[27],stage1_37[83],stage1_36[127],stage1_35[162]}
   );
   gpc606_5 gpc1410 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438], stage0_35[439]},
      {stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78], stage0_37[79]},
      {stage1_39[12],stage1_38[28],stage1_37[84],stage1_36[128],stage1_35[163]}
   );
   gpc606_5 gpc1411 (
      {stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443], stage0_35[444], stage0_35[445]},
      {stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84], stage0_37[85]},
      {stage1_39[13],stage1_38[29],stage1_37[85],stage1_36[129],stage1_35[164]}
   );
   gpc606_5 gpc1412 (
      {stage0_35[446], stage0_35[447], stage0_35[448], stage0_35[449], stage0_35[450], stage0_35[451]},
      {stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90], stage0_37[91]},
      {stage1_39[14],stage1_38[30],stage1_37[86],stage1_36[130],stage1_35[165]}
   );
   gpc606_5 gpc1413 (
      {stage0_35[452], stage0_35[453], stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457]},
      {stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96], stage0_37[97]},
      {stage1_39[15],stage1_38[31],stage1_37[87],stage1_36[131],stage1_35[166]}
   );
   gpc606_5 gpc1414 (
      {stage0_35[458], stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102], stage0_37[103]},
      {stage1_39[16],stage1_38[32],stage1_37[88],stage1_36[132],stage1_35[167]}
   );
   gpc606_5 gpc1415 (
      {stage0_35[464], stage0_35[465], stage0_35[466], stage0_35[467], stage0_35[468], stage0_35[469]},
      {stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108], stage0_37[109]},
      {stage1_39[17],stage1_38[33],stage1_37[89],stage1_36[133],stage1_35[168]}
   );
   gpc615_5 gpc1416 (
      {stage0_35[470], stage0_35[471], stage0_35[472], stage0_35[473], stage0_35[474]},
      {stage0_36[86]},
      {stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114], stage0_37[115]},
      {stage1_39[18],stage1_38[34],stage1_37[90],stage1_36[134],stage1_35[169]}
   );
   gpc615_5 gpc1417 (
      {stage0_35[475], stage0_35[476], stage0_35[477], stage0_35[478], stage0_35[479]},
      {stage0_36[87]},
      {stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120], stage0_37[121]},
      {stage1_39[19],stage1_38[35],stage1_37[91],stage1_36[135],stage1_35[170]}
   );
   gpc615_5 gpc1418 (
      {stage0_35[480], stage0_35[481], stage0_35[482], stage0_35[483], stage0_35[484]},
      {stage0_36[88]},
      {stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126], stage0_37[127]},
      {stage1_39[20],stage1_38[36],stage1_37[92],stage1_36[136],stage1_35[171]}
   );
   gpc615_5 gpc1419 (
      {stage0_35[485], stage0_35[486], stage0_35[487], stage0_35[488], stage0_35[489]},
      {stage0_36[89]},
      {stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132], stage0_37[133]},
      {stage1_39[21],stage1_38[37],stage1_37[93],stage1_36[137],stage1_35[172]}
   );
   gpc615_5 gpc1420 (
      {stage0_35[490], stage0_35[491], stage0_35[492], stage0_35[493], stage0_35[494]},
      {stage0_36[90]},
      {stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138], stage0_37[139]},
      {stage1_39[22],stage1_38[38],stage1_37[94],stage1_36[138],stage1_35[173]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[23],stage1_38[39],stage1_37[95],stage1_36[139]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[97], stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[24],stage1_38[40],stage1_37[96],stage1_36[140]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[25],stage1_38[41],stage1_37[97],stage1_36[141]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[109], stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[26],stage1_38[42],stage1_37[98],stage1_36[142]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[115], stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[27],stage1_38[43],stage1_37[99],stage1_36[143]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[121], stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[28],stage1_38[44],stage1_37[100],stage1_36[144]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[127], stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[29],stage1_38[45],stage1_37[101],stage1_36[145]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[133], stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[30],stage1_38[46],stage1_37[102],stage1_36[146]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[139], stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[31],stage1_38[47],stage1_37[103],stage1_36[147]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[145], stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[32],stage1_38[48],stage1_37[104],stage1_36[148]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[151], stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[33],stage1_38[49],stage1_37[105],stage1_36[149]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[157], stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[34],stage1_38[50],stage1_37[106],stage1_36[150]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[163], stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[35],stage1_38[51],stage1_37[107],stage1_36[151]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[169], stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[36],stage1_38[52],stage1_37[108],stage1_36[152]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[175], stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[37],stage1_38[53],stage1_37[109],stage1_36[153]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[181], stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[38],stage1_38[54],stage1_37[110],stage1_36[154]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[187], stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[39],stage1_38[55],stage1_37[111],stage1_36[155]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[193], stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[40],stage1_38[56],stage1_37[112],stage1_36[156]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[199], stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[41],stage1_38[57],stage1_37[113],stage1_36[157]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[205], stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[42],stage1_38[58],stage1_37[114],stage1_36[158]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[211], stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[43],stage1_38[59],stage1_37[115],stage1_36[159]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[217], stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[44],stage1_38[60],stage1_37[116],stage1_36[160]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[223], stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[45],stage1_38[61],stage1_37[117],stage1_36[161]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[229], stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[46],stage1_38[62],stage1_37[118],stage1_36[162]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[235], stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[47],stage1_38[63],stage1_37[119],stage1_36[163]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[241], stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[48],stage1_38[64],stage1_37[120],stage1_36[164]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[247], stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[49],stage1_38[65],stage1_37[121],stage1_36[165]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[253], stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[50],stage1_38[66],stage1_37[122],stage1_36[166]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[259], stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[51],stage1_38[67],stage1_37[123],stage1_36[167]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[265], stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[52],stage1_38[68],stage1_37[124],stage1_36[168]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[271], stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[53],stage1_38[69],stage1_37[125],stage1_36[169]}
   );
   gpc606_5 gpc1452 (
      {stage0_36[277], stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[54],stage1_38[70],stage1_37[126],stage1_36[170]}
   );
   gpc606_5 gpc1453 (
      {stage0_36[283], stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[55],stage1_38[71],stage1_37[127],stage1_36[171]}
   );
   gpc606_5 gpc1454 (
      {stage0_36[289], stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[56],stage1_38[72],stage1_37[128],stage1_36[172]}
   );
   gpc606_5 gpc1455 (
      {stage0_36[295], stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[57],stage1_38[73],stage1_37[129],stage1_36[173]}
   );
   gpc606_5 gpc1456 (
      {stage0_36[301], stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[58],stage1_38[74],stage1_37[130],stage1_36[174]}
   );
   gpc606_5 gpc1457 (
      {stage0_36[307], stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[59],stage1_38[75],stage1_37[131],stage1_36[175]}
   );
   gpc606_5 gpc1458 (
      {stage0_36[313], stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[60],stage1_38[76],stage1_37[132],stage1_36[176]}
   );
   gpc606_5 gpc1459 (
      {stage0_36[319], stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[61],stage1_38[77],stage1_37[133],stage1_36[177]}
   );
   gpc606_5 gpc1460 (
      {stage0_36[325], stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[62],stage1_38[78],stage1_37[134],stage1_36[178]}
   );
   gpc606_5 gpc1461 (
      {stage0_36[331], stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[63],stage1_38[79],stage1_37[135],stage1_36[179]}
   );
   gpc615_5 gpc1462 (
      {stage0_36[337], stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341]},
      {stage0_37[140]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[64],stage1_38[80],stage1_37[136],stage1_36[180]}
   );
   gpc615_5 gpc1463 (
      {stage0_36[342], stage0_36[343], stage0_36[344], stage0_36[345], stage0_36[346]},
      {stage0_37[141]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[65],stage1_38[81],stage1_37[137],stage1_36[181]}
   );
   gpc615_5 gpc1464 (
      {stage0_36[347], stage0_36[348], stage0_36[349], stage0_36[350], stage0_36[351]},
      {stage0_37[142]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[66],stage1_38[82],stage1_37[138],stage1_36[182]}
   );
   gpc615_5 gpc1465 (
      {stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355], stage0_36[356]},
      {stage0_37[143]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[67],stage1_38[83],stage1_37[139],stage1_36[183]}
   );
   gpc615_5 gpc1466 (
      {stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_37[144]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[68],stage1_38[84],stage1_37[140],stage1_36[184]}
   );
   gpc615_5 gpc1467 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366]},
      {stage0_37[145]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[69],stage1_38[85],stage1_37[141],stage1_36[185]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150], stage0_37[151]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[47],stage1_39[70],stage1_38[86],stage1_37[142]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156], stage0_37[157]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[48],stage1_39[71],stage1_38[87],stage1_37[143]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162], stage0_37[163]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[49],stage1_39[72],stage1_38[88],stage1_37[144]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168], stage0_37[169]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[50],stage1_39[73],stage1_38[89],stage1_37[145]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174], stage0_37[175]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[51],stage1_39[74],stage1_38[90],stage1_37[146]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180], stage0_37[181]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[52],stage1_39[75],stage1_38[91],stage1_37[147]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186], stage0_37[187]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[53],stage1_39[76],stage1_38[92],stage1_37[148]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192], stage0_37[193]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[54],stage1_39[77],stage1_38[93],stage1_37[149]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198], stage0_37[199]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[55],stage1_39[78],stage1_38[94],stage1_37[150]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204], stage0_37[205]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[56],stage1_39[79],stage1_38[95],stage1_37[151]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210], stage0_37[211]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[57],stage1_39[80],stage1_38[96],stage1_37[152]}
   );
   gpc606_5 gpc1479 (
      {stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216], stage0_37[217]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[58],stage1_39[81],stage1_38[97],stage1_37[153]}
   );
   gpc606_5 gpc1480 (
      {stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222], stage0_37[223]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[59],stage1_39[82],stage1_38[98],stage1_37[154]}
   );
   gpc606_5 gpc1481 (
      {stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228], stage0_37[229]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[60],stage1_39[83],stage1_38[99],stage1_37[155]}
   );
   gpc606_5 gpc1482 (
      {stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234], stage0_37[235]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[61],stage1_39[84],stage1_38[100],stage1_37[156]}
   );
   gpc606_5 gpc1483 (
      {stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240], stage0_37[241]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[62],stage1_39[85],stage1_38[101],stage1_37[157]}
   );
   gpc606_5 gpc1484 (
      {stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246], stage0_37[247]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[63],stage1_39[86],stage1_38[102],stage1_37[158]}
   );
   gpc606_5 gpc1485 (
      {stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252], stage0_37[253]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[64],stage1_39[87],stage1_38[103],stage1_37[159]}
   );
   gpc606_5 gpc1486 (
      {stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258], stage0_37[259]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[65],stage1_39[88],stage1_38[104],stage1_37[160]}
   );
   gpc606_5 gpc1487 (
      {stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264], stage0_37[265]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[66],stage1_39[89],stage1_38[105],stage1_37[161]}
   );
   gpc606_5 gpc1488 (
      {stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270], stage0_37[271]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[67],stage1_39[90],stage1_38[106],stage1_37[162]}
   );
   gpc606_5 gpc1489 (
      {stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276], stage0_37[277]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[68],stage1_39[91],stage1_38[107],stage1_37[163]}
   );
   gpc606_5 gpc1490 (
      {stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282], stage0_37[283]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[69],stage1_39[92],stage1_38[108],stage1_37[164]}
   );
   gpc606_5 gpc1491 (
      {stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288], stage0_37[289]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[70],stage1_39[93],stage1_38[109],stage1_37[165]}
   );
   gpc606_5 gpc1492 (
      {stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294], stage0_37[295]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[71],stage1_39[94],stage1_38[110],stage1_37[166]}
   );
   gpc606_5 gpc1493 (
      {stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300], stage0_37[301]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[72],stage1_39[95],stage1_38[111],stage1_37[167]}
   );
   gpc606_5 gpc1494 (
      {stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306], stage0_37[307]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[73],stage1_39[96],stage1_38[112],stage1_37[168]}
   );
   gpc606_5 gpc1495 (
      {stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312], stage0_37[313]},
      {stage0_39[162], stage0_39[163], stage0_39[164], stage0_39[165], stage0_39[166], stage0_39[167]},
      {stage1_41[27],stage1_40[74],stage1_39[97],stage1_38[113],stage1_37[169]}
   );
   gpc606_5 gpc1496 (
      {stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318], stage0_37[319]},
      {stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171], stage0_39[172], stage0_39[173]},
      {stage1_41[28],stage1_40[75],stage1_39[98],stage1_38[114],stage1_37[170]}
   );
   gpc606_5 gpc1497 (
      {stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324], stage0_37[325]},
      {stage0_39[174], stage0_39[175], stage0_39[176], stage0_39[177], stage0_39[178], stage0_39[179]},
      {stage1_41[29],stage1_40[76],stage1_39[99],stage1_38[115],stage1_37[171]}
   );
   gpc606_5 gpc1498 (
      {stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330], stage0_37[331]},
      {stage0_39[180], stage0_39[181], stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185]},
      {stage1_41[30],stage1_40[77],stage1_39[100],stage1_38[116],stage1_37[172]}
   );
   gpc606_5 gpc1499 (
      {stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336], stage0_37[337]},
      {stage0_39[186], stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage1_41[31],stage1_40[78],stage1_39[101],stage1_38[117],stage1_37[173]}
   );
   gpc606_5 gpc1500 (
      {stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342], stage0_37[343]},
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196], stage0_39[197]},
      {stage1_41[32],stage1_40[79],stage1_39[102],stage1_38[118],stage1_37[174]}
   );
   gpc606_5 gpc1501 (
      {stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348], stage0_37[349]},
      {stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201], stage0_39[202], stage0_39[203]},
      {stage1_41[33],stage1_40[80],stage1_39[103],stage1_38[119],stage1_37[175]}
   );
   gpc606_5 gpc1502 (
      {stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354], stage0_37[355]},
      {stage0_39[204], stage0_39[205], stage0_39[206], stage0_39[207], stage0_39[208], stage0_39[209]},
      {stage1_41[34],stage1_40[81],stage1_39[104],stage1_38[120],stage1_37[176]}
   );
   gpc606_5 gpc1503 (
      {stage0_37[356], stage0_37[357], stage0_37[358], stage0_37[359], stage0_37[360], stage0_37[361]},
      {stage0_39[210], stage0_39[211], stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215]},
      {stage1_41[35],stage1_40[82],stage1_39[105],stage1_38[121],stage1_37[177]}
   );
   gpc606_5 gpc1504 (
      {stage0_37[362], stage0_37[363], stage0_37[364], stage0_37[365], stage0_37[366], stage0_37[367]},
      {stage0_39[216], stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage1_41[36],stage1_40[83],stage1_39[106],stage1_38[122],stage1_37[178]}
   );
   gpc606_5 gpc1505 (
      {stage0_37[368], stage0_37[369], stage0_37[370], stage0_37[371], stage0_37[372], stage0_37[373]},
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226], stage0_39[227]},
      {stage1_41[37],stage1_40[84],stage1_39[107],stage1_38[123],stage1_37[179]}
   );
   gpc606_5 gpc1506 (
      {stage0_37[374], stage0_37[375], stage0_37[376], stage0_37[377], stage0_37[378], stage0_37[379]},
      {stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231], stage0_39[232], stage0_39[233]},
      {stage1_41[38],stage1_40[85],stage1_39[108],stage1_38[124],stage1_37[180]}
   );
   gpc606_5 gpc1507 (
      {stage0_37[380], stage0_37[381], stage0_37[382], stage0_37[383], stage0_37[384], stage0_37[385]},
      {stage0_39[234], stage0_39[235], stage0_39[236], stage0_39[237], stage0_39[238], stage0_39[239]},
      {stage1_41[39],stage1_40[86],stage1_39[109],stage1_38[125],stage1_37[181]}
   );
   gpc606_5 gpc1508 (
      {stage0_37[386], stage0_37[387], stage0_37[388], stage0_37[389], stage0_37[390], stage0_37[391]},
      {stage0_39[240], stage0_39[241], stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245]},
      {stage1_41[40],stage1_40[87],stage1_39[110],stage1_38[126],stage1_37[182]}
   );
   gpc615_5 gpc1509 (
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286]},
      {stage0_39[246]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[41],stage1_40[88],stage1_39[111],stage1_38[127]}
   );
   gpc615_5 gpc1510 (
      {stage0_38[287], stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291]},
      {stage0_39[247]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[42],stage1_40[89],stage1_39[112],stage1_38[128]}
   );
   gpc615_5 gpc1511 (
      {stage0_38[292], stage0_38[293], stage0_38[294], stage0_38[295], stage0_38[296]},
      {stage0_39[248]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[43],stage1_40[90],stage1_39[113],stage1_38[129]}
   );
   gpc615_5 gpc1512 (
      {stage0_38[297], stage0_38[298], stage0_38[299], stage0_38[300], stage0_38[301]},
      {stage0_39[249]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[44],stage1_40[91],stage1_39[114],stage1_38[130]}
   );
   gpc615_5 gpc1513 (
      {stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305], stage0_38[306]},
      {stage0_39[250]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[45],stage1_40[92],stage1_39[115],stage1_38[131]}
   );
   gpc615_5 gpc1514 (
      {stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage0_39[251]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[46],stage1_40[93],stage1_39[116],stage1_38[132]}
   );
   gpc615_5 gpc1515 (
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316]},
      {stage0_39[252]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[47],stage1_40[94],stage1_39[117],stage1_38[133]}
   );
   gpc615_5 gpc1516 (
      {stage0_38[317], stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321]},
      {stage0_39[253]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[48],stage1_40[95],stage1_39[118],stage1_38[134]}
   );
   gpc615_5 gpc1517 (
      {stage0_38[322], stage0_38[323], stage0_38[324], stage0_38[325], stage0_38[326]},
      {stage0_39[254]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[49],stage1_40[96],stage1_39[119],stage1_38[135]}
   );
   gpc615_5 gpc1518 (
      {stage0_38[327], stage0_38[328], stage0_38[329], stage0_38[330], stage0_38[331]},
      {stage0_39[255]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[50],stage1_40[97],stage1_39[120],stage1_38[136]}
   );
   gpc615_5 gpc1519 (
      {stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335], stage0_38[336]},
      {stage0_39[256]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[51],stage1_40[98],stage1_39[121],stage1_38[137]}
   );
   gpc615_5 gpc1520 (
      {stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage0_39[257]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[52],stage1_40[99],stage1_39[122],stage1_38[138]}
   );
   gpc615_5 gpc1521 (
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346]},
      {stage0_39[258]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[53],stage1_40[100],stage1_39[123],stage1_38[139]}
   );
   gpc615_5 gpc1522 (
      {stage0_38[347], stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351]},
      {stage0_39[259]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[54],stage1_40[101],stage1_39[124],stage1_38[140]}
   );
   gpc615_5 gpc1523 (
      {stage0_38[352], stage0_38[353], stage0_38[354], stage0_38[355], stage0_38[356]},
      {stage0_39[260]},
      {stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89]},
      {stage1_42[14],stage1_41[55],stage1_40[102],stage1_39[125],stage1_38[141]}
   );
   gpc615_5 gpc1524 (
      {stage0_38[357], stage0_38[358], stage0_38[359], stage0_38[360], stage0_38[361]},
      {stage0_39[261]},
      {stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95]},
      {stage1_42[15],stage1_41[56],stage1_40[103],stage1_39[126],stage1_38[142]}
   );
   gpc615_5 gpc1525 (
      {stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365], stage0_38[366]},
      {stage0_39[262]},
      {stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101]},
      {stage1_42[16],stage1_41[57],stage1_40[104],stage1_39[127],stage1_38[143]}
   );
   gpc615_5 gpc1526 (
      {stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370], stage0_38[371]},
      {stage0_39[263]},
      {stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107]},
      {stage1_42[17],stage1_41[58],stage1_40[105],stage1_39[128],stage1_38[144]}
   );
   gpc615_5 gpc1527 (
      {stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375], stage0_38[376]},
      {stage0_39[264]},
      {stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113]},
      {stage1_42[18],stage1_41[59],stage1_40[106],stage1_39[129],stage1_38[145]}
   );
   gpc615_5 gpc1528 (
      {stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380], stage0_38[381]},
      {stage0_39[265]},
      {stage0_40[114], stage0_40[115], stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119]},
      {stage1_42[19],stage1_41[60],stage1_40[107],stage1_39[130],stage1_38[146]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[266], stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270]},
      {stage0_40[120]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[20],stage1_41[61],stage1_40[108],stage1_39[131]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[271], stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275]},
      {stage0_40[121]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[21],stage1_41[62],stage1_40[109],stage1_39[132]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[276], stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280]},
      {stage0_40[122]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[22],stage1_41[63],stage1_40[110],stage1_39[133]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[281], stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285]},
      {stage0_40[123]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[23],stage1_41[64],stage1_40[111],stage1_39[134]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[286], stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290]},
      {stage0_40[124]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[24],stage1_41[65],stage1_40[112],stage1_39[135]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[291], stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295]},
      {stage0_40[125]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[25],stage1_41[66],stage1_40[113],stage1_39[136]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[296], stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300]},
      {stage0_40[126]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[26],stage1_41[67],stage1_40[114],stage1_39[137]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[301], stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305]},
      {stage0_40[127]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[27],stage1_41[68],stage1_40[115],stage1_39[138]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[306], stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310]},
      {stage0_40[128]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[28],stage1_41[69],stage1_40[116],stage1_39[139]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[311], stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315]},
      {stage0_40[129]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[29],stage1_41[70],stage1_40[117],stage1_39[140]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[316], stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320]},
      {stage0_40[130]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[30],stage1_41[71],stage1_40[118],stage1_39[141]}
   );
   gpc615_5 gpc1540 (
      {stage0_39[321], stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325]},
      {stage0_40[131]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[31],stage1_41[72],stage1_40[119],stage1_39[142]}
   );
   gpc615_5 gpc1541 (
      {stage0_39[326], stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330]},
      {stage0_40[132]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[32],stage1_41[73],stage1_40[120],stage1_39[143]}
   );
   gpc615_5 gpc1542 (
      {stage0_39[331], stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335]},
      {stage0_40[133]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[33],stage1_41[74],stage1_40[121],stage1_39[144]}
   );
   gpc615_5 gpc1543 (
      {stage0_39[336], stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340]},
      {stage0_40[134]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[34],stage1_41[75],stage1_40[122],stage1_39[145]}
   );
   gpc615_5 gpc1544 (
      {stage0_39[341], stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345]},
      {stage0_40[135]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[35],stage1_41[76],stage1_40[123],stage1_39[146]}
   );
   gpc615_5 gpc1545 (
      {stage0_39[346], stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350]},
      {stage0_40[136]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[36],stage1_41[77],stage1_40[124],stage1_39[147]}
   );
   gpc615_5 gpc1546 (
      {stage0_39[351], stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355]},
      {stage0_40[137]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[37],stage1_41[78],stage1_40[125],stage1_39[148]}
   );
   gpc615_5 gpc1547 (
      {stage0_39[356], stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360]},
      {stage0_40[138]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[38],stage1_41[79],stage1_40[126],stage1_39[149]}
   );
   gpc615_5 gpc1548 (
      {stage0_39[361], stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365]},
      {stage0_40[139]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[39],stage1_41[80],stage1_40[127],stage1_39[150]}
   );
   gpc615_5 gpc1549 (
      {stage0_39[366], stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370]},
      {stage0_40[140]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[40],stage1_41[81],stage1_40[128],stage1_39[151]}
   );
   gpc615_5 gpc1550 (
      {stage0_39[371], stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375]},
      {stage0_40[141]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[41],stage1_41[82],stage1_40[129],stage1_39[152]}
   );
   gpc615_5 gpc1551 (
      {stage0_39[376], stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380]},
      {stage0_40[142]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[42],stage1_41[83],stage1_40[130],stage1_39[153]}
   );
   gpc615_5 gpc1552 (
      {stage0_39[381], stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385]},
      {stage0_40[143]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[43],stage1_41[84],stage1_40[131],stage1_39[154]}
   );
   gpc615_5 gpc1553 (
      {stage0_39[386], stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390]},
      {stage0_40[144]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[44],stage1_41[85],stage1_40[132],stage1_39[155]}
   );
   gpc615_5 gpc1554 (
      {stage0_39[391], stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395]},
      {stage0_40[145]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[45],stage1_41[86],stage1_40[133],stage1_39[156]}
   );
   gpc615_5 gpc1555 (
      {stage0_39[396], stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400]},
      {stage0_40[146]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[46],stage1_41[87],stage1_40[134],stage1_39[157]}
   );
   gpc615_5 gpc1556 (
      {stage0_39[401], stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405]},
      {stage0_40[147]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[47],stage1_41[88],stage1_40[135],stage1_39[158]}
   );
   gpc615_5 gpc1557 (
      {stage0_39[406], stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410]},
      {stage0_40[148]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[48],stage1_41[89],stage1_40[136],stage1_39[159]}
   );
   gpc615_5 gpc1558 (
      {stage0_39[411], stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415]},
      {stage0_40[149]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[49],stage1_41[90],stage1_40[137],stage1_39[160]}
   );
   gpc615_5 gpc1559 (
      {stage0_39[416], stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420]},
      {stage0_40[150]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[50],stage1_41[91],stage1_40[138],stage1_39[161]}
   );
   gpc615_5 gpc1560 (
      {stage0_39[421], stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425]},
      {stage0_40[151]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[51],stage1_41[92],stage1_40[139],stage1_39[162]}
   );
   gpc615_5 gpc1561 (
      {stage0_39[426], stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430]},
      {stage0_40[152]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[52],stage1_41[93],stage1_40[140],stage1_39[163]}
   );
   gpc615_5 gpc1562 (
      {stage0_39[431], stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435]},
      {stage0_40[153]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[53],stage1_41[94],stage1_40[141],stage1_39[164]}
   );
   gpc615_5 gpc1563 (
      {stage0_39[436], stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440]},
      {stage0_40[154]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[54],stage1_41[95],stage1_40[142],stage1_39[165]}
   );
   gpc615_5 gpc1564 (
      {stage0_39[441], stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445]},
      {stage0_40[155]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[55],stage1_41[96],stage1_40[143],stage1_39[166]}
   );
   gpc615_5 gpc1565 (
      {stage0_39[446], stage0_39[447], stage0_39[448], stage0_39[449], stage0_39[450]},
      {stage0_40[156]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[56],stage1_41[97],stage1_40[144],stage1_39[167]}
   );
   gpc615_5 gpc1566 (
      {stage0_39[451], stage0_39[452], stage0_39[453], stage0_39[454], stage0_39[455]},
      {stage0_40[157]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[57],stage1_41[98],stage1_40[145],stage1_39[168]}
   );
   gpc615_5 gpc1567 (
      {stage0_39[456], stage0_39[457], stage0_39[458], stage0_39[459], stage0_39[460]},
      {stage0_40[158]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[58],stage1_41[99],stage1_40[146],stage1_39[169]}
   );
   gpc615_5 gpc1568 (
      {stage0_39[461], stage0_39[462], stage0_39[463], stage0_39[464], stage0_39[465]},
      {stage0_40[159]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[59],stage1_41[100],stage1_40[147],stage1_39[170]}
   );
   gpc615_5 gpc1569 (
      {stage0_39[466], stage0_39[467], stage0_39[468], stage0_39[469], stage0_39[470]},
      {stage0_40[160]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[60],stage1_41[101],stage1_40[148],stage1_39[171]}
   );
   gpc615_5 gpc1570 (
      {stage0_39[471], stage0_39[472], stage0_39[473], stage0_39[474], stage0_39[475]},
      {stage0_40[161]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[61],stage1_41[102],stage1_40[149],stage1_39[172]}
   );
   gpc615_5 gpc1571 (
      {stage0_39[476], stage0_39[477], stage0_39[478], stage0_39[479], stage0_39[480]},
      {stage0_40[162]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[62],stage1_41[103],stage1_40[150],stage1_39[173]}
   );
   gpc615_5 gpc1572 (
      {stage0_39[481], stage0_39[482], stage0_39[483], stage0_39[484], stage0_39[485]},
      {stage0_40[163]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[63],stage1_41[104],stage1_40[151],stage1_39[174]}
   );
   gpc615_5 gpc1573 (
      {stage0_39[486], stage0_39[487], stage0_39[488], stage0_39[489], stage0_39[490]},
      {stage0_40[164]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[64],stage1_41[105],stage1_40[152],stage1_39[175]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169], stage0_40[170]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[45],stage1_42[65],stage1_41[106],stage1_40[153]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175], stage0_40[176]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[46],stage1_42[66],stage1_41[107],stage1_40[154]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181], stage0_40[182]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[47],stage1_42[67],stage1_41[108],stage1_40[155]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187], stage0_40[188]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[48],stage1_42[68],stage1_41[109],stage1_40[156]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193], stage0_40[194]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[49],stage1_42[69],stage1_41[110],stage1_40[157]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199], stage0_40[200]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[50],stage1_42[70],stage1_41[111],stage1_40[158]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205], stage0_40[206]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[51],stage1_42[71],stage1_41[112],stage1_40[159]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211], stage0_40[212]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[52],stage1_42[72],stage1_41[113],stage1_40[160]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217], stage0_40[218]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[53],stage1_42[73],stage1_41[114],stage1_40[161]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223], stage0_40[224]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[54],stage1_42[74],stage1_41[115],stage1_40[162]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229], stage0_40[230]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[55],stage1_42[75],stage1_41[116],stage1_40[163]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235], stage0_40[236]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[56],stage1_42[76],stage1_41[117],stage1_40[164]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241], stage0_40[242]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[57],stage1_42[77],stage1_41[118],stage1_40[165]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247], stage0_40[248]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[58],stage1_42[78],stage1_41[119],stage1_40[166]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253], stage0_40[254]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[59],stage1_42[79],stage1_41[120],stage1_40[167]}
   );
   gpc606_5 gpc1589 (
      {stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259], stage0_40[260]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[60],stage1_42[80],stage1_41[121],stage1_40[168]}
   );
   gpc606_5 gpc1590 (
      {stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265], stage0_40[266]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[61],stage1_42[81],stage1_41[122],stage1_40[169]}
   );
   gpc606_5 gpc1591 (
      {stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271], stage0_40[272]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[62],stage1_42[82],stage1_41[123],stage1_40[170]}
   );
   gpc606_5 gpc1592 (
      {stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277], stage0_40[278]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[63],stage1_42[83],stage1_41[124],stage1_40[171]}
   );
   gpc606_5 gpc1593 (
      {stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283], stage0_40[284]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[64],stage1_42[84],stage1_41[125],stage1_40[172]}
   );
   gpc606_5 gpc1594 (
      {stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289], stage0_40[290]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[65],stage1_42[85],stage1_41[126],stage1_40[173]}
   );
   gpc606_5 gpc1595 (
      {stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295], stage0_40[296]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[66],stage1_42[86],stage1_41[127],stage1_40[174]}
   );
   gpc606_5 gpc1596 (
      {stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301], stage0_40[302]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[67],stage1_42[87],stage1_41[128],stage1_40[175]}
   );
   gpc606_5 gpc1597 (
      {stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307], stage0_40[308]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[68],stage1_42[88],stage1_41[129],stage1_40[176]}
   );
   gpc606_5 gpc1598 (
      {stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313], stage0_40[314]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[69],stage1_42[89],stage1_41[130],stage1_40[177]}
   );
   gpc606_5 gpc1599 (
      {stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319], stage0_40[320]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[70],stage1_42[90],stage1_41[131],stage1_40[178]}
   );
   gpc606_5 gpc1600 (
      {stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325], stage0_40[326]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[71],stage1_42[91],stage1_41[132],stage1_40[179]}
   );
   gpc606_5 gpc1601 (
      {stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331], stage0_40[332]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[72],stage1_42[92],stage1_41[133],stage1_40[180]}
   );
   gpc606_5 gpc1602 (
      {stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337], stage0_40[338]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[73],stage1_42[93],stage1_41[134],stage1_40[181]}
   );
   gpc606_5 gpc1603 (
      {stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343], stage0_40[344]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[74],stage1_42[94],stage1_41[135],stage1_40[182]}
   );
   gpc606_5 gpc1604 (
      {stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349], stage0_40[350]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[75],stage1_42[95],stage1_41[136],stage1_40[183]}
   );
   gpc606_5 gpc1605 (
      {stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355], stage0_40[356]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[76],stage1_42[96],stage1_41[137],stage1_40[184]}
   );
   gpc606_5 gpc1606 (
      {stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361], stage0_40[362]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[77],stage1_42[97],stage1_41[138],stage1_40[185]}
   );
   gpc606_5 gpc1607 (
      {stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367], stage0_40[368]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[78],stage1_42[98],stage1_41[139],stage1_40[186]}
   );
   gpc606_5 gpc1608 (
      {stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373], stage0_40[374]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[79],stage1_42[99],stage1_41[140],stage1_40[187]}
   );
   gpc606_5 gpc1609 (
      {stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379], stage0_40[380]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[80],stage1_42[100],stage1_41[141],stage1_40[188]}
   );
   gpc606_5 gpc1610 (
      {stage0_40[381], stage0_40[382], stage0_40[383], stage0_40[384], stage0_40[385], stage0_40[386]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[81],stage1_42[101],stage1_41[142],stage1_40[189]}
   );
   gpc606_5 gpc1611 (
      {stage0_40[387], stage0_40[388], stage0_40[389], stage0_40[390], stage0_40[391], stage0_40[392]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[82],stage1_42[102],stage1_41[143],stage1_40[190]}
   );
   gpc606_5 gpc1612 (
      {stage0_40[393], stage0_40[394], stage0_40[395], stage0_40[396], stage0_40[397], stage0_40[398]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[83],stage1_42[103],stage1_41[144],stage1_40[191]}
   );
   gpc606_5 gpc1613 (
      {stage0_40[399], stage0_40[400], stage0_40[401], stage0_40[402], stage0_40[403], stage0_40[404]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[84],stage1_42[104],stage1_41[145],stage1_40[192]}
   );
   gpc606_5 gpc1614 (
      {stage0_40[405], stage0_40[406], stage0_40[407], stage0_40[408], stage0_40[409], stage0_40[410]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[85],stage1_42[105],stage1_41[146],stage1_40[193]}
   );
   gpc606_5 gpc1615 (
      {stage0_40[411], stage0_40[412], stage0_40[413], stage0_40[414], stage0_40[415], stage0_40[416]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[86],stage1_42[106],stage1_41[147],stage1_40[194]}
   );
   gpc606_5 gpc1616 (
      {stage0_40[417], stage0_40[418], stage0_40[419], stage0_40[420], stage0_40[421], stage0_40[422]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[87],stage1_42[107],stage1_41[148],stage1_40[195]}
   );
   gpc606_5 gpc1617 (
      {stage0_40[423], stage0_40[424], stage0_40[425], stage0_40[426], stage0_40[427], stage0_40[428]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[88],stage1_42[108],stage1_41[149],stage1_40[196]}
   );
   gpc606_5 gpc1618 (
      {stage0_40[429], stage0_40[430], stage0_40[431], stage0_40[432], stage0_40[433], stage0_40[434]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[89],stage1_42[109],stage1_41[150],stage1_40[197]}
   );
   gpc606_5 gpc1619 (
      {stage0_40[435], stage0_40[436], stage0_40[437], stage0_40[438], stage0_40[439], stage0_40[440]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[90],stage1_42[110],stage1_41[151],stage1_40[198]}
   );
   gpc606_5 gpc1620 (
      {stage0_40[441], stage0_40[442], stage0_40[443], stage0_40[444], stage0_40[445], stage0_40[446]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[91],stage1_42[111],stage1_41[152],stage1_40[199]}
   );
   gpc606_5 gpc1621 (
      {stage0_40[447], stage0_40[448], stage0_40[449], stage0_40[450], stage0_40[451], stage0_40[452]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[92],stage1_42[112],stage1_41[153],stage1_40[200]}
   );
   gpc606_5 gpc1622 (
      {stage0_40[453], stage0_40[454], stage0_40[455], stage0_40[456], stage0_40[457], stage0_40[458]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[93],stage1_42[113],stage1_41[154],stage1_40[201]}
   );
   gpc606_5 gpc1623 (
      {stage0_40[459], stage0_40[460], stage0_40[461], stage0_40[462], stage0_40[463], stage0_40[464]},
      {stage0_42[294], stage0_42[295], stage0_42[296], stage0_42[297], stage0_42[298], stage0_42[299]},
      {stage1_44[49],stage1_43[94],stage1_42[114],stage1_41[155],stage1_40[202]}
   );
   gpc606_5 gpc1624 (
      {stage0_40[465], stage0_40[466], stage0_40[467], stage0_40[468], stage0_40[469], stage0_40[470]},
      {stage0_42[300], stage0_42[301], stage0_42[302], stage0_42[303], stage0_42[304], stage0_42[305]},
      {stage1_44[50],stage1_43[95],stage1_42[115],stage1_41[156],stage1_40[203]}
   );
   gpc606_5 gpc1625 (
      {stage0_40[471], stage0_40[472], stage0_40[473], stage0_40[474], stage0_40[475], stage0_40[476]},
      {stage0_42[306], stage0_42[307], stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311]},
      {stage1_44[51],stage1_43[96],stage1_42[116],stage1_41[157],stage1_40[204]}
   );
   gpc606_5 gpc1626 (
      {stage0_40[477], stage0_40[478], stage0_40[479], stage0_40[480], stage0_40[481], stage0_40[482]},
      {stage0_42[312], stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage1_44[52],stage1_43[97],stage1_42[117],stage1_41[158],stage1_40[205]}
   );
   gpc606_5 gpc1627 (
      {stage0_40[483], stage0_40[484], stage0_40[485], stage0_40[486], stage0_40[487], stage0_40[488]},
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322], stage0_42[323]},
      {stage1_44[53],stage1_43[98],stage1_42[118],stage1_41[159],stage1_40[206]}
   );
   gpc606_5 gpc1628 (
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[54],stage1_43[99],stage1_42[119],stage1_41[160]}
   );
   gpc606_5 gpc1629 (
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[55],stage1_43[100],stage1_42[120],stage1_41[161]}
   );
   gpc606_5 gpc1630 (
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[56],stage1_43[101],stage1_42[121],stage1_41[162]}
   );
   gpc606_5 gpc1631 (
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[57],stage1_43[102],stage1_42[122],stage1_41[163]}
   );
   gpc606_5 gpc1632 (
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[58],stage1_43[103],stage1_42[123],stage1_41[164]}
   );
   gpc606_5 gpc1633 (
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[59],stage1_43[104],stage1_42[124],stage1_41[165]}
   );
   gpc606_5 gpc1634 (
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[60],stage1_43[105],stage1_42[125],stage1_41[166]}
   );
   gpc606_5 gpc1635 (
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[61],stage1_43[106],stage1_42[126],stage1_41[167]}
   );
   gpc606_5 gpc1636 (
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[62],stage1_43[107],stage1_42[127],stage1_41[168]}
   );
   gpc606_5 gpc1637 (
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[63],stage1_43[108],stage1_42[128],stage1_41[169]}
   );
   gpc606_5 gpc1638 (
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[64],stage1_43[109],stage1_42[129],stage1_41[170]}
   );
   gpc606_5 gpc1639 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[65],stage1_43[110],stage1_42[130],stage1_41[171]}
   );
   gpc606_5 gpc1640 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[66],stage1_43[111],stage1_42[131],stage1_41[172]}
   );
   gpc606_5 gpc1641 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[67],stage1_43[112],stage1_42[132],stage1_41[173]}
   );
   gpc606_5 gpc1642 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[68],stage1_43[113],stage1_42[133],stage1_41[174]}
   );
   gpc606_5 gpc1643 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[69],stage1_43[114],stage1_42[134],stage1_41[175]}
   );
   gpc606_5 gpc1644 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[70],stage1_43[115],stage1_42[135],stage1_41[176]}
   );
   gpc606_5 gpc1645 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[71],stage1_43[116],stage1_42[136],stage1_41[177]}
   );
   gpc606_5 gpc1646 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[72],stage1_43[117],stage1_42[137],stage1_41[178]}
   );
   gpc606_5 gpc1647 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[73],stage1_43[118],stage1_42[138],stage1_41[179]}
   );
   gpc606_5 gpc1648 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[74],stage1_43[119],stage1_42[139],stage1_41[180]}
   );
   gpc606_5 gpc1649 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[75],stage1_43[120],stage1_42[140],stage1_41[181]}
   );
   gpc606_5 gpc1650 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[76],stage1_43[121],stage1_42[141],stage1_41[182]}
   );
   gpc606_5 gpc1651 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[77],stage1_43[122],stage1_42[142],stage1_41[183]}
   );
   gpc606_5 gpc1652 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[78],stage1_43[123],stage1_42[143],stage1_41[184]}
   );
   gpc606_5 gpc1653 (
      {stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327], stage0_42[328], stage0_42[329]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[79],stage1_43[124],stage1_42[144]}
   );
   gpc606_5 gpc1654 (
      {stage0_42[330], stage0_42[331], stage0_42[332], stage0_42[333], stage0_42[334], stage0_42[335]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[80],stage1_43[125],stage1_42[145]}
   );
   gpc606_5 gpc1655 (
      {stage0_42[336], stage0_42[337], stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[81],stage1_43[126],stage1_42[146]}
   );
   gpc606_5 gpc1656 (
      {stage0_42[342], stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[82],stage1_43[127],stage1_42[147]}
   );
   gpc606_5 gpc1657 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352], stage0_42[353]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[83],stage1_43[128],stage1_42[148]}
   );
   gpc606_5 gpc1658 (
      {stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357], stage0_42[358], stage0_42[359]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[84],stage1_43[129],stage1_42[149]}
   );
   gpc606_5 gpc1659 (
      {stage0_42[360], stage0_42[361], stage0_42[362], stage0_42[363], stage0_42[364], stage0_42[365]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[85],stage1_43[130],stage1_42[150]}
   );
   gpc615_5 gpc1660 (
      {stage0_42[366], stage0_42[367], stage0_42[368], stage0_42[369], stage0_42[370]},
      {stage0_43[150]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[86],stage1_43[131],stage1_42[151]}
   );
   gpc615_5 gpc1661 (
      {stage0_42[371], stage0_42[372], stage0_42[373], stage0_42[374], stage0_42[375]},
      {stage0_43[151]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[87],stage1_43[132],stage1_42[152]}
   );
   gpc615_5 gpc1662 (
      {stage0_42[376], stage0_42[377], stage0_42[378], stage0_42[379], stage0_42[380]},
      {stage0_43[152]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[88],stage1_43[133],stage1_42[153]}
   );
   gpc615_5 gpc1663 (
      {stage0_42[381], stage0_42[382], stage0_42[383], stage0_42[384], stage0_42[385]},
      {stage0_43[153]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[89],stage1_43[134],stage1_42[154]}
   );
   gpc615_5 gpc1664 (
      {stage0_42[386], stage0_42[387], stage0_42[388], stage0_42[389], stage0_42[390]},
      {stage0_43[154]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[90],stage1_43[135],stage1_42[155]}
   );
   gpc615_5 gpc1665 (
      {stage0_42[391], stage0_42[392], stage0_42[393], stage0_42[394], stage0_42[395]},
      {stage0_43[155]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[91],stage1_43[136],stage1_42[156]}
   );
   gpc615_5 gpc1666 (
      {stage0_42[396], stage0_42[397], stage0_42[398], stage0_42[399], stage0_42[400]},
      {stage0_43[156]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[92],stage1_43[137],stage1_42[157]}
   );
   gpc615_5 gpc1667 (
      {stage0_42[401], stage0_42[402], stage0_42[403], stage0_42[404], stage0_42[405]},
      {stage0_43[157]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[93],stage1_43[138],stage1_42[158]}
   );
   gpc615_5 gpc1668 (
      {stage0_42[406], stage0_42[407], stage0_42[408], stage0_42[409], stage0_42[410]},
      {stage0_43[158]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[94],stage1_43[139],stage1_42[159]}
   );
   gpc615_5 gpc1669 (
      {stage0_42[411], stage0_42[412], stage0_42[413], stage0_42[414], stage0_42[415]},
      {stage0_43[159]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[95],stage1_43[140],stage1_42[160]}
   );
   gpc615_5 gpc1670 (
      {stage0_42[416], stage0_42[417], stage0_42[418], stage0_42[419], stage0_42[420]},
      {stage0_43[160]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[96],stage1_43[141],stage1_42[161]}
   );
   gpc615_5 gpc1671 (
      {stage0_42[421], stage0_42[422], stage0_42[423], stage0_42[424], stage0_42[425]},
      {stage0_43[161]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[97],stage1_43[142],stage1_42[162]}
   );
   gpc615_5 gpc1672 (
      {stage0_42[426], stage0_42[427], stage0_42[428], stage0_42[429], stage0_42[430]},
      {stage0_43[162]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[98],stage1_43[143],stage1_42[163]}
   );
   gpc615_5 gpc1673 (
      {stage0_42[431], stage0_42[432], stage0_42[433], stage0_42[434], stage0_42[435]},
      {stage0_43[163]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[99],stage1_43[144],stage1_42[164]}
   );
   gpc615_5 gpc1674 (
      {stage0_42[436], stage0_42[437], stage0_42[438], stage0_42[439], stage0_42[440]},
      {stage0_43[164]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[100],stage1_43[145],stage1_42[165]}
   );
   gpc615_5 gpc1675 (
      {stage0_42[441], stage0_42[442], stage0_42[443], stage0_42[444], stage0_42[445]},
      {stage0_43[165]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[101],stage1_43[146],stage1_42[166]}
   );
   gpc615_5 gpc1676 (
      {stage0_42[446], stage0_42[447], stage0_42[448], stage0_42[449], stage0_42[450]},
      {stage0_43[166]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[102],stage1_43[147],stage1_42[167]}
   );
   gpc606_5 gpc1677 (
      {stage0_43[167], stage0_43[168], stage0_43[169], stage0_43[170], stage0_43[171], stage0_43[172]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[24],stage1_45[49],stage1_44[103],stage1_43[148]}
   );
   gpc606_5 gpc1678 (
      {stage0_43[173], stage0_43[174], stage0_43[175], stage0_43[176], stage0_43[177], stage0_43[178]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[25],stage1_45[50],stage1_44[104],stage1_43[149]}
   );
   gpc606_5 gpc1679 (
      {stage0_43[179], stage0_43[180], stage0_43[181], stage0_43[182], stage0_43[183], stage0_43[184]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[26],stage1_45[51],stage1_44[105],stage1_43[150]}
   );
   gpc606_5 gpc1680 (
      {stage0_43[185], stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[27],stage1_45[52],stage1_44[106],stage1_43[151]}
   );
   gpc606_5 gpc1681 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195], stage0_43[196]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[28],stage1_45[53],stage1_44[107],stage1_43[152]}
   );
   gpc606_5 gpc1682 (
      {stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200], stage0_43[201], stage0_43[202]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[29],stage1_45[54],stage1_44[108],stage1_43[153]}
   );
   gpc606_5 gpc1683 (
      {stage0_43[203], stage0_43[204], stage0_43[205], stage0_43[206], stage0_43[207], stage0_43[208]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[30],stage1_45[55],stage1_44[109],stage1_43[154]}
   );
   gpc606_5 gpc1684 (
      {stage0_43[209], stage0_43[210], stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[31],stage1_45[56],stage1_44[110],stage1_43[155]}
   );
   gpc606_5 gpc1685 (
      {stage0_43[215], stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[32],stage1_45[57],stage1_44[111],stage1_43[156]}
   );
   gpc606_5 gpc1686 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225], stage0_43[226]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[33],stage1_45[58],stage1_44[112],stage1_43[157]}
   );
   gpc606_5 gpc1687 (
      {stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230], stage0_43[231], stage0_43[232]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[34],stage1_45[59],stage1_44[113],stage1_43[158]}
   );
   gpc606_5 gpc1688 (
      {stage0_43[233], stage0_43[234], stage0_43[235], stage0_43[236], stage0_43[237], stage0_43[238]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[35],stage1_45[60],stage1_44[114],stage1_43[159]}
   );
   gpc606_5 gpc1689 (
      {stage0_43[239], stage0_43[240], stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[36],stage1_45[61],stage1_44[115],stage1_43[160]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[245], stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249]},
      {stage0_44[144]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[37],stage1_45[62],stage1_44[116],stage1_43[161]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[250], stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254]},
      {stage0_44[145]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[38],stage1_45[63],stage1_44[117],stage1_43[162]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[255], stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259]},
      {stage0_44[146]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[39],stage1_45[64],stage1_44[118],stage1_43[163]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[260], stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264]},
      {stage0_44[147]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[40],stage1_45[65],stage1_44[119],stage1_43[164]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[265], stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269]},
      {stage0_44[148]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[41],stage1_45[66],stage1_44[120],stage1_43[165]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[270], stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274]},
      {stage0_44[149]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[42],stage1_45[67],stage1_44[121],stage1_43[166]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[275], stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279]},
      {stage0_44[150]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[43],stage1_45[68],stage1_44[122],stage1_43[167]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[280], stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284]},
      {stage0_44[151]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[44],stage1_45[69],stage1_44[123],stage1_43[168]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[285], stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289]},
      {stage0_44[152]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[45],stage1_45[70],stage1_44[124],stage1_43[169]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[290], stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294]},
      {stage0_44[153]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[46],stage1_45[71],stage1_44[125],stage1_43[170]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[295], stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299]},
      {stage0_44[154]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[47],stage1_45[72],stage1_44[126],stage1_43[171]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[300], stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304]},
      {stage0_44[155]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[48],stage1_45[73],stage1_44[127],stage1_43[172]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[305], stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309]},
      {stage0_44[156]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[49],stage1_45[74],stage1_44[128],stage1_43[173]}
   );
   gpc615_5 gpc1703 (
      {stage0_43[310], stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314]},
      {stage0_44[157]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[50],stage1_45[75],stage1_44[129],stage1_43[174]}
   );
   gpc615_5 gpc1704 (
      {stage0_43[315], stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319]},
      {stage0_44[158]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[51],stage1_45[76],stage1_44[130],stage1_43[175]}
   );
   gpc615_5 gpc1705 (
      {stage0_43[320], stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324]},
      {stage0_44[159]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[52],stage1_45[77],stage1_44[131],stage1_43[176]}
   );
   gpc615_5 gpc1706 (
      {stage0_43[325], stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329]},
      {stage0_44[160]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[53],stage1_45[78],stage1_44[132],stage1_43[177]}
   );
   gpc615_5 gpc1707 (
      {stage0_43[330], stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334]},
      {stage0_44[161]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[54],stage1_45[79],stage1_44[133],stage1_43[178]}
   );
   gpc615_5 gpc1708 (
      {stage0_43[335], stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339]},
      {stage0_44[162]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[55],stage1_45[80],stage1_44[134],stage1_43[179]}
   );
   gpc615_5 gpc1709 (
      {stage0_43[340], stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344]},
      {stage0_44[163]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[56],stage1_45[81],stage1_44[135],stage1_43[180]}
   );
   gpc615_5 gpc1710 (
      {stage0_43[345], stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349]},
      {stage0_44[164]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[57],stage1_45[82],stage1_44[136],stage1_43[181]}
   );
   gpc615_5 gpc1711 (
      {stage0_43[350], stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354]},
      {stage0_44[165]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[58],stage1_45[83],stage1_44[137],stage1_43[182]}
   );
   gpc615_5 gpc1712 (
      {stage0_43[355], stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359]},
      {stage0_44[166]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[59],stage1_45[84],stage1_44[138],stage1_43[183]}
   );
   gpc615_5 gpc1713 (
      {stage0_43[360], stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364]},
      {stage0_44[167]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[60],stage1_45[85],stage1_44[139],stage1_43[184]}
   );
   gpc615_5 gpc1714 (
      {stage0_43[365], stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369]},
      {stage0_44[168]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[61],stage1_45[86],stage1_44[140],stage1_43[185]}
   );
   gpc615_5 gpc1715 (
      {stage0_43[370], stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374]},
      {stage0_44[169]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[62],stage1_45[87],stage1_44[141],stage1_43[186]}
   );
   gpc615_5 gpc1716 (
      {stage0_43[375], stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379]},
      {stage0_44[170]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[63],stage1_45[88],stage1_44[142],stage1_43[187]}
   );
   gpc615_5 gpc1717 (
      {stage0_43[380], stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384]},
      {stage0_44[171]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[64],stage1_45[89],stage1_44[143],stage1_43[188]}
   );
   gpc615_5 gpc1718 (
      {stage0_43[385], stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389]},
      {stage0_44[172]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[65],stage1_45[90],stage1_44[144],stage1_43[189]}
   );
   gpc615_5 gpc1719 (
      {stage0_43[390], stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394]},
      {stage0_44[173]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[66],stage1_45[91],stage1_44[145],stage1_43[190]}
   );
   gpc615_5 gpc1720 (
      {stage0_43[395], stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399]},
      {stage0_44[174]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[67],stage1_45[92],stage1_44[146],stage1_43[191]}
   );
   gpc615_5 gpc1721 (
      {stage0_43[400], stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404]},
      {stage0_44[175]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[68],stage1_45[93],stage1_44[147],stage1_43[192]}
   );
   gpc615_5 gpc1722 (
      {stage0_43[405], stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409]},
      {stage0_44[176]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[69],stage1_45[94],stage1_44[148],stage1_43[193]}
   );
   gpc615_5 gpc1723 (
      {stage0_43[410], stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414]},
      {stage0_44[177]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[70],stage1_45[95],stage1_44[149],stage1_43[194]}
   );
   gpc615_5 gpc1724 (
      {stage0_43[415], stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419]},
      {stage0_44[178]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[71],stage1_45[96],stage1_44[150],stage1_43[195]}
   );
   gpc615_5 gpc1725 (
      {stage0_43[420], stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424]},
      {stage0_44[179]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[72],stage1_45[97],stage1_44[151],stage1_43[196]}
   );
   gpc615_5 gpc1726 (
      {stage0_43[425], stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429]},
      {stage0_44[180]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[73],stage1_45[98],stage1_44[152],stage1_43[197]}
   );
   gpc615_5 gpc1727 (
      {stage0_43[430], stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434]},
      {stage0_44[181]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[74],stage1_45[99],stage1_44[153],stage1_43[198]}
   );
   gpc615_5 gpc1728 (
      {stage0_43[435], stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439]},
      {stage0_44[182]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[75],stage1_45[100],stage1_44[154],stage1_43[199]}
   );
   gpc615_5 gpc1729 (
      {stage0_43[440], stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444]},
      {stage0_44[183]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[76],stage1_45[101],stage1_44[155],stage1_43[200]}
   );
   gpc615_5 gpc1730 (
      {stage0_43[445], stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449]},
      {stage0_44[184]},
      {stage0_45[318], stage0_45[319], stage0_45[320], stage0_45[321], stage0_45[322], stage0_45[323]},
      {stage1_47[53],stage1_46[77],stage1_45[102],stage1_44[156],stage1_43[201]}
   );
   gpc615_5 gpc1731 (
      {stage0_43[450], stage0_43[451], stage0_43[452], stage0_43[453], stage0_43[454]},
      {stage0_44[185]},
      {stage0_45[324], stage0_45[325], stage0_45[326], stage0_45[327], stage0_45[328], stage0_45[329]},
      {stage1_47[54],stage1_46[78],stage1_45[103],stage1_44[157],stage1_43[202]}
   );
   gpc615_5 gpc1732 (
      {stage0_43[455], stage0_43[456], stage0_43[457], stage0_43[458], stage0_43[459]},
      {stage0_44[186]},
      {stage0_45[330], stage0_45[331], stage0_45[332], stage0_45[333], stage0_45[334], stage0_45[335]},
      {stage1_47[55],stage1_46[79],stage1_45[104],stage1_44[158],stage1_43[203]}
   );
   gpc615_5 gpc1733 (
      {stage0_43[460], stage0_43[461], stage0_43[462], stage0_43[463], stage0_43[464]},
      {stage0_44[187]},
      {stage0_45[336], stage0_45[337], stage0_45[338], stage0_45[339], stage0_45[340], stage0_45[341]},
      {stage1_47[56],stage1_46[80],stage1_45[105],stage1_44[159],stage1_43[204]}
   );
   gpc615_5 gpc1734 (
      {stage0_43[465], stage0_43[466], stage0_43[467], stage0_43[468], stage0_43[469]},
      {stage0_44[188]},
      {stage0_45[342], stage0_45[343], stage0_45[344], stage0_45[345], stage0_45[346], stage0_45[347]},
      {stage1_47[57],stage1_46[81],stage1_45[106],stage1_44[160],stage1_43[205]}
   );
   gpc615_5 gpc1735 (
      {stage0_43[470], stage0_43[471], stage0_43[472], stage0_43[473], stage0_43[474]},
      {stage0_44[189]},
      {stage0_45[348], stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353]},
      {stage1_47[58],stage1_46[82],stage1_45[107],stage1_44[161],stage1_43[206]}
   );
   gpc606_5 gpc1736 (
      {stage0_44[190], stage0_44[191], stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[59],stage1_46[83],stage1_45[108],stage1_44[162]}
   );
   gpc606_5 gpc1737 (
      {stage0_44[196], stage0_44[197], stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[60],stage1_46[84],stage1_45[109],stage1_44[163]}
   );
   gpc606_5 gpc1738 (
      {stage0_44[202], stage0_44[203], stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[61],stage1_46[85],stage1_45[110],stage1_44[164]}
   );
   gpc606_5 gpc1739 (
      {stage0_44[208], stage0_44[209], stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[62],stage1_46[86],stage1_45[111],stage1_44[165]}
   );
   gpc606_5 gpc1740 (
      {stage0_44[214], stage0_44[215], stage0_44[216], stage0_44[217], stage0_44[218], stage0_44[219]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[63],stage1_46[87],stage1_45[112],stage1_44[166]}
   );
   gpc606_5 gpc1741 (
      {stage0_44[220], stage0_44[221], stage0_44[222], stage0_44[223], stage0_44[224], stage0_44[225]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[64],stage1_46[88],stage1_45[113],stage1_44[167]}
   );
   gpc606_5 gpc1742 (
      {stage0_44[226], stage0_44[227], stage0_44[228], stage0_44[229], stage0_44[230], stage0_44[231]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[65],stage1_46[89],stage1_45[114],stage1_44[168]}
   );
   gpc606_5 gpc1743 (
      {stage0_44[232], stage0_44[233], stage0_44[234], stage0_44[235], stage0_44[236], stage0_44[237]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[66],stage1_46[90],stage1_45[115],stage1_44[169]}
   );
   gpc606_5 gpc1744 (
      {stage0_44[238], stage0_44[239], stage0_44[240], stage0_44[241], stage0_44[242], stage0_44[243]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[67],stage1_46[91],stage1_45[116],stage1_44[170]}
   );
   gpc606_5 gpc1745 (
      {stage0_44[244], stage0_44[245], stage0_44[246], stage0_44[247], stage0_44[248], stage0_44[249]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[68],stage1_46[92],stage1_45[117],stage1_44[171]}
   );
   gpc606_5 gpc1746 (
      {stage0_44[250], stage0_44[251], stage0_44[252], stage0_44[253], stage0_44[254], stage0_44[255]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[69],stage1_46[93],stage1_45[118],stage1_44[172]}
   );
   gpc606_5 gpc1747 (
      {stage0_44[256], stage0_44[257], stage0_44[258], stage0_44[259], stage0_44[260], stage0_44[261]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[70],stage1_46[94],stage1_45[119],stage1_44[173]}
   );
   gpc606_5 gpc1748 (
      {stage0_44[262], stage0_44[263], stage0_44[264], stage0_44[265], stage0_44[266], stage0_44[267]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[71],stage1_46[95],stage1_45[120],stage1_44[174]}
   );
   gpc606_5 gpc1749 (
      {stage0_44[268], stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[72],stage1_46[96],stage1_45[121],stage1_44[175]}
   );
   gpc606_5 gpc1750 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278], stage0_44[279]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[73],stage1_46[97],stage1_45[122],stage1_44[176]}
   );
   gpc606_5 gpc1751 (
      {stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283], stage0_44[284], stage0_44[285]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[74],stage1_46[98],stage1_45[123],stage1_44[177]}
   );
   gpc606_5 gpc1752 (
      {stage0_44[286], stage0_44[287], stage0_44[288], stage0_44[289], stage0_44[290], stage0_44[291]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[75],stage1_46[99],stage1_45[124],stage1_44[178]}
   );
   gpc606_5 gpc1753 (
      {stage0_44[292], stage0_44[293], stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[76],stage1_46[100],stage1_45[125],stage1_44[179]}
   );
   gpc606_5 gpc1754 (
      {stage0_44[298], stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[77],stage1_46[101],stage1_45[126],stage1_44[180]}
   );
   gpc606_5 gpc1755 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308], stage0_44[309]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[78],stage1_46[102],stage1_45[127],stage1_44[181]}
   );
   gpc606_5 gpc1756 (
      {stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313], stage0_44[314], stage0_44[315]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[79],stage1_46[103],stage1_45[128],stage1_44[182]}
   );
   gpc606_5 gpc1757 (
      {stage0_44[316], stage0_44[317], stage0_44[318], stage0_44[319], stage0_44[320], stage0_44[321]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[80],stage1_46[104],stage1_45[129],stage1_44[183]}
   );
   gpc606_5 gpc1758 (
      {stage0_44[322], stage0_44[323], stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[81],stage1_46[105],stage1_45[130],stage1_44[184]}
   );
   gpc606_5 gpc1759 (
      {stage0_44[328], stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[82],stage1_46[106],stage1_45[131],stage1_44[185]}
   );
   gpc606_5 gpc1760 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338], stage0_44[339]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[83],stage1_46[107],stage1_45[132],stage1_44[186]}
   );
   gpc606_5 gpc1761 (
      {stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343], stage0_44[344], stage0_44[345]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[84],stage1_46[108],stage1_45[133],stage1_44[187]}
   );
   gpc606_5 gpc1762 (
      {stage0_44[346], stage0_44[347], stage0_44[348], stage0_44[349], stage0_44[350], stage0_44[351]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[85],stage1_46[109],stage1_45[134],stage1_44[188]}
   );
   gpc606_5 gpc1763 (
      {stage0_44[352], stage0_44[353], stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[86],stage1_46[110],stage1_45[135],stage1_44[189]}
   );
   gpc606_5 gpc1764 (
      {stage0_44[358], stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[87],stage1_46[111],stage1_45[136],stage1_44[190]}
   );
   gpc606_5 gpc1765 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368], stage0_44[369]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[88],stage1_46[112],stage1_45[137],stage1_44[191]}
   );
   gpc606_5 gpc1766 (
      {stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373], stage0_44[374], stage0_44[375]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[89],stage1_46[113],stage1_45[138],stage1_44[192]}
   );
   gpc606_5 gpc1767 (
      {stage0_44[376], stage0_44[377], stage0_44[378], stage0_44[379], stage0_44[380], stage0_44[381]},
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190], stage0_46[191]},
      {stage1_48[31],stage1_47[90],stage1_46[114],stage1_45[139],stage1_44[193]}
   );
   gpc606_5 gpc1768 (
      {stage0_44[382], stage0_44[383], stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387]},
      {stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195], stage0_46[196], stage0_46[197]},
      {stage1_48[32],stage1_47[91],stage1_46[115],stage1_45[140],stage1_44[194]}
   );
   gpc606_5 gpc1769 (
      {stage0_44[388], stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_46[198], stage0_46[199], stage0_46[200], stage0_46[201], stage0_46[202], stage0_46[203]},
      {stage1_48[33],stage1_47[92],stage1_46[116],stage1_45[141],stage1_44[195]}
   );
   gpc606_5 gpc1770 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398], stage0_44[399]},
      {stage0_46[204], stage0_46[205], stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209]},
      {stage1_48[34],stage1_47[93],stage1_46[117],stage1_45[142],stage1_44[196]}
   );
   gpc606_5 gpc1771 (
      {stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403], stage0_44[404], stage0_44[405]},
      {stage0_46[210], stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage1_48[35],stage1_47[94],stage1_46[118],stage1_45[143],stage1_44[197]}
   );
   gpc606_5 gpc1772 (
      {stage0_44[406], stage0_44[407], stage0_44[408], stage0_44[409], stage0_44[410], stage0_44[411]},
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220], stage0_46[221]},
      {stage1_48[36],stage1_47[95],stage1_46[119],stage1_45[144],stage1_44[198]}
   );
   gpc606_5 gpc1773 (
      {stage0_44[412], stage0_44[413], stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417]},
      {stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225], stage0_46[226], stage0_46[227]},
      {stage1_48[37],stage1_47[96],stage1_46[120],stage1_45[145],stage1_44[199]}
   );
   gpc606_5 gpc1774 (
      {stage0_44[418], stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_46[228], stage0_46[229], stage0_46[230], stage0_46[231], stage0_46[232], stage0_46[233]},
      {stage1_48[38],stage1_47[97],stage1_46[121],stage1_45[146],stage1_44[200]}
   );
   gpc606_5 gpc1775 (
      {stage0_44[424], stage0_44[425], stage0_44[426], stage0_44[427], stage0_44[428], stage0_44[429]},
      {stage0_46[234], stage0_46[235], stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239]},
      {stage1_48[39],stage1_47[98],stage1_46[122],stage1_45[147],stage1_44[201]}
   );
   gpc606_5 gpc1776 (
      {stage0_44[430], stage0_44[431], stage0_44[432], stage0_44[433], stage0_44[434], stage0_44[435]},
      {stage0_46[240], stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage1_48[40],stage1_47[99],stage1_46[123],stage1_45[148],stage1_44[202]}
   );
   gpc606_5 gpc1777 (
      {stage0_44[436], stage0_44[437], stage0_44[438], stage0_44[439], stage0_44[440], stage0_44[441]},
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250], stage0_46[251]},
      {stage1_48[41],stage1_47[100],stage1_46[124],stage1_45[149],stage1_44[203]}
   );
   gpc606_5 gpc1778 (
      {stage0_44[442], stage0_44[443], stage0_44[444], stage0_44[445], stage0_44[446], stage0_44[447]},
      {stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255], stage0_46[256], stage0_46[257]},
      {stage1_48[42],stage1_47[101],stage1_46[125],stage1_45[150],stage1_44[204]}
   );
   gpc606_5 gpc1779 (
      {stage0_45[354], stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[43],stage1_47[102],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1780 (
      {stage0_45[360], stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[44],stage1_47[103],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1781 (
      {stage0_45[366], stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[45],stage1_47[104],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1782 (
      {stage0_45[372], stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[46],stage1_47[105],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1783 (
      {stage0_45[378], stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[47],stage1_47[106],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1784 (
      {stage0_45[384], stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[48],stage1_47[107],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1785 (
      {stage0_45[390], stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[49],stage1_47[108],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1786 (
      {stage0_45[396], stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[50],stage1_47[109],stage1_46[133],stage1_45[158]}
   );
   gpc606_5 gpc1787 (
      {stage0_45[402], stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[51],stage1_47[110],stage1_46[134],stage1_45[159]}
   );
   gpc606_5 gpc1788 (
      {stage0_45[408], stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[52],stage1_47[111],stage1_46[135],stage1_45[160]}
   );
   gpc606_5 gpc1789 (
      {stage0_45[414], stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[53],stage1_47[112],stage1_46[136],stage1_45[161]}
   );
   gpc606_5 gpc1790 (
      {stage0_45[420], stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[54],stage1_47[113],stage1_46[137],stage1_45[162]}
   );
   gpc606_5 gpc1791 (
      {stage0_45[426], stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[55],stage1_47[114],stage1_46[138],stage1_45[163]}
   );
   gpc606_5 gpc1792 (
      {stage0_45[432], stage0_45[433], stage0_45[434], stage0_45[435], stage0_45[436], stage0_45[437]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[56],stage1_47[115],stage1_46[139],stage1_45[164]}
   );
   gpc606_5 gpc1793 (
      {stage0_45[438], stage0_45[439], stage0_45[440], stage0_45[441], stage0_45[442], stage0_45[443]},
      {stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage1_49[14],stage1_48[57],stage1_47[116],stage1_46[140],stage1_45[165]}
   );
   gpc606_5 gpc1794 (
      {stage0_45[444], stage0_45[445], stage0_45[446], stage0_45[447], stage0_45[448], stage0_45[449]},
      {stage0_47[90], stage0_47[91], stage0_47[92], stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage1_49[15],stage1_48[58],stage1_47[117],stage1_46[141],stage1_45[166]}
   );
   gpc606_5 gpc1795 (
      {stage0_45[450], stage0_45[451], stage0_45[452], stage0_45[453], stage0_45[454], stage0_45[455]},
      {stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage1_49[16],stage1_48[59],stage1_47[118],stage1_46[142],stage1_45[167]}
   );
   gpc606_5 gpc1796 (
      {stage0_45[456], stage0_45[457], stage0_45[458], stage0_45[459], stage0_45[460], stage0_45[461]},
      {stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage1_49[17],stage1_48[60],stage1_47[119],stage1_46[143],stage1_45[168]}
   );
   gpc606_5 gpc1797 (
      {stage0_45[462], stage0_45[463], stage0_45[464], stage0_45[465], stage0_45[466], stage0_45[467]},
      {stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage1_49[18],stage1_48[61],stage1_47[120],stage1_46[144],stage1_45[169]}
   );
   gpc606_5 gpc1798 (
      {stage0_45[468], stage0_45[469], stage0_45[470], stage0_45[471], stage0_45[472], stage0_45[473]},
      {stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117], stage0_47[118], stage0_47[119]},
      {stage1_49[19],stage1_48[62],stage1_47[121],stage1_46[145],stage1_45[170]}
   );
   gpc606_5 gpc1799 (
      {stage0_45[474], stage0_45[475], stage0_45[476], stage0_45[477], stage0_45[478], stage0_45[479]},
      {stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123], stage0_47[124], stage0_47[125]},
      {stage1_49[20],stage1_48[63],stage1_47[122],stage1_46[146],stage1_45[171]}
   );
   gpc606_5 gpc1800 (
      {stage0_45[480], stage0_45[481], stage0_45[482], stage0_45[483], stage0_45[484], stage0_45[485]},
      {stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129], stage0_47[130], stage0_47[131]},
      {stage1_49[21],stage1_48[64],stage1_47[123],stage1_46[147],stage1_45[172]}
   );
   gpc606_5 gpc1801 (
      {stage0_45[486], stage0_45[487], stage0_45[488], stage0_45[489], stage0_45[490], stage0_45[491]},
      {stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135], stage0_47[136], stage0_47[137]},
      {stage1_49[22],stage1_48[65],stage1_47[124],stage1_46[148],stage1_45[173]}
   );
   gpc606_5 gpc1802 (
      {stage0_45[492], stage0_45[493], stage0_45[494], stage0_45[495], stage0_45[496], stage0_45[497]},
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142], stage0_47[143]},
      {stage1_49[23],stage1_48[66],stage1_47[125],stage1_46[149],stage1_45[174]}
   );
   gpc615_5 gpc1803 (
      {stage0_46[258], stage0_46[259], stage0_46[260], stage0_46[261], stage0_46[262]},
      {stage0_47[144]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[24],stage1_48[67],stage1_47[126],stage1_46[150]}
   );
   gpc615_5 gpc1804 (
      {stage0_46[263], stage0_46[264], stage0_46[265], stage0_46[266], stage0_46[267]},
      {stage0_47[145]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[25],stage1_48[68],stage1_47[127],stage1_46[151]}
   );
   gpc615_5 gpc1805 (
      {stage0_46[268], stage0_46[269], stage0_46[270], stage0_46[271], stage0_46[272]},
      {stage0_47[146]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[26],stage1_48[69],stage1_47[128],stage1_46[152]}
   );
   gpc615_5 gpc1806 (
      {stage0_46[273], stage0_46[274], stage0_46[275], stage0_46[276], stage0_46[277]},
      {stage0_47[147]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[27],stage1_48[70],stage1_47[129],stage1_46[153]}
   );
   gpc615_5 gpc1807 (
      {stage0_46[278], stage0_46[279], stage0_46[280], stage0_46[281], stage0_46[282]},
      {stage0_47[148]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[28],stage1_48[71],stage1_47[130],stage1_46[154]}
   );
   gpc615_5 gpc1808 (
      {stage0_46[283], stage0_46[284], stage0_46[285], stage0_46[286], stage0_46[287]},
      {stage0_47[149]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[29],stage1_48[72],stage1_47[131],stage1_46[155]}
   );
   gpc615_5 gpc1809 (
      {stage0_46[288], stage0_46[289], stage0_46[290], stage0_46[291], stage0_46[292]},
      {stage0_47[150]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[30],stage1_48[73],stage1_47[132],stage1_46[156]}
   );
   gpc615_5 gpc1810 (
      {stage0_46[293], stage0_46[294], stage0_46[295], stage0_46[296], stage0_46[297]},
      {stage0_47[151]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[31],stage1_48[74],stage1_47[133],stage1_46[157]}
   );
   gpc615_5 gpc1811 (
      {stage0_46[298], stage0_46[299], stage0_46[300], stage0_46[301], stage0_46[302]},
      {stage0_47[152]},
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage1_50[8],stage1_49[32],stage1_48[75],stage1_47[134],stage1_46[158]}
   );
   gpc615_5 gpc1812 (
      {stage0_46[303], stage0_46[304], stage0_46[305], stage0_46[306], stage0_46[307]},
      {stage0_47[153]},
      {stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58], stage0_48[59]},
      {stage1_50[9],stage1_49[33],stage1_48[76],stage1_47[135],stage1_46[159]}
   );
   gpc615_5 gpc1813 (
      {stage0_46[308], stage0_46[309], stage0_46[310], stage0_46[311], stage0_46[312]},
      {stage0_47[154]},
      {stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64], stage0_48[65]},
      {stage1_50[10],stage1_49[34],stage1_48[77],stage1_47[136],stage1_46[160]}
   );
   gpc615_5 gpc1814 (
      {stage0_46[313], stage0_46[314], stage0_46[315], stage0_46[316], stage0_46[317]},
      {stage0_47[155]},
      {stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70], stage0_48[71]},
      {stage1_50[11],stage1_49[35],stage1_48[78],stage1_47[137],stage1_46[161]}
   );
   gpc615_5 gpc1815 (
      {stage0_46[318], stage0_46[319], stage0_46[320], stage0_46[321], stage0_46[322]},
      {stage0_47[156]},
      {stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75], stage0_48[76], stage0_48[77]},
      {stage1_50[12],stage1_49[36],stage1_48[79],stage1_47[138],stage1_46[162]}
   );
   gpc615_5 gpc1816 (
      {stage0_46[323], stage0_46[324], stage0_46[325], stage0_46[326], stage0_46[327]},
      {stage0_47[157]},
      {stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81], stage0_48[82], stage0_48[83]},
      {stage1_50[13],stage1_49[37],stage1_48[80],stage1_47[139],stage1_46[163]}
   );
   gpc615_5 gpc1817 (
      {stage0_46[328], stage0_46[329], stage0_46[330], stage0_46[331], stage0_46[332]},
      {stage0_47[158]},
      {stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89]},
      {stage1_50[14],stage1_49[38],stage1_48[81],stage1_47[140],stage1_46[164]}
   );
   gpc615_5 gpc1818 (
      {stage0_46[333], stage0_46[334], stage0_46[335], stage0_46[336], stage0_46[337]},
      {stage0_47[159]},
      {stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage1_50[15],stage1_49[39],stage1_48[82],stage1_47[141],stage1_46[165]}
   );
   gpc615_5 gpc1819 (
      {stage0_46[338], stage0_46[339], stage0_46[340], stage0_46[341], stage0_46[342]},
      {stage0_47[160]},
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100], stage0_48[101]},
      {stage1_50[16],stage1_49[40],stage1_48[83],stage1_47[142],stage1_46[166]}
   );
   gpc615_5 gpc1820 (
      {stage0_46[343], stage0_46[344], stage0_46[345], stage0_46[346], stage0_46[347]},
      {stage0_47[161]},
      {stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105], stage0_48[106], stage0_48[107]},
      {stage1_50[17],stage1_49[41],stage1_48[84],stage1_47[143],stage1_46[167]}
   );
   gpc615_5 gpc1821 (
      {stage0_46[348], stage0_46[349], stage0_46[350], stage0_46[351], stage0_46[352]},
      {stage0_47[162]},
      {stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111], stage0_48[112], stage0_48[113]},
      {stage1_50[18],stage1_49[42],stage1_48[85],stage1_47[144],stage1_46[168]}
   );
   gpc615_5 gpc1822 (
      {stage0_46[353], stage0_46[354], stage0_46[355], stage0_46[356], stage0_46[357]},
      {stage0_47[163]},
      {stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119]},
      {stage1_50[19],stage1_49[43],stage1_48[86],stage1_47[145],stage1_46[169]}
   );
   gpc615_5 gpc1823 (
      {stage0_46[358], stage0_46[359], stage0_46[360], stage0_46[361], stage0_46[362]},
      {stage0_47[164]},
      {stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage1_50[20],stage1_49[44],stage1_48[87],stage1_47[146],stage1_46[170]}
   );
   gpc615_5 gpc1824 (
      {stage0_46[363], stage0_46[364], stage0_46[365], stage0_46[366], stage0_46[367]},
      {stage0_47[165]},
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130], stage0_48[131]},
      {stage1_50[21],stage1_49[45],stage1_48[88],stage1_47[147],stage1_46[171]}
   );
   gpc615_5 gpc1825 (
      {stage0_46[368], stage0_46[369], stage0_46[370], stage0_46[371], stage0_46[372]},
      {stage0_47[166]},
      {stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135], stage0_48[136], stage0_48[137]},
      {stage1_50[22],stage1_49[46],stage1_48[89],stage1_47[148],stage1_46[172]}
   );
   gpc615_5 gpc1826 (
      {stage0_46[373], stage0_46[374], stage0_46[375], stage0_46[376], stage0_46[377]},
      {stage0_47[167]},
      {stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141], stage0_48[142], stage0_48[143]},
      {stage1_50[23],stage1_49[47],stage1_48[90],stage1_47[149],stage1_46[173]}
   );
   gpc615_5 gpc1827 (
      {stage0_46[378], stage0_46[379], stage0_46[380], stage0_46[381], stage0_46[382]},
      {stage0_47[168]},
      {stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149]},
      {stage1_50[24],stage1_49[48],stage1_48[91],stage1_47[150],stage1_46[174]}
   );
   gpc615_5 gpc1828 (
      {stage0_46[383], stage0_46[384], stage0_46[385], stage0_46[386], stage0_46[387]},
      {stage0_47[169]},
      {stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage1_50[25],stage1_49[49],stage1_48[92],stage1_47[151],stage1_46[175]}
   );
   gpc606_5 gpc1829 (
      {stage0_47[170], stage0_47[171], stage0_47[172], stage0_47[173], stage0_47[174], stage0_47[175]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[26],stage1_49[50],stage1_48[93],stage1_47[152]}
   );
   gpc606_5 gpc1830 (
      {stage0_47[176], stage0_47[177], stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[27],stage1_49[51],stage1_48[94],stage1_47[153]}
   );
   gpc606_5 gpc1831 (
      {stage0_47[182], stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[28],stage1_49[52],stage1_48[95],stage1_47[154]}
   );
   gpc606_5 gpc1832 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192], stage0_47[193]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[29],stage1_49[53],stage1_48[96],stage1_47[155]}
   );
   gpc606_5 gpc1833 (
      {stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197], stage0_47[198], stage0_47[199]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[30],stage1_49[54],stage1_48[97],stage1_47[156]}
   );
   gpc606_5 gpc1834 (
      {stage0_47[200], stage0_47[201], stage0_47[202], stage0_47[203], stage0_47[204], stage0_47[205]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[31],stage1_49[55],stage1_48[98],stage1_47[157]}
   );
   gpc606_5 gpc1835 (
      {stage0_47[206], stage0_47[207], stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[32],stage1_49[56],stage1_48[99],stage1_47[158]}
   );
   gpc606_5 gpc1836 (
      {stage0_47[212], stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[33],stage1_49[57],stage1_48[100],stage1_47[159]}
   );
   gpc606_5 gpc1837 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222], stage0_47[223]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[34],stage1_49[58],stage1_48[101],stage1_47[160]}
   );
   gpc606_5 gpc1838 (
      {stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227], stage0_47[228], stage0_47[229]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[35],stage1_49[59],stage1_48[102],stage1_47[161]}
   );
   gpc606_5 gpc1839 (
      {stage0_47[230], stage0_47[231], stage0_47[232], stage0_47[233], stage0_47[234], stage0_47[235]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[36],stage1_49[60],stage1_48[103],stage1_47[162]}
   );
   gpc606_5 gpc1840 (
      {stage0_47[236], stage0_47[237], stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[37],stage1_49[61],stage1_48[104],stage1_47[163]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[242], stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246]},
      {stage0_48[156]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[38],stage1_49[62],stage1_48[105],stage1_47[164]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[247], stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251]},
      {stage0_48[157]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[39],stage1_49[63],stage1_48[106],stage1_47[165]}
   );
   gpc615_5 gpc1843 (
      {stage0_47[252], stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256]},
      {stage0_48[158]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[40],stage1_49[64],stage1_48[107],stage1_47[166]}
   );
   gpc615_5 gpc1844 (
      {stage0_47[257], stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261]},
      {stage0_48[159]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[41],stage1_49[65],stage1_48[108],stage1_47[167]}
   );
   gpc615_5 gpc1845 (
      {stage0_47[262], stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266]},
      {stage0_48[160]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[42],stage1_49[66],stage1_48[109],stage1_47[168]}
   );
   gpc615_5 gpc1846 (
      {stage0_47[267], stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271]},
      {stage0_48[161]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[43],stage1_49[67],stage1_48[110],stage1_47[169]}
   );
   gpc615_5 gpc1847 (
      {stage0_47[272], stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276]},
      {stage0_48[162]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[44],stage1_49[68],stage1_48[111],stage1_47[170]}
   );
   gpc615_5 gpc1848 (
      {stage0_47[277], stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281]},
      {stage0_48[163]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[45],stage1_49[69],stage1_48[112],stage1_47[171]}
   );
   gpc615_5 gpc1849 (
      {stage0_47[282], stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286]},
      {stage0_48[164]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[46],stage1_49[70],stage1_48[113],stage1_47[172]}
   );
   gpc615_5 gpc1850 (
      {stage0_47[287], stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291]},
      {stage0_48[165]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[47],stage1_49[71],stage1_48[114],stage1_47[173]}
   );
   gpc615_5 gpc1851 (
      {stage0_47[292], stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296]},
      {stage0_48[166]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[48],stage1_49[72],stage1_48[115],stage1_47[174]}
   );
   gpc615_5 gpc1852 (
      {stage0_47[297], stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301]},
      {stage0_48[167]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[49],stage1_49[73],stage1_48[116],stage1_47[175]}
   );
   gpc615_5 gpc1853 (
      {stage0_47[302], stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306]},
      {stage0_48[168]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[50],stage1_49[74],stage1_48[117],stage1_47[176]}
   );
   gpc615_5 gpc1854 (
      {stage0_47[307], stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311]},
      {stage0_48[169]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[51],stage1_49[75],stage1_48[118],stage1_47[177]}
   );
   gpc615_5 gpc1855 (
      {stage0_47[312], stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316]},
      {stage0_48[170]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[52],stage1_49[76],stage1_48[119],stage1_47[178]}
   );
   gpc615_5 gpc1856 (
      {stage0_47[317], stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321]},
      {stage0_48[171]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[53],stage1_49[77],stage1_48[120],stage1_47[179]}
   );
   gpc615_5 gpc1857 (
      {stage0_47[322], stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326]},
      {stage0_48[172]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[54],stage1_49[78],stage1_48[121],stage1_47[180]}
   );
   gpc615_5 gpc1858 (
      {stage0_47[327], stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331]},
      {stage0_48[173]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[55],stage1_49[79],stage1_48[122],stage1_47[181]}
   );
   gpc615_5 gpc1859 (
      {stage0_47[332], stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336]},
      {stage0_48[174]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[56],stage1_49[80],stage1_48[123],stage1_47[182]}
   );
   gpc615_5 gpc1860 (
      {stage0_47[337], stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341]},
      {stage0_48[175]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[57],stage1_49[81],stage1_48[124],stage1_47[183]}
   );
   gpc615_5 gpc1861 (
      {stage0_47[342], stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346]},
      {stage0_48[176]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[58],stage1_49[82],stage1_48[125],stage1_47[184]}
   );
   gpc615_5 gpc1862 (
      {stage0_47[347], stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351]},
      {stage0_48[177]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[59],stage1_49[83],stage1_48[126],stage1_47[185]}
   );
   gpc615_5 gpc1863 (
      {stage0_47[352], stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356]},
      {stage0_48[178]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[60],stage1_49[84],stage1_48[127],stage1_47[186]}
   );
   gpc615_5 gpc1864 (
      {stage0_47[357], stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361]},
      {stage0_48[179]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[61],stage1_49[85],stage1_48[128],stage1_47[187]}
   );
   gpc615_5 gpc1865 (
      {stage0_47[362], stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366]},
      {stage0_48[180]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[62],stage1_49[86],stage1_48[129],stage1_47[188]}
   );
   gpc615_5 gpc1866 (
      {stage0_47[367], stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371]},
      {stage0_48[181]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[63],stage1_49[87],stage1_48[130],stage1_47[189]}
   );
   gpc615_5 gpc1867 (
      {stage0_47[372], stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376]},
      {stage0_48[182]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[64],stage1_49[88],stage1_48[131],stage1_47[190]}
   );
   gpc615_5 gpc1868 (
      {stage0_47[377], stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381]},
      {stage0_48[183]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[65],stage1_49[89],stage1_48[132],stage1_47[191]}
   );
   gpc615_5 gpc1869 (
      {stage0_47[382], stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386]},
      {stage0_48[184]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[66],stage1_49[90],stage1_48[133],stage1_47[192]}
   );
   gpc615_5 gpc1870 (
      {stage0_47[387], stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391]},
      {stage0_48[185]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[67],stage1_49[91],stage1_48[134],stage1_47[193]}
   );
   gpc615_5 gpc1871 (
      {stage0_47[392], stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396]},
      {stage0_48[186]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[68],stage1_49[92],stage1_48[135],stage1_47[194]}
   );
   gpc615_5 gpc1872 (
      {stage0_47[397], stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401]},
      {stage0_48[187]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[69],stage1_49[93],stage1_48[136],stage1_47[195]}
   );
   gpc615_5 gpc1873 (
      {stage0_47[402], stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406]},
      {stage0_48[188]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[70],stage1_49[94],stage1_48[137],stage1_47[196]}
   );
   gpc615_5 gpc1874 (
      {stage0_47[407], stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411]},
      {stage0_48[189]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[71],stage1_49[95],stage1_48[138],stage1_47[197]}
   );
   gpc615_5 gpc1875 (
      {stage0_47[412], stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416]},
      {stage0_48[190]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[72],stage1_49[96],stage1_48[139],stage1_47[198]}
   );
   gpc615_5 gpc1876 (
      {stage0_47[417], stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421]},
      {stage0_48[191]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[73],stage1_49[97],stage1_48[140],stage1_47[199]}
   );
   gpc615_5 gpc1877 (
      {stage0_47[422], stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426]},
      {stage0_48[192]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[74],stage1_49[98],stage1_48[141],stage1_47[200]}
   );
   gpc615_5 gpc1878 (
      {stage0_47[427], stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431]},
      {stage0_48[193]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[75],stage1_49[99],stage1_48[142],stage1_47[201]}
   );
   gpc615_5 gpc1879 (
      {stage0_47[432], stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436]},
      {stage0_48[194]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[76],stage1_49[100],stage1_48[143],stage1_47[202]}
   );
   gpc606_5 gpc1880 (
      {stage0_48[195], stage0_48[196], stage0_48[197], stage0_48[198], stage0_48[199], stage0_48[200]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[51],stage1_50[77],stage1_49[101],stage1_48[144]}
   );
   gpc606_5 gpc1881 (
      {stage0_48[201], stage0_48[202], stage0_48[203], stage0_48[204], stage0_48[205], stage0_48[206]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[52],stage1_50[78],stage1_49[102],stage1_48[145]}
   );
   gpc606_5 gpc1882 (
      {stage0_48[207], stage0_48[208], stage0_48[209], stage0_48[210], stage0_48[211], stage0_48[212]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[53],stage1_50[79],stage1_49[103],stage1_48[146]}
   );
   gpc606_5 gpc1883 (
      {stage0_48[213], stage0_48[214], stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[54],stage1_50[80],stage1_49[104],stage1_48[147]}
   );
   gpc606_5 gpc1884 (
      {stage0_48[219], stage0_48[220], stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[55],stage1_50[81],stage1_49[105],stage1_48[148]}
   );
   gpc606_5 gpc1885 (
      {stage0_48[225], stage0_48[226], stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[56],stage1_50[82],stage1_49[106],stage1_48[149]}
   );
   gpc606_5 gpc1886 (
      {stage0_48[231], stage0_48[232], stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[57],stage1_50[83],stage1_49[107],stage1_48[150]}
   );
   gpc606_5 gpc1887 (
      {stage0_48[237], stage0_48[238], stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[58],stage1_50[84],stage1_49[108],stage1_48[151]}
   );
   gpc606_5 gpc1888 (
      {stage0_48[243], stage0_48[244], stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[59],stage1_50[85],stage1_49[109],stage1_48[152]}
   );
   gpc606_5 gpc1889 (
      {stage0_48[249], stage0_48[250], stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[60],stage1_50[86],stage1_49[110],stage1_48[153]}
   );
   gpc606_5 gpc1890 (
      {stage0_48[255], stage0_48[256], stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[61],stage1_50[87],stage1_49[111],stage1_48[154]}
   );
   gpc606_5 gpc1891 (
      {stage0_48[261], stage0_48[262], stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[62],stage1_50[88],stage1_49[112],stage1_48[155]}
   );
   gpc606_5 gpc1892 (
      {stage0_48[267], stage0_48[268], stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[63],stage1_50[89],stage1_49[113],stage1_48[156]}
   );
   gpc606_5 gpc1893 (
      {stage0_48[273], stage0_48[274], stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[64],stage1_50[90],stage1_49[114],stage1_48[157]}
   );
   gpc606_5 gpc1894 (
      {stage0_48[279], stage0_48[280], stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[65],stage1_50[91],stage1_49[115],stage1_48[158]}
   );
   gpc606_5 gpc1895 (
      {stage0_48[285], stage0_48[286], stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[66],stage1_50[92],stage1_49[116],stage1_48[159]}
   );
   gpc606_5 gpc1896 (
      {stage0_48[291], stage0_48[292], stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[67],stage1_50[93],stage1_49[117],stage1_48[160]}
   );
   gpc606_5 gpc1897 (
      {stage0_48[297], stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[68],stage1_50[94],stage1_49[118],stage1_48[161]}
   );
   gpc606_5 gpc1898 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307], stage0_48[308]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[69],stage1_50[95],stage1_49[119],stage1_48[162]}
   );
   gpc606_5 gpc1899 (
      {stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312], stage0_48[313], stage0_48[314]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[70],stage1_50[96],stage1_49[120],stage1_48[163]}
   );
   gpc606_5 gpc1900 (
      {stage0_48[315], stage0_48[316], stage0_48[317], stage0_48[318], stage0_48[319], stage0_48[320]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[71],stage1_50[97],stage1_49[121],stage1_48[164]}
   );
   gpc606_5 gpc1901 (
      {stage0_48[321], stage0_48[322], stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[72],stage1_50[98],stage1_49[122],stage1_48[165]}
   );
   gpc606_5 gpc1902 (
      {stage0_48[327], stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[73],stage1_50[99],stage1_49[123],stage1_48[166]}
   );
   gpc606_5 gpc1903 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337], stage0_48[338]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[74],stage1_50[100],stage1_49[124],stage1_48[167]}
   );
   gpc606_5 gpc1904 (
      {stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342], stage0_48[343], stage0_48[344]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[75],stage1_50[101],stage1_49[125],stage1_48[168]}
   );
   gpc606_5 gpc1905 (
      {stage0_48[345], stage0_48[346], stage0_48[347], stage0_48[348], stage0_48[349], stage0_48[350]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[76],stage1_50[102],stage1_49[126],stage1_48[169]}
   );
   gpc606_5 gpc1906 (
      {stage0_48[351], stage0_48[352], stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[77],stage1_50[103],stage1_49[127],stage1_48[170]}
   );
   gpc606_5 gpc1907 (
      {stage0_48[357], stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[78],stage1_50[104],stage1_49[128],stage1_48[171]}
   );
   gpc606_5 gpc1908 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367], stage0_48[368]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[79],stage1_50[105],stage1_49[129],stage1_48[172]}
   );
   gpc606_5 gpc1909 (
      {stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372], stage0_48[373], stage0_48[374]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[80],stage1_50[106],stage1_49[130],stage1_48[173]}
   );
   gpc606_5 gpc1910 (
      {stage0_48[375], stage0_48[376], stage0_48[377], stage0_48[378], stage0_48[379], stage0_48[380]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[81],stage1_50[107],stage1_49[131],stage1_48[174]}
   );
   gpc606_5 gpc1911 (
      {stage0_48[381], stage0_48[382], stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[82],stage1_50[108],stage1_49[132],stage1_48[175]}
   );
   gpc606_5 gpc1912 (
      {stage0_48[387], stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[83],stage1_50[109],stage1_49[133],stage1_48[176]}
   );
   gpc606_5 gpc1913 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397], stage0_48[398]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[84],stage1_50[110],stage1_49[134],stage1_48[177]}
   );
   gpc606_5 gpc1914 (
      {stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402], stage0_48[403], stage0_48[404]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[85],stage1_50[111],stage1_49[135],stage1_48[178]}
   );
   gpc606_5 gpc1915 (
      {stage0_48[405], stage0_48[406], stage0_48[407], stage0_48[408], stage0_48[409], stage0_48[410]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[86],stage1_50[112],stage1_49[136],stage1_48[179]}
   );
   gpc606_5 gpc1916 (
      {stage0_48[411], stage0_48[412], stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[87],stage1_50[113],stage1_49[137],stage1_48[180]}
   );
   gpc606_5 gpc1917 (
      {stage0_48[417], stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[88],stage1_50[114],stage1_49[138],stage1_48[181]}
   );
   gpc606_5 gpc1918 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427], stage0_48[428]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[89],stage1_50[115],stage1_49[139],stage1_48[182]}
   );
   gpc606_5 gpc1919 (
      {stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432], stage0_48[433], stage0_48[434]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[90],stage1_50[116],stage1_49[140],stage1_48[183]}
   );
   gpc606_5 gpc1920 (
      {stage0_48[435], stage0_48[436], stage0_48[437], stage0_48[438], stage0_48[439], stage0_48[440]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[91],stage1_50[117],stage1_49[141],stage1_48[184]}
   );
   gpc606_5 gpc1921 (
      {stage0_48[441], stage0_48[442], stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[92],stage1_50[118],stage1_49[142],stage1_48[185]}
   );
   gpc606_5 gpc1922 (
      {stage0_48[447], stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[93],stage1_50[119],stage1_49[143],stage1_48[186]}
   );
   gpc606_5 gpc1923 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457], stage0_48[458]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[94],stage1_50[120],stage1_49[144],stage1_48[187]}
   );
   gpc606_5 gpc1924 (
      {stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462], stage0_48[463], stage0_48[464]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[95],stage1_50[121],stage1_49[145],stage1_48[188]}
   );
   gpc606_5 gpc1925 (
      {stage0_48[465], stage0_48[466], stage0_48[467], stage0_48[468], stage0_48[469], stage0_48[470]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[96],stage1_50[122],stage1_49[146],stage1_48[189]}
   );
   gpc606_5 gpc1926 (
      {stage0_48[471], stage0_48[472], stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[97],stage1_50[123],stage1_49[147],stage1_48[190]}
   );
   gpc606_5 gpc1927 (
      {stage0_48[477], stage0_48[478], stage0_48[479], stage0_48[480], stage0_48[481], stage0_48[482]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[98],stage1_50[124],stage1_49[148],stage1_48[191]}
   );
   gpc606_5 gpc1928 (
      {stage0_48[483], stage0_48[484], stage0_48[485], stage0_48[486], stage0_48[487], stage0_48[488]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[99],stage1_50[125],stage1_49[149],stage1_48[192]}
   );
   gpc606_5 gpc1929 (
      {stage0_48[489], stage0_48[490], stage0_48[491], stage0_48[492], stage0_48[493], stage0_48[494]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[100],stage1_50[126],stage1_49[150],stage1_48[193]}
   );
   gpc606_5 gpc1930 (
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[101],stage1_50[127],stage1_49[151]}
   );
   gpc606_5 gpc1931 (
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[102],stage1_50[128],stage1_49[152]}
   );
   gpc606_5 gpc1932 (
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[103],stage1_50[129],stage1_49[153]}
   );
   gpc606_5 gpc1933 (
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[104],stage1_50[130],stage1_49[154]}
   );
   gpc606_5 gpc1934 (
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[105],stage1_50[131],stage1_49[155]}
   );
   gpc606_5 gpc1935 (
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[106],stage1_50[132],stage1_49[156]}
   );
   gpc606_5 gpc1936 (
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[107],stage1_50[133],stage1_49[157]}
   );
   gpc606_5 gpc1937 (
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[108],stage1_50[134],stage1_49[158]}
   );
   gpc606_5 gpc1938 (
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[109],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1939 (
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[110],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1940 (
      {stage0_49[366], stage0_49[367], stage0_49[368], stage0_49[369], stage0_49[370], stage0_49[371]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[111],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1941 (
      {stage0_49[372], stage0_49[373], stage0_49[374], stage0_49[375], stage0_49[376], stage0_49[377]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[112],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1942 (
      {stage0_49[378], stage0_49[379], stage0_49[380], stage0_49[381], stage0_49[382], stage0_49[383]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[113],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1943 (
      {stage0_49[384], stage0_49[385], stage0_49[386], stage0_49[387], stage0_49[388], stage0_49[389]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[114],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1944 (
      {stage0_49[390], stage0_49[391], stage0_49[392], stage0_49[393], stage0_49[394], stage0_49[395]},
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage1_53[14],stage1_52[64],stage1_51[115],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1945 (
      {stage0_49[396], stage0_49[397], stage0_49[398], stage0_49[399], stage0_49[400], stage0_49[401]},
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage1_53[15],stage1_52[65],stage1_51[116],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1946 (
      {stage0_49[402], stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407]},
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage1_53[16],stage1_52[66],stage1_51[117],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1947 (
      {stage0_49[408], stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413]},
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage1_53[17],stage1_52[67],stage1_51[118],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1948 (
      {stage0_49[414], stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419]},
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage1_53[18],stage1_52[68],stage1_51[119],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1949 (
      {stage0_49[420], stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425]},
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage1_53[19],stage1_52[69],stage1_51[120],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1950 (
      {stage0_49[426], stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431]},
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage1_53[20],stage1_52[70],stage1_51[121],stage1_50[147],stage1_49[171]}
   );
   gpc606_5 gpc1951 (
      {stage0_49[432], stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437]},
      {stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129], stage0_51[130], stage0_51[131]},
      {stage1_53[21],stage1_52[71],stage1_51[122],stage1_50[148],stage1_49[172]}
   );
   gpc606_5 gpc1952 (
      {stage0_49[438], stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443]},
      {stage0_51[132], stage0_51[133], stage0_51[134], stage0_51[135], stage0_51[136], stage0_51[137]},
      {stage1_53[22],stage1_52[72],stage1_51[123],stage1_50[149],stage1_49[173]}
   );
   gpc606_5 gpc1953 (
      {stage0_50[300], stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[23],stage1_52[73],stage1_51[124],stage1_50[150]}
   );
   gpc606_5 gpc1954 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310], stage0_50[311]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[24],stage1_52[74],stage1_51[125],stage1_50[151]}
   );
   gpc606_5 gpc1955 (
      {stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315], stage0_50[316], stage0_50[317]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[25],stage1_52[75],stage1_51[126],stage1_50[152]}
   );
   gpc606_5 gpc1956 (
      {stage0_50[318], stage0_50[319], stage0_50[320], stage0_50[321], stage0_50[322], stage0_50[323]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[26],stage1_52[76],stage1_51[127],stage1_50[153]}
   );
   gpc606_5 gpc1957 (
      {stage0_50[324], stage0_50[325], stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[27],stage1_52[77],stage1_51[128],stage1_50[154]}
   );
   gpc606_5 gpc1958 (
      {stage0_50[330], stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[28],stage1_52[78],stage1_51[129],stage1_50[155]}
   );
   gpc606_5 gpc1959 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340], stage0_50[341]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[29],stage1_52[79],stage1_51[130],stage1_50[156]}
   );
   gpc606_5 gpc1960 (
      {stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345], stage0_50[346], stage0_50[347]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[30],stage1_52[80],stage1_51[131],stage1_50[157]}
   );
   gpc606_5 gpc1961 (
      {stage0_50[348], stage0_50[349], stage0_50[350], stage0_50[351], stage0_50[352], stage0_50[353]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[31],stage1_52[81],stage1_51[132],stage1_50[158]}
   );
   gpc606_5 gpc1962 (
      {stage0_50[354], stage0_50[355], stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[32],stage1_52[82],stage1_51[133],stage1_50[159]}
   );
   gpc606_5 gpc1963 (
      {stage0_50[360], stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[33],stage1_52[83],stage1_51[134],stage1_50[160]}
   );
   gpc606_5 gpc1964 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370], stage0_50[371]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[34],stage1_52[84],stage1_51[135],stage1_50[161]}
   );
   gpc606_5 gpc1965 (
      {stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375], stage0_50[376], stage0_50[377]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[35],stage1_52[85],stage1_51[136],stage1_50[162]}
   );
   gpc606_5 gpc1966 (
      {stage0_50[378], stage0_50[379], stage0_50[380], stage0_50[381], stage0_50[382], stage0_50[383]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[36],stage1_52[86],stage1_51[137],stage1_50[163]}
   );
   gpc606_5 gpc1967 (
      {stage0_50[384], stage0_50[385], stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[37],stage1_52[87],stage1_51[138],stage1_50[164]}
   );
   gpc606_5 gpc1968 (
      {stage0_50[390], stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[38],stage1_52[88],stage1_51[139],stage1_50[165]}
   );
   gpc606_5 gpc1969 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400], stage0_50[401]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[39],stage1_52[89],stage1_51[140],stage1_50[166]}
   );
   gpc606_5 gpc1970 (
      {stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405], stage0_50[406], stage0_50[407]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[40],stage1_52[90],stage1_51[141],stage1_50[167]}
   );
   gpc606_5 gpc1971 (
      {stage0_50[408], stage0_50[409], stage0_50[410], stage0_50[411], stage0_50[412], stage0_50[413]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[41],stage1_52[91],stage1_51[142],stage1_50[168]}
   );
   gpc606_5 gpc1972 (
      {stage0_50[414], stage0_50[415], stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[42],stage1_52[92],stage1_51[143],stage1_50[169]}
   );
   gpc606_5 gpc1973 (
      {stage0_50[420], stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[43],stage1_52[93],stage1_51[144],stage1_50[170]}
   );
   gpc606_5 gpc1974 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430], stage0_50[431]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[44],stage1_52[94],stage1_51[145],stage1_50[171]}
   );
   gpc606_5 gpc1975 (
      {stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435], stage0_50[436], stage0_50[437]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[45],stage1_52[95],stage1_51[146],stage1_50[172]}
   );
   gpc606_5 gpc1976 (
      {stage0_50[438], stage0_50[439], stage0_50[440], stage0_50[441], stage0_50[442], stage0_50[443]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[46],stage1_52[96],stage1_51[147],stage1_50[173]}
   );
   gpc606_5 gpc1977 (
      {stage0_50[444], stage0_50[445], stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[47],stage1_52[97],stage1_51[148],stage1_50[174]}
   );
   gpc606_5 gpc1978 (
      {stage0_50[450], stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[48],stage1_52[98],stage1_51[149],stage1_50[175]}
   );
   gpc606_5 gpc1979 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460], stage0_50[461]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[49],stage1_52[99],stage1_51[150],stage1_50[176]}
   );
   gpc606_5 gpc1980 (
      {stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465], stage0_50[466], stage0_50[467]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[50],stage1_52[100],stage1_51[151],stage1_50[177]}
   );
   gpc606_5 gpc1981 (
      {stage0_50[468], stage0_50[469], stage0_50[470], stage0_50[471], stage0_50[472], stage0_50[473]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[51],stage1_52[101],stage1_51[152],stage1_50[178]}
   );
   gpc606_5 gpc1982 (
      {stage0_51[138], stage0_51[139], stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[29],stage1_53[52],stage1_52[102],stage1_51[153]}
   );
   gpc606_5 gpc1983 (
      {stage0_51[144], stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[30],stage1_53[53],stage1_52[103],stage1_51[154]}
   );
   gpc606_5 gpc1984 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154], stage0_51[155]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[31],stage1_53[54],stage1_52[104],stage1_51[155]}
   );
   gpc606_5 gpc1985 (
      {stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159], stage0_51[160], stage0_51[161]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[32],stage1_53[55],stage1_52[105],stage1_51[156]}
   );
   gpc606_5 gpc1986 (
      {stage0_51[162], stage0_51[163], stage0_51[164], stage0_51[165], stage0_51[166], stage0_51[167]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[33],stage1_53[56],stage1_52[106],stage1_51[157]}
   );
   gpc606_5 gpc1987 (
      {stage0_51[168], stage0_51[169], stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[34],stage1_53[57],stage1_52[107],stage1_51[158]}
   );
   gpc606_5 gpc1988 (
      {stage0_51[174], stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[35],stage1_53[58],stage1_52[108],stage1_51[159]}
   );
   gpc606_5 gpc1989 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184], stage0_51[185]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[36],stage1_53[59],stage1_52[109],stage1_51[160]}
   );
   gpc606_5 gpc1990 (
      {stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189], stage0_51[190], stage0_51[191]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[37],stage1_53[60],stage1_52[110],stage1_51[161]}
   );
   gpc606_5 gpc1991 (
      {stage0_51[192], stage0_51[193], stage0_51[194], stage0_51[195], stage0_51[196], stage0_51[197]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[38],stage1_53[61],stage1_52[111],stage1_51[162]}
   );
   gpc606_5 gpc1992 (
      {stage0_51[198], stage0_51[199], stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[39],stage1_53[62],stage1_52[112],stage1_51[163]}
   );
   gpc606_5 gpc1993 (
      {stage0_51[204], stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[40],stage1_53[63],stage1_52[113],stage1_51[164]}
   );
   gpc606_5 gpc1994 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214], stage0_51[215]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[41],stage1_53[64],stage1_52[114],stage1_51[165]}
   );
   gpc606_5 gpc1995 (
      {stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219], stage0_51[220], stage0_51[221]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[42],stage1_53[65],stage1_52[115],stage1_51[166]}
   );
   gpc606_5 gpc1996 (
      {stage0_51[222], stage0_51[223], stage0_51[224], stage0_51[225], stage0_51[226], stage0_51[227]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[43],stage1_53[66],stage1_52[116],stage1_51[167]}
   );
   gpc606_5 gpc1997 (
      {stage0_51[228], stage0_51[229], stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[44],stage1_53[67],stage1_52[117],stage1_51[168]}
   );
   gpc606_5 gpc1998 (
      {stage0_51[234], stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[45],stage1_53[68],stage1_52[118],stage1_51[169]}
   );
   gpc606_5 gpc1999 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244], stage0_51[245]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[46],stage1_53[69],stage1_52[119],stage1_51[170]}
   );
   gpc606_5 gpc2000 (
      {stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249], stage0_51[250], stage0_51[251]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[47],stage1_53[70],stage1_52[120],stage1_51[171]}
   );
   gpc606_5 gpc2001 (
      {stage0_51[252], stage0_51[253], stage0_51[254], stage0_51[255], stage0_51[256], stage0_51[257]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[48],stage1_53[71],stage1_52[121],stage1_51[172]}
   );
   gpc606_5 gpc2002 (
      {stage0_51[258], stage0_51[259], stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[49],stage1_53[72],stage1_52[122],stage1_51[173]}
   );
   gpc606_5 gpc2003 (
      {stage0_51[264], stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[50],stage1_53[73],stage1_52[123],stage1_51[174]}
   );
   gpc606_5 gpc2004 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274], stage0_51[275]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[51],stage1_53[74],stage1_52[124],stage1_51[175]}
   );
   gpc606_5 gpc2005 (
      {stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279], stage0_51[280], stage0_51[281]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[52],stage1_53[75],stage1_52[125],stage1_51[176]}
   );
   gpc606_5 gpc2006 (
      {stage0_51[282], stage0_51[283], stage0_51[284], stage0_51[285], stage0_51[286], stage0_51[287]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[53],stage1_53[76],stage1_52[126],stage1_51[177]}
   );
   gpc606_5 gpc2007 (
      {stage0_51[288], stage0_51[289], stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[54],stage1_53[77],stage1_52[127],stage1_51[178]}
   );
   gpc606_5 gpc2008 (
      {stage0_51[294], stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[55],stage1_53[78],stage1_52[128],stage1_51[179]}
   );
   gpc606_5 gpc2009 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304], stage0_51[305]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[56],stage1_53[79],stage1_52[129],stage1_51[180]}
   );
   gpc606_5 gpc2010 (
      {stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309], stage0_51[310], stage0_51[311]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[57],stage1_53[80],stage1_52[130],stage1_51[181]}
   );
   gpc606_5 gpc2011 (
      {stage0_51[312], stage0_51[313], stage0_51[314], stage0_51[315], stage0_51[316], stage0_51[317]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[58],stage1_53[81],stage1_52[131],stage1_51[182]}
   );
   gpc606_5 gpc2012 (
      {stage0_51[318], stage0_51[319], stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[59],stage1_53[82],stage1_52[132],stage1_51[183]}
   );
   gpc606_5 gpc2013 (
      {stage0_51[324], stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[60],stage1_53[83],stage1_52[133],stage1_51[184]}
   );
   gpc606_5 gpc2014 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334], stage0_51[335]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[61],stage1_53[84],stage1_52[134],stage1_51[185]}
   );
   gpc606_5 gpc2015 (
      {stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339], stage0_51[340], stage0_51[341]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[62],stage1_53[85],stage1_52[135],stage1_51[186]}
   );
   gpc606_5 gpc2016 (
      {stage0_51[342], stage0_51[343], stage0_51[344], stage0_51[345], stage0_51[346], stage0_51[347]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[63],stage1_53[86],stage1_52[136],stage1_51[187]}
   );
   gpc606_5 gpc2017 (
      {stage0_51[348], stage0_51[349], stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[64],stage1_53[87],stage1_52[137],stage1_51[188]}
   );
   gpc606_5 gpc2018 (
      {stage0_51[354], stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[65],stage1_53[88],stage1_52[138],stage1_51[189]}
   );
   gpc606_5 gpc2019 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364], stage0_51[365]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[66],stage1_53[89],stage1_52[139],stage1_51[190]}
   );
   gpc606_5 gpc2020 (
      {stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369], stage0_51[370], stage0_51[371]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[67],stage1_53[90],stage1_52[140],stage1_51[191]}
   );
   gpc606_5 gpc2021 (
      {stage0_51[372], stage0_51[373], stage0_51[374], stage0_51[375], stage0_51[376], stage0_51[377]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[68],stage1_53[91],stage1_52[141],stage1_51[192]}
   );
   gpc606_5 gpc2022 (
      {stage0_51[378], stage0_51[379], stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[69],stage1_53[92],stage1_52[142],stage1_51[193]}
   );
   gpc606_5 gpc2023 (
      {stage0_51[384], stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[70],stage1_53[93],stage1_52[143],stage1_51[194]}
   );
   gpc606_5 gpc2024 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394], stage0_51[395]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[71],stage1_53[94],stage1_52[144],stage1_51[195]}
   );
   gpc606_5 gpc2025 (
      {stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399], stage0_51[400], stage0_51[401]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[72],stage1_53[95],stage1_52[145],stage1_51[196]}
   );
   gpc606_5 gpc2026 (
      {stage0_51[402], stage0_51[403], stage0_51[404], stage0_51[405], stage0_51[406], stage0_51[407]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[73],stage1_53[96],stage1_52[146],stage1_51[197]}
   );
   gpc606_5 gpc2027 (
      {stage0_51[408], stage0_51[409], stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[74],stage1_53[97],stage1_52[147],stage1_51[198]}
   );
   gpc606_5 gpc2028 (
      {stage0_51[414], stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[75],stage1_53[98],stage1_52[148],stage1_51[199]}
   );
   gpc606_5 gpc2029 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424], stage0_51[425]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[76],stage1_53[99],stage1_52[149],stage1_51[200]}
   );
   gpc606_5 gpc2030 (
      {stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429], stage0_51[430], stage0_51[431]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[77],stage1_53[100],stage1_52[150],stage1_51[201]}
   );
   gpc606_5 gpc2031 (
      {stage0_51[432], stage0_51[433], stage0_51[434], stage0_51[435], stage0_51[436], stage0_51[437]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[78],stage1_53[101],stage1_52[151],stage1_51[202]}
   );
   gpc615_5 gpc2032 (
      {stage0_51[438], stage0_51[439], stage0_51[440], stage0_51[441], stage0_51[442]},
      {stage0_52[174]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[79],stage1_53[102],stage1_52[152],stage1_51[203]}
   );
   gpc615_5 gpc2033 (
      {stage0_51[443], stage0_51[444], stage0_51[445], stage0_51[446], stage0_51[447]},
      {stage0_52[175]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[80],stage1_53[103],stage1_52[153],stage1_51[204]}
   );
   gpc615_5 gpc2034 (
      {stage0_51[448], stage0_51[449], stage0_51[450], stage0_51[451], stage0_51[452]},
      {stage0_52[176]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[81],stage1_53[104],stage1_52[154],stage1_51[205]}
   );
   gpc615_5 gpc2035 (
      {stage0_51[453], stage0_51[454], stage0_51[455], stage0_51[456], stage0_51[457]},
      {stage0_52[177]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[82],stage1_53[105],stage1_52[155],stage1_51[206]}
   );
   gpc615_5 gpc2036 (
      {stage0_51[458], stage0_51[459], stage0_51[460], stage0_51[461], stage0_51[462]},
      {stage0_52[178]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[83],stage1_53[106],stage1_52[156],stage1_51[207]}
   );
   gpc615_5 gpc2037 (
      {stage0_51[463], stage0_51[464], stage0_51[465], stage0_51[466], stage0_51[467]},
      {stage0_52[179]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[84],stage1_53[107],stage1_52[157],stage1_51[208]}
   );
   gpc615_5 gpc2038 (
      {stage0_51[468], stage0_51[469], stage0_51[470], stage0_51[471], stage0_51[472]},
      {stage0_52[180]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[85],stage1_53[108],stage1_52[158],stage1_51[209]}
   );
   gpc615_5 gpc2039 (
      {stage0_51[473], stage0_51[474], stage0_51[475], stage0_51[476], stage0_51[477]},
      {stage0_52[181]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[86],stage1_53[109],stage1_52[159],stage1_51[210]}
   );
   gpc615_5 gpc2040 (
      {stage0_51[478], stage0_51[479], stage0_51[480], stage0_51[481], stage0_51[482]},
      {stage0_52[182]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[87],stage1_53[110],stage1_52[160],stage1_51[211]}
   );
   gpc615_5 gpc2041 (
      {stage0_51[483], stage0_51[484], stage0_51[485], stage0_51[486], stage0_51[487]},
      {stage0_52[183]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[88],stage1_53[111],stage1_52[161],stage1_51[212]}
   );
   gpc615_5 gpc2042 (
      {stage0_51[488], stage0_51[489], stage0_51[490], stage0_51[491], stage0_51[492]},
      {stage0_52[184]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[89],stage1_53[112],stage1_52[162],stage1_51[213]}
   );
   gpc615_5 gpc2043 (
      {stage0_51[493], stage0_51[494], stage0_51[495], stage0_51[496], stage0_51[497]},
      {stage0_52[185]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[90],stage1_53[113],stage1_52[163],stage1_51[214]}
   );
   gpc623_5 gpc2044 (
      {stage0_51[498], stage0_51[499], stage0_51[500]},
      {stage0_52[186], stage0_52[187]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[91],stage1_53[114],stage1_52[164],stage1_51[215]}
   );
   gpc606_5 gpc2045 (
      {stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191], stage0_52[192], stage0_52[193]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[92],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2046 (
      {stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197], stage0_52[198], stage0_52[199]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[93],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2047 (
      {stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203], stage0_52[204], stage0_52[205]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[94],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2048 (
      {stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209], stage0_52[210], stage0_52[211]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[95],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2049 (
      {stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215], stage0_52[216], stage0_52[217]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[96],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2050 (
      {stage0_52[218], stage0_52[219], stage0_52[220], stage0_52[221], stage0_52[222], stage0_52[223]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[97],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2051 (
      {stage0_52[224], stage0_52[225], stage0_52[226], stage0_52[227], stage0_52[228], stage0_52[229]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[98],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2052 (
      {stage0_52[230], stage0_52[231], stage0_52[232], stage0_52[233], stage0_52[234], stage0_52[235]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[99],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2053 (
      {stage0_52[236], stage0_52[237], stage0_52[238], stage0_52[239], stage0_52[240], stage0_52[241]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[100],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2054 (
      {stage0_52[242], stage0_52[243], stage0_52[244], stage0_52[245], stage0_52[246], stage0_52[247]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[101],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2055 (
      {stage0_52[248], stage0_52[249], stage0_52[250], stage0_52[251], stage0_52[252], stage0_52[253]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[102],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2056 (
      {stage0_52[254], stage0_52[255], stage0_52[256], stage0_52[257], stage0_52[258], stage0_52[259]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[103],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2057 (
      {stage0_52[260], stage0_52[261], stage0_52[262], stage0_52[263], stage0_52[264], stage0_52[265]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[104],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2058 (
      {stage0_52[266], stage0_52[267], stage0_52[268], stage0_52[269], stage0_52[270], stage0_52[271]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[105],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2059 (
      {stage0_52[272], stage0_52[273], stage0_52[274], stage0_52[275], stage0_52[276], stage0_52[277]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[106],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2060 (
      {stage0_52[278], stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[107],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2061 (
      {stage0_52[284], stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[108],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2062 (
      {stage0_52[290], stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[109],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2063 (
      {stage0_52[296], stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[110],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2064 (
      {stage0_52[302], stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[111],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2065 (
      {stage0_52[308], stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[112],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2066 (
      {stage0_52[314], stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[113],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2067 (
      {stage0_52[320], stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[114],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2068 (
      {stage0_52[326], stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[115],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2069 (
      {stage0_52[332], stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[116],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2070 (
      {stage0_52[338], stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[117],stage1_53[140],stage1_52[190]}
   );
   gpc606_5 gpc2071 (
      {stage0_52[344], stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[118],stage1_53[141],stage1_52[191]}
   );
   gpc606_5 gpc2072 (
      {stage0_52[350], stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[119],stage1_53[142],stage1_52[192]}
   );
   gpc606_5 gpc2073 (
      {stage0_52[356], stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[120],stage1_53[143],stage1_52[193]}
   );
   gpc606_5 gpc2074 (
      {stage0_52[362], stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[121],stage1_53[144],stage1_52[194]}
   );
   gpc606_5 gpc2075 (
      {stage0_52[368], stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[122],stage1_53[145],stage1_52[195]}
   );
   gpc606_5 gpc2076 (
      {stage0_52[374], stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[123],stage1_53[146],stage1_52[196]}
   );
   gpc606_5 gpc2077 (
      {stage0_52[380], stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[124],stage1_53[147],stage1_52[197]}
   );
   gpc606_5 gpc2078 (
      {stage0_52[386], stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[125],stage1_53[148],stage1_52[198]}
   );
   gpc606_5 gpc2079 (
      {stage0_52[392], stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[126],stage1_53[149],stage1_52[199]}
   );
   gpc606_5 gpc2080 (
      {stage0_52[398], stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[127],stage1_53[150],stage1_52[200]}
   );
   gpc606_5 gpc2081 (
      {stage0_52[404], stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409]},
      {stage0_54[216], stage0_54[217], stage0_54[218], stage0_54[219], stage0_54[220], stage0_54[221]},
      {stage1_56[36],stage1_55[99],stage1_54[128],stage1_53[151],stage1_52[201]}
   );
   gpc606_5 gpc2082 (
      {stage0_53[378], stage0_53[379], stage0_53[380], stage0_53[381], stage0_53[382], stage0_53[383]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[37],stage1_55[100],stage1_54[129],stage1_53[152]}
   );
   gpc606_5 gpc2083 (
      {stage0_53[384], stage0_53[385], stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[38],stage1_55[101],stage1_54[130],stage1_53[153]}
   );
   gpc606_5 gpc2084 (
      {stage0_53[390], stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[39],stage1_55[102],stage1_54[131],stage1_53[154]}
   );
   gpc606_5 gpc2085 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400], stage0_53[401]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[40],stage1_55[103],stage1_54[132],stage1_53[155]}
   );
   gpc606_5 gpc2086 (
      {stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405], stage0_53[406], stage0_53[407]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[41],stage1_55[104],stage1_54[133],stage1_53[156]}
   );
   gpc606_5 gpc2087 (
      {stage0_53[408], stage0_53[409], stage0_53[410], stage0_53[411], stage0_53[412], stage0_53[413]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[42],stage1_55[105],stage1_54[134],stage1_53[157]}
   );
   gpc606_5 gpc2088 (
      {stage0_53[414], stage0_53[415], stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[43],stage1_55[106],stage1_54[135],stage1_53[158]}
   );
   gpc606_5 gpc2089 (
      {stage0_53[420], stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[44],stage1_55[107],stage1_54[136],stage1_53[159]}
   );
   gpc606_5 gpc2090 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430], stage0_53[431]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[45],stage1_55[108],stage1_54[137],stage1_53[160]}
   );
   gpc606_5 gpc2091 (
      {stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435], stage0_53[436], stage0_53[437]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[46],stage1_55[109],stage1_54[138],stage1_53[161]}
   );
   gpc606_5 gpc2092 (
      {stage0_53[438], stage0_53[439], stage0_53[440], stage0_53[441], stage0_53[442], stage0_53[443]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[47],stage1_55[110],stage1_54[139],stage1_53[162]}
   );
   gpc606_5 gpc2093 (
      {stage0_53[444], stage0_53[445], stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[48],stage1_55[111],stage1_54[140],stage1_53[163]}
   );
   gpc606_5 gpc2094 (
      {stage0_53[450], stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[49],stage1_55[112],stage1_54[141],stage1_53[164]}
   );
   gpc606_5 gpc2095 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460], stage0_53[461]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[50],stage1_55[113],stage1_54[142],stage1_53[165]}
   );
   gpc606_5 gpc2096 (
      {stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465], stage0_53[466], stage0_53[467]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[51],stage1_55[114],stage1_54[143],stage1_53[166]}
   );
   gpc606_5 gpc2097 (
      {stage0_53[468], stage0_53[469], stage0_53[470], stage0_53[471], stage0_53[472], stage0_53[473]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[52],stage1_55[115],stage1_54[144],stage1_53[167]}
   );
   gpc606_5 gpc2098 (
      {stage0_53[474], stage0_53[475], stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[53],stage1_55[116],stage1_54[145],stage1_53[168]}
   );
   gpc606_5 gpc2099 (
      {stage0_53[480], stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[54],stage1_55[117],stage1_54[146],stage1_53[169]}
   );
   gpc606_5 gpc2100 (
      {stage0_53[486], stage0_53[487], stage0_53[488], stage0_53[489], stage0_53[490], stage0_53[491]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[55],stage1_55[118],stage1_54[147],stage1_53[170]}
   );
   gpc615_5 gpc2101 (
      {stage0_53[492], stage0_53[493], stage0_53[494], stage0_53[495], stage0_53[496]},
      {stage0_54[222]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[56],stage1_55[119],stage1_54[148],stage1_53[171]}
   );
   gpc606_5 gpc2102 (
      {stage0_54[223], stage0_54[224], stage0_54[225], stage0_54[226], stage0_54[227], stage0_54[228]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[20],stage1_56[57],stage1_55[120],stage1_54[149]}
   );
   gpc606_5 gpc2103 (
      {stage0_54[229], stage0_54[230], stage0_54[231], stage0_54[232], stage0_54[233], stage0_54[234]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[21],stage1_56[58],stage1_55[121],stage1_54[150]}
   );
   gpc606_5 gpc2104 (
      {stage0_54[235], stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[22],stage1_56[59],stage1_55[122],stage1_54[151]}
   );
   gpc615_5 gpc2105 (
      {stage0_54[241], stage0_54[242], stage0_54[243], stage0_54[244], stage0_54[245]},
      {stage0_55[120]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[23],stage1_56[60],stage1_55[123],stage1_54[152]}
   );
   gpc615_5 gpc2106 (
      {stage0_54[246], stage0_54[247], stage0_54[248], stage0_54[249], stage0_54[250]},
      {stage0_55[121]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[24],stage1_56[61],stage1_55[124],stage1_54[153]}
   );
   gpc615_5 gpc2107 (
      {stage0_54[251], stage0_54[252], stage0_54[253], stage0_54[254], stage0_54[255]},
      {stage0_55[122]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[25],stage1_56[62],stage1_55[125],stage1_54[154]}
   );
   gpc615_5 gpc2108 (
      {stage0_54[256], stage0_54[257], stage0_54[258], stage0_54[259], stage0_54[260]},
      {stage0_55[123]},
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage1_58[6],stage1_57[26],stage1_56[63],stage1_55[126],stage1_54[155]}
   );
   gpc615_5 gpc2109 (
      {stage0_54[261], stage0_54[262], stage0_54[263], stage0_54[264], stage0_54[265]},
      {stage0_55[124]},
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage1_58[7],stage1_57[27],stage1_56[64],stage1_55[127],stage1_54[156]}
   );
   gpc615_5 gpc2110 (
      {stage0_54[266], stage0_54[267], stage0_54[268], stage0_54[269], stage0_54[270]},
      {stage0_55[125]},
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage1_58[8],stage1_57[28],stage1_56[65],stage1_55[128],stage1_54[157]}
   );
   gpc615_5 gpc2111 (
      {stage0_54[271], stage0_54[272], stage0_54[273], stage0_54[274], stage0_54[275]},
      {stage0_55[126]},
      {stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59]},
      {stage1_58[9],stage1_57[29],stage1_56[66],stage1_55[129],stage1_54[158]}
   );
   gpc615_5 gpc2112 (
      {stage0_54[276], stage0_54[277], stage0_54[278], stage0_54[279], stage0_54[280]},
      {stage0_55[127]},
      {stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65]},
      {stage1_58[10],stage1_57[30],stage1_56[67],stage1_55[130],stage1_54[159]}
   );
   gpc615_5 gpc2113 (
      {stage0_54[281], stage0_54[282], stage0_54[283], stage0_54[284], stage0_54[285]},
      {stage0_55[128]},
      {stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71]},
      {stage1_58[11],stage1_57[31],stage1_56[68],stage1_55[131],stage1_54[160]}
   );
   gpc615_5 gpc2114 (
      {stage0_54[286], stage0_54[287], stage0_54[288], stage0_54[289], stage0_54[290]},
      {stage0_55[129]},
      {stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77]},
      {stage1_58[12],stage1_57[32],stage1_56[69],stage1_55[132],stage1_54[161]}
   );
   gpc615_5 gpc2115 (
      {stage0_54[291], stage0_54[292], stage0_54[293], stage0_54[294], stage0_54[295]},
      {stage0_55[130]},
      {stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83]},
      {stage1_58[13],stage1_57[33],stage1_56[70],stage1_55[133],stage1_54[162]}
   );
   gpc615_5 gpc2116 (
      {stage0_54[296], stage0_54[297], stage0_54[298], stage0_54[299], stage0_54[300]},
      {stage0_55[131]},
      {stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89]},
      {stage1_58[14],stage1_57[34],stage1_56[71],stage1_55[134],stage1_54[163]}
   );
   gpc615_5 gpc2117 (
      {stage0_54[301], stage0_54[302], stage0_54[303], stage0_54[304], stage0_54[305]},
      {stage0_55[132]},
      {stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95]},
      {stage1_58[15],stage1_57[35],stage1_56[72],stage1_55[135],stage1_54[164]}
   );
   gpc615_5 gpc2118 (
      {stage0_54[306], stage0_54[307], stage0_54[308], stage0_54[309], stage0_54[310]},
      {stage0_55[133]},
      {stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101]},
      {stage1_58[16],stage1_57[36],stage1_56[73],stage1_55[136],stage1_54[165]}
   );
   gpc615_5 gpc2119 (
      {stage0_54[311], stage0_54[312], stage0_54[313], stage0_54[314], stage0_54[315]},
      {stage0_55[134]},
      {stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107]},
      {stage1_58[17],stage1_57[37],stage1_56[74],stage1_55[137],stage1_54[166]}
   );
   gpc615_5 gpc2120 (
      {stage0_54[316], stage0_54[317], stage0_54[318], stage0_54[319], stage0_54[320]},
      {stage0_55[135]},
      {stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113]},
      {stage1_58[18],stage1_57[38],stage1_56[75],stage1_55[138],stage1_54[167]}
   );
   gpc615_5 gpc2121 (
      {stage0_54[321], stage0_54[322], stage0_54[323], stage0_54[324], stage0_54[325]},
      {stage0_55[136]},
      {stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119]},
      {stage1_58[19],stage1_57[39],stage1_56[76],stage1_55[139],stage1_54[168]}
   );
   gpc615_5 gpc2122 (
      {stage0_54[326], stage0_54[327], stage0_54[328], stage0_54[329], stage0_54[330]},
      {stage0_55[137]},
      {stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125]},
      {stage1_58[20],stage1_57[40],stage1_56[77],stage1_55[140],stage1_54[169]}
   );
   gpc615_5 gpc2123 (
      {stage0_54[331], stage0_54[332], stage0_54[333], stage0_54[334], stage0_54[335]},
      {stage0_55[138]},
      {stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131]},
      {stage1_58[21],stage1_57[41],stage1_56[78],stage1_55[141],stage1_54[170]}
   );
   gpc615_5 gpc2124 (
      {stage0_54[336], stage0_54[337], stage0_54[338], stage0_54[339], stage0_54[340]},
      {stage0_55[139]},
      {stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137]},
      {stage1_58[22],stage1_57[42],stage1_56[79],stage1_55[142],stage1_54[171]}
   );
   gpc615_5 gpc2125 (
      {stage0_54[341], stage0_54[342], stage0_54[343], stage0_54[344], stage0_54[345]},
      {stage0_55[140]},
      {stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143]},
      {stage1_58[23],stage1_57[43],stage1_56[80],stage1_55[143],stage1_54[172]}
   );
   gpc615_5 gpc2126 (
      {stage0_54[346], stage0_54[347], stage0_54[348], stage0_54[349], stage0_54[350]},
      {stage0_55[141]},
      {stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149]},
      {stage1_58[24],stage1_57[44],stage1_56[81],stage1_55[144],stage1_54[173]}
   );
   gpc615_5 gpc2127 (
      {stage0_54[351], stage0_54[352], stage0_54[353], stage0_54[354], stage0_54[355]},
      {stage0_55[142]},
      {stage0_56[150], stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155]},
      {stage1_58[25],stage1_57[45],stage1_56[82],stage1_55[145],stage1_54[174]}
   );
   gpc615_5 gpc2128 (
      {stage0_54[356], stage0_54[357], stage0_54[358], stage0_54[359], stage0_54[360]},
      {stage0_55[143]},
      {stage0_56[156], stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161]},
      {stage1_58[26],stage1_57[46],stage1_56[83],stage1_55[146],stage1_54[175]}
   );
   gpc615_5 gpc2129 (
      {stage0_54[361], stage0_54[362], stage0_54[363], stage0_54[364], stage0_54[365]},
      {stage0_55[144]},
      {stage0_56[162], stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167]},
      {stage1_58[27],stage1_57[47],stage1_56[84],stage1_55[147],stage1_54[176]}
   );
   gpc615_5 gpc2130 (
      {stage0_54[366], stage0_54[367], stage0_54[368], stage0_54[369], stage0_54[370]},
      {stage0_55[145]},
      {stage0_56[168], stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173]},
      {stage1_58[28],stage1_57[48],stage1_56[85],stage1_55[148],stage1_54[177]}
   );
   gpc615_5 gpc2131 (
      {stage0_54[371], stage0_54[372], stage0_54[373], stage0_54[374], stage0_54[375]},
      {stage0_55[146]},
      {stage0_56[174], stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179]},
      {stage1_58[29],stage1_57[49],stage1_56[86],stage1_55[149],stage1_54[178]}
   );
   gpc615_5 gpc2132 (
      {stage0_54[376], stage0_54[377], stage0_54[378], stage0_54[379], stage0_54[380]},
      {stage0_55[147]},
      {stage0_56[180], stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185]},
      {stage1_58[30],stage1_57[50],stage1_56[87],stage1_55[150],stage1_54[179]}
   );
   gpc615_5 gpc2133 (
      {stage0_54[381], stage0_54[382], stage0_54[383], stage0_54[384], stage0_54[385]},
      {stage0_55[148]},
      {stage0_56[186], stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191]},
      {stage1_58[31],stage1_57[51],stage1_56[88],stage1_55[151],stage1_54[180]}
   );
   gpc615_5 gpc2134 (
      {stage0_54[386], stage0_54[387], stage0_54[388], stage0_54[389], stage0_54[390]},
      {stage0_55[149]},
      {stage0_56[192], stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197]},
      {stage1_58[32],stage1_57[52],stage1_56[89],stage1_55[152],stage1_54[181]}
   );
   gpc615_5 gpc2135 (
      {stage0_54[391], stage0_54[392], stage0_54[393], stage0_54[394], stage0_54[395]},
      {stage0_55[150]},
      {stage0_56[198], stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203]},
      {stage1_58[33],stage1_57[53],stage1_56[90],stage1_55[153],stage1_54[182]}
   );
   gpc615_5 gpc2136 (
      {stage0_54[396], stage0_54[397], stage0_54[398], stage0_54[399], stage0_54[400]},
      {stage0_55[151]},
      {stage0_56[204], stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209]},
      {stage1_58[34],stage1_57[54],stage1_56[91],stage1_55[154],stage1_54[183]}
   );
   gpc615_5 gpc2137 (
      {stage0_54[401], stage0_54[402], stage0_54[403], stage0_54[404], stage0_54[405]},
      {stage0_55[152]},
      {stage0_56[210], stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215]},
      {stage1_58[35],stage1_57[55],stage1_56[92],stage1_55[155],stage1_54[184]}
   );
   gpc615_5 gpc2138 (
      {stage0_54[406], stage0_54[407], stage0_54[408], stage0_54[409], stage0_54[410]},
      {stage0_55[153]},
      {stage0_56[216], stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221]},
      {stage1_58[36],stage1_57[56],stage1_56[93],stage1_55[156],stage1_54[185]}
   );
   gpc615_5 gpc2139 (
      {stage0_54[411], stage0_54[412], stage0_54[413], stage0_54[414], stage0_54[415]},
      {stage0_55[154]},
      {stage0_56[222], stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227]},
      {stage1_58[37],stage1_57[57],stage1_56[94],stage1_55[157],stage1_54[186]}
   );
   gpc615_5 gpc2140 (
      {stage0_54[416], stage0_54[417], stage0_54[418], stage0_54[419], stage0_54[420]},
      {stage0_55[155]},
      {stage0_56[228], stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233]},
      {stage1_58[38],stage1_57[58],stage1_56[95],stage1_55[158],stage1_54[187]}
   );
   gpc615_5 gpc2141 (
      {stage0_54[421], stage0_54[422], stage0_54[423], stage0_54[424], stage0_54[425]},
      {stage0_55[156]},
      {stage0_56[234], stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239]},
      {stage1_58[39],stage1_57[59],stage1_56[96],stage1_55[159],stage1_54[188]}
   );
   gpc615_5 gpc2142 (
      {stage0_54[426], stage0_54[427], stage0_54[428], stage0_54[429], stage0_54[430]},
      {stage0_55[157]},
      {stage0_56[240], stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245]},
      {stage1_58[40],stage1_57[60],stage1_56[97],stage1_55[160],stage1_54[189]}
   );
   gpc615_5 gpc2143 (
      {stage0_54[431], stage0_54[432], stage0_54[433], stage0_54[434], stage0_54[435]},
      {stage0_55[158]},
      {stage0_56[246], stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251]},
      {stage1_58[41],stage1_57[61],stage1_56[98],stage1_55[161],stage1_54[190]}
   );
   gpc615_5 gpc2144 (
      {stage0_54[436], stage0_54[437], stage0_54[438], stage0_54[439], stage0_54[440]},
      {stage0_55[159]},
      {stage0_56[252], stage0_56[253], stage0_56[254], stage0_56[255], stage0_56[256], stage0_56[257]},
      {stage1_58[42],stage1_57[62],stage1_56[99],stage1_55[162],stage1_54[191]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[160], stage0_55[161], stage0_55[162], stage0_55[163], stage0_55[164], stage0_55[165]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[43],stage1_57[63],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[166], stage0_55[167], stage0_55[168], stage0_55[169], stage0_55[170], stage0_55[171]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[44],stage1_57[64],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2147 (
      {stage0_55[172], stage0_55[173], stage0_55[174], stage0_55[175], stage0_55[176], stage0_55[177]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[45],stage1_57[65],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2148 (
      {stage0_55[178], stage0_55[179], stage0_55[180], stage0_55[181], stage0_55[182], stage0_55[183]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[46],stage1_57[66],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2149 (
      {stage0_55[184], stage0_55[185], stage0_55[186], stage0_55[187], stage0_55[188], stage0_55[189]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[47],stage1_57[67],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2150 (
      {stage0_55[190], stage0_55[191], stage0_55[192], stage0_55[193], stage0_55[194], stage0_55[195]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[48],stage1_57[68],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2151 (
      {stage0_55[196], stage0_55[197], stage0_55[198], stage0_55[199], stage0_55[200], stage0_55[201]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[49],stage1_57[69],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2152 (
      {stage0_55[202], stage0_55[203], stage0_55[204], stage0_55[205], stage0_55[206], stage0_55[207]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[50],stage1_57[70],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2153 (
      {stage0_55[208], stage0_55[209], stage0_55[210], stage0_55[211], stage0_55[212], stage0_55[213]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[51],stage1_57[71],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2154 (
      {stage0_55[214], stage0_55[215], stage0_55[216], stage0_55[217], stage0_55[218], stage0_55[219]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[52],stage1_57[72],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2155 (
      {stage0_55[220], stage0_55[221], stage0_55[222], stage0_55[223], stage0_55[224], stage0_55[225]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[53],stage1_57[73],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2156 (
      {stage0_55[226], stage0_55[227], stage0_55[228], stage0_55[229], stage0_55[230], stage0_55[231]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[54],stage1_57[74],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2157 (
      {stage0_55[232], stage0_55[233], stage0_55[234], stage0_55[235], stage0_55[236], stage0_55[237]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[55],stage1_57[75],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2158 (
      {stage0_55[238], stage0_55[239], stage0_55[240], stage0_55[241], stage0_55[242], stage0_55[243]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[56],stage1_57[76],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2159 (
      {stage0_55[244], stage0_55[245], stage0_55[246], stage0_55[247], stage0_55[248], stage0_55[249]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[57],stage1_57[77],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2160 (
      {stage0_55[250], stage0_55[251], stage0_55[252], stage0_55[253], stage0_55[254], stage0_55[255]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[58],stage1_57[78],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2161 (
      {stage0_55[256], stage0_55[257], stage0_55[258], stage0_55[259], stage0_55[260], stage0_55[261]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[59],stage1_57[79],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2162 (
      {stage0_55[262], stage0_55[263], stage0_55[264], stage0_55[265], stage0_55[266], stage0_55[267]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[60],stage1_57[80],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2163 (
      {stage0_55[268], stage0_55[269], stage0_55[270], stage0_55[271], stage0_55[272], stage0_55[273]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[61],stage1_57[81],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2164 (
      {stage0_55[274], stage0_55[275], stage0_55[276], stage0_55[277], stage0_55[278], stage0_55[279]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[62],stage1_57[82],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2165 (
      {stage0_55[280], stage0_55[281], stage0_55[282], stage0_55[283], stage0_55[284], stage0_55[285]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[63],stage1_57[83],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2166 (
      {stage0_55[286], stage0_55[287], stage0_55[288], stage0_55[289], stage0_55[290], stage0_55[291]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[64],stage1_57[84],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2167 (
      {stage0_55[292], stage0_55[293], stage0_55[294], stage0_55[295], stage0_55[296], stage0_55[297]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[65],stage1_57[85],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2168 (
      {stage0_55[298], stage0_55[299], stage0_55[300], stage0_55[301], stage0_55[302], stage0_55[303]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[66],stage1_57[86],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2169 (
      {stage0_55[304], stage0_55[305], stage0_55[306], stage0_55[307], stage0_55[308], stage0_55[309]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[67],stage1_57[87],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2170 (
      {stage0_55[310], stage0_55[311], stage0_55[312], stage0_55[313], stage0_55[314], stage0_55[315]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[68],stage1_57[88],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2171 (
      {stage0_55[316], stage0_55[317], stage0_55[318], stage0_55[319], stage0_55[320], stage0_55[321]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[69],stage1_57[89],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2172 (
      {stage0_55[322], stage0_55[323], stage0_55[324], stage0_55[325], stage0_55[326], stage0_55[327]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[70],stage1_57[90],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2173 (
      {stage0_55[328], stage0_55[329], stage0_55[330], stage0_55[331], stage0_55[332], stage0_55[333]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[71],stage1_57[91],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2174 (
      {stage0_55[334], stage0_55[335], stage0_55[336], stage0_55[337], stage0_55[338], stage0_55[339]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[72],stage1_57[92],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2175 (
      {stage0_55[340], stage0_55[341], stage0_55[342], stage0_55[343], stage0_55[344], stage0_55[345]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[73],stage1_57[93],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2176 (
      {stage0_55[346], stage0_55[347], stage0_55[348], stage0_55[349], stage0_55[350], stage0_55[351]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[74],stage1_57[94],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2177 (
      {stage0_55[352], stage0_55[353], stage0_55[354], stage0_55[355], stage0_55[356], stage0_55[357]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[75],stage1_57[95],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2178 (
      {stage0_55[358], stage0_55[359], stage0_55[360], stage0_55[361], stage0_55[362], stage0_55[363]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[76],stage1_57[96],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2179 (
      {stage0_55[364], stage0_55[365], stage0_55[366], stage0_55[367], stage0_55[368], stage0_55[369]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[77],stage1_57[97],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2180 (
      {stage0_55[370], stage0_55[371], stage0_55[372], stage0_55[373], stage0_55[374], stage0_55[375]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[78],stage1_57[98],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2181 (
      {stage0_55[376], stage0_55[377], stage0_55[378], stage0_55[379], stage0_55[380], stage0_55[381]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[79],stage1_57[99],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2182 (
      {stage0_55[382], stage0_55[383], stage0_55[384], stage0_55[385], stage0_55[386], stage0_55[387]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[80],stage1_57[100],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2183 (
      {stage0_55[388], stage0_55[389], stage0_55[390], stage0_55[391], stage0_55[392], stage0_55[393]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[81],stage1_57[101],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2184 (
      {stage0_55[394], stage0_55[395], stage0_55[396], stage0_55[397], stage0_55[398], stage0_55[399]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[82],stage1_57[102],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2185 (
      {stage0_55[400], stage0_55[401], stage0_55[402], stage0_55[403], stage0_55[404], stage0_55[405]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[83],stage1_57[103],stage1_56[140],stage1_55[203]}
   );
   gpc606_5 gpc2186 (
      {stage0_55[406], stage0_55[407], stage0_55[408], stage0_55[409], stage0_55[410], stage0_55[411]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[84],stage1_57[104],stage1_56[141],stage1_55[204]}
   );
   gpc606_5 gpc2187 (
      {stage0_55[412], stage0_55[413], stage0_55[414], stage0_55[415], stage0_55[416], stage0_55[417]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[85],stage1_57[105],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2188 (
      {stage0_55[418], stage0_55[419], stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[86],stage1_57[106],stage1_56[143],stage1_55[206]}
   );
   gpc606_5 gpc2189 (
      {stage0_55[424], stage0_55[425], stage0_55[426], stage0_55[427], stage0_55[428], stage0_55[429]},
      {stage0_57[264], stage0_57[265], stage0_57[266], stage0_57[267], stage0_57[268], stage0_57[269]},
      {stage1_59[44],stage1_58[87],stage1_57[107],stage1_56[144],stage1_55[207]}
   );
   gpc606_5 gpc2190 (
      {stage0_55[430], stage0_55[431], stage0_55[432], stage0_55[433], stage0_55[434], stage0_55[435]},
      {stage0_57[270], stage0_57[271], stage0_57[272], stage0_57[273], stage0_57[274], stage0_57[275]},
      {stage1_59[45],stage1_58[88],stage1_57[108],stage1_56[145],stage1_55[208]}
   );
   gpc606_5 gpc2191 (
      {stage0_55[436], stage0_55[437], stage0_55[438], stage0_55[439], stage0_55[440], stage0_55[441]},
      {stage0_57[276], stage0_57[277], stage0_57[278], stage0_57[279], stage0_57[280], stage0_57[281]},
      {stage1_59[46],stage1_58[89],stage1_57[109],stage1_56[146],stage1_55[209]}
   );
   gpc606_5 gpc2192 (
      {stage0_55[442], stage0_55[443], stage0_55[444], stage0_55[445], stage0_55[446], stage0_55[447]},
      {stage0_57[282], stage0_57[283], stage0_57[284], stage0_57[285], stage0_57[286], stage0_57[287]},
      {stage1_59[47],stage1_58[90],stage1_57[110],stage1_56[147],stage1_55[210]}
   );
   gpc606_5 gpc2193 (
      {stage0_55[448], stage0_55[449], stage0_55[450], stage0_55[451], stage0_55[452], stage0_55[453]},
      {stage0_57[288], stage0_57[289], stage0_57[290], stage0_57[291], stage0_57[292], stage0_57[293]},
      {stage1_59[48],stage1_58[91],stage1_57[111],stage1_56[148],stage1_55[211]}
   );
   gpc606_5 gpc2194 (
      {stage0_55[454], stage0_55[455], stage0_55[456], stage0_55[457], stage0_55[458], stage0_55[459]},
      {stage0_57[294], stage0_57[295], stage0_57[296], stage0_57[297], stage0_57[298], stage0_57[299]},
      {stage1_59[49],stage1_58[92],stage1_57[112],stage1_56[149],stage1_55[212]}
   );
   gpc606_5 gpc2195 (
      {stage0_55[460], stage0_55[461], stage0_55[462], stage0_55[463], stage0_55[464], stage0_55[465]},
      {stage0_57[300], stage0_57[301], stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305]},
      {stage1_59[50],stage1_58[93],stage1_57[113],stage1_56[150],stage1_55[213]}
   );
   gpc606_5 gpc2196 (
      {stage0_55[466], stage0_55[467], stage0_55[468], stage0_55[469], stage0_55[470], stage0_55[471]},
      {stage0_57[306], stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage1_59[51],stage1_58[94],stage1_57[114],stage1_56[151],stage1_55[214]}
   );
   gpc606_5 gpc2197 (
      {stage0_55[472], stage0_55[473], stage0_55[474], stage0_55[475], stage0_55[476], stage0_55[477]},
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316], stage0_57[317]},
      {stage1_59[52],stage1_58[95],stage1_57[115],stage1_56[152],stage1_55[215]}
   );
   gpc615_5 gpc2198 (
      {stage0_55[478], stage0_55[479], stage0_55[480], stage0_55[481], stage0_55[482]},
      {stage0_56[258]},
      {stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321], stage0_57[322], stage0_57[323]},
      {stage1_59[53],stage1_58[96],stage1_57[116],stage1_56[153],stage1_55[216]}
   );
   gpc615_5 gpc2199 (
      {stage0_55[483], stage0_55[484], stage0_55[485], stage0_55[486], stage0_55[487]},
      {stage0_56[259]},
      {stage0_57[324], stage0_57[325], stage0_57[326], stage0_57[327], stage0_57[328], stage0_57[329]},
      {stage1_59[54],stage1_58[97],stage1_57[117],stage1_56[154],stage1_55[217]}
   );
   gpc615_5 gpc2200 (
      {stage0_55[488], stage0_55[489], stage0_55[490], stage0_55[491], stage0_55[492]},
      {stage0_56[260]},
      {stage0_57[330], stage0_57[331], stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335]},
      {stage1_59[55],stage1_58[98],stage1_57[118],stage1_56[155],stage1_55[218]}
   );
   gpc615_5 gpc2201 (
      {stage0_55[493], stage0_55[494], stage0_55[495], stage0_55[496], stage0_55[497]},
      {stage0_56[261]},
      {stage0_57[336], stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage1_59[56],stage1_58[99],stage1_57[119],stage1_56[156],stage1_55[219]}
   );
   gpc615_5 gpc2202 (
      {stage0_55[498], stage0_55[499], stage0_55[500], stage0_55[501], stage0_55[502]},
      {stage0_56[262]},
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346], stage0_57[347]},
      {stage1_59[57],stage1_58[100],stage1_57[120],stage1_56[157],stage1_55[220]}
   );
   gpc615_5 gpc2203 (
      {stage0_55[503], stage0_55[504], stage0_55[505], stage0_55[506], stage0_55[507]},
      {stage0_56[263]},
      {stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351], stage0_57[352], stage0_57[353]},
      {stage1_59[58],stage1_58[101],stage1_57[121],stage1_56[158],stage1_55[221]}
   );
   gpc606_5 gpc2204 (
      {stage0_56[264], stage0_56[265], stage0_56[266], stage0_56[267], stage0_56[268], stage0_56[269]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[59],stage1_58[102],stage1_57[122],stage1_56[159]}
   );
   gpc606_5 gpc2205 (
      {stage0_56[270], stage0_56[271], stage0_56[272], stage0_56[273], stage0_56[274], stage0_56[275]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[60],stage1_58[103],stage1_57[123],stage1_56[160]}
   );
   gpc606_5 gpc2206 (
      {stage0_56[276], stage0_56[277], stage0_56[278], stage0_56[279], stage0_56[280], stage0_56[281]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[61],stage1_58[104],stage1_57[124],stage1_56[161]}
   );
   gpc606_5 gpc2207 (
      {stage0_56[282], stage0_56[283], stage0_56[284], stage0_56[285], stage0_56[286], stage0_56[287]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[62],stage1_58[105],stage1_57[125],stage1_56[162]}
   );
   gpc606_5 gpc2208 (
      {stage0_56[288], stage0_56[289], stage0_56[290], stage0_56[291], stage0_56[292], stage0_56[293]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[63],stage1_58[106],stage1_57[126],stage1_56[163]}
   );
   gpc606_5 gpc2209 (
      {stage0_56[294], stage0_56[295], stage0_56[296], stage0_56[297], stage0_56[298], stage0_56[299]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[64],stage1_58[107],stage1_57[127],stage1_56[164]}
   );
   gpc606_5 gpc2210 (
      {stage0_56[300], stage0_56[301], stage0_56[302], stage0_56[303], stage0_56[304], stage0_56[305]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[65],stage1_58[108],stage1_57[128],stage1_56[165]}
   );
   gpc606_5 gpc2211 (
      {stage0_56[306], stage0_56[307], stage0_56[308], stage0_56[309], stage0_56[310], stage0_56[311]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[66],stage1_58[109],stage1_57[129],stage1_56[166]}
   );
   gpc606_5 gpc2212 (
      {stage0_56[312], stage0_56[313], stage0_56[314], stage0_56[315], stage0_56[316], stage0_56[317]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[67],stage1_58[110],stage1_57[130],stage1_56[167]}
   );
   gpc606_5 gpc2213 (
      {stage0_56[318], stage0_56[319], stage0_56[320], stage0_56[321], stage0_56[322], stage0_56[323]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[68],stage1_58[111],stage1_57[131],stage1_56[168]}
   );
   gpc606_5 gpc2214 (
      {stage0_56[324], stage0_56[325], stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[69],stage1_58[112],stage1_57[132],stage1_56[169]}
   );
   gpc606_5 gpc2215 (
      {stage0_56[330], stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[70],stage1_58[113],stage1_57[133],stage1_56[170]}
   );
   gpc606_5 gpc2216 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340], stage0_56[341]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[71],stage1_58[114],stage1_57[134],stage1_56[171]}
   );
   gpc606_5 gpc2217 (
      {stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345], stage0_56[346], stage0_56[347]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[72],stage1_58[115],stage1_57[135],stage1_56[172]}
   );
   gpc606_5 gpc2218 (
      {stage0_56[348], stage0_56[349], stage0_56[350], stage0_56[351], stage0_56[352], stage0_56[353]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[73],stage1_58[116],stage1_57[136],stage1_56[173]}
   );
   gpc606_5 gpc2219 (
      {stage0_56[354], stage0_56[355], stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[74],stage1_58[117],stage1_57[137],stage1_56[174]}
   );
   gpc606_5 gpc2220 (
      {stage0_56[360], stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[75],stage1_58[118],stage1_57[138],stage1_56[175]}
   );
   gpc606_5 gpc2221 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370], stage0_56[371]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[76],stage1_58[119],stage1_57[139],stage1_56[176]}
   );
   gpc606_5 gpc2222 (
      {stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375], stage0_56[376], stage0_56[377]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[77],stage1_58[120],stage1_57[140],stage1_56[177]}
   );
   gpc606_5 gpc2223 (
      {stage0_56[378], stage0_56[379], stage0_56[380], stage0_56[381], stage0_56[382], stage0_56[383]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[78],stage1_58[121],stage1_57[141],stage1_56[178]}
   );
   gpc606_5 gpc2224 (
      {stage0_56[384], stage0_56[385], stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[79],stage1_58[122],stage1_57[142],stage1_56[179]}
   );
   gpc606_5 gpc2225 (
      {stage0_56[390], stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[80],stage1_58[123],stage1_57[143],stage1_56[180]}
   );
   gpc606_5 gpc2226 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400], stage0_56[401]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[81],stage1_58[124],stage1_57[144],stage1_56[181]}
   );
   gpc606_5 gpc2227 (
      {stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405], stage0_56[406], stage0_56[407]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[82],stage1_58[125],stage1_57[145],stage1_56[182]}
   );
   gpc606_5 gpc2228 (
      {stage0_56[408], stage0_56[409], stage0_56[410], stage0_56[411], stage0_56[412], stage0_56[413]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[83],stage1_58[126],stage1_57[146],stage1_56[183]}
   );
   gpc606_5 gpc2229 (
      {stage0_56[414], stage0_56[415], stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[84],stage1_58[127],stage1_57[147],stage1_56[184]}
   );
   gpc606_5 gpc2230 (
      {stage0_56[420], stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[85],stage1_58[128],stage1_57[148],stage1_56[185]}
   );
   gpc606_5 gpc2231 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430], stage0_56[431]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[86],stage1_58[129],stage1_57[149],stage1_56[186]}
   );
   gpc606_5 gpc2232 (
      {stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435], stage0_56[436], stage0_56[437]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[87],stage1_58[130],stage1_57[150],stage1_56[187]}
   );
   gpc606_5 gpc2233 (
      {stage0_56[438], stage0_56[439], stage0_56[440], stage0_56[441], stage0_56[442], stage0_56[443]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[88],stage1_58[131],stage1_57[151],stage1_56[188]}
   );
   gpc606_5 gpc2234 (
      {stage0_57[354], stage0_57[355], stage0_57[356], stage0_57[357], stage0_57[358], stage0_57[359]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[30],stage1_59[89],stage1_58[132],stage1_57[152]}
   );
   gpc606_5 gpc2235 (
      {stage0_57[360], stage0_57[361], stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[31],stage1_59[90],stage1_58[133],stage1_57[153]}
   );
   gpc606_5 gpc2236 (
      {stage0_57[366], stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[32],stage1_59[91],stage1_58[134],stage1_57[154]}
   );
   gpc606_5 gpc2237 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376], stage0_57[377]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[33],stage1_59[92],stage1_58[135],stage1_57[155]}
   );
   gpc606_5 gpc2238 (
      {stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381], stage0_57[382], stage0_57[383]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[34],stage1_59[93],stage1_58[136],stage1_57[156]}
   );
   gpc606_5 gpc2239 (
      {stage0_57[384], stage0_57[385], stage0_57[386], stage0_57[387], stage0_57[388], stage0_57[389]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[35],stage1_59[94],stage1_58[137],stage1_57[157]}
   );
   gpc606_5 gpc2240 (
      {stage0_57[390], stage0_57[391], stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[36],stage1_59[95],stage1_58[138],stage1_57[158]}
   );
   gpc606_5 gpc2241 (
      {stage0_57[396], stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[37],stage1_59[96],stage1_58[139],stage1_57[159]}
   );
   gpc606_5 gpc2242 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406], stage0_57[407]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[38],stage1_59[97],stage1_58[140],stage1_57[160]}
   );
   gpc606_5 gpc2243 (
      {stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411], stage0_57[412], stage0_57[413]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[39],stage1_59[98],stage1_58[141],stage1_57[161]}
   );
   gpc606_5 gpc2244 (
      {stage0_57[414], stage0_57[415], stage0_57[416], stage0_57[417], stage0_57[418], stage0_57[419]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[40],stage1_59[99],stage1_58[142],stage1_57[162]}
   );
   gpc606_5 gpc2245 (
      {stage0_57[420], stage0_57[421], stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[41],stage1_59[100],stage1_58[143],stage1_57[163]}
   );
   gpc606_5 gpc2246 (
      {stage0_57[426], stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[42],stage1_59[101],stage1_58[144],stage1_57[164]}
   );
   gpc606_5 gpc2247 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436], stage0_57[437]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[43],stage1_59[102],stage1_58[145],stage1_57[165]}
   );
   gpc606_5 gpc2248 (
      {stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441], stage0_57[442], stage0_57[443]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[44],stage1_59[103],stage1_58[146],stage1_57[166]}
   );
   gpc606_5 gpc2249 (
      {stage0_57[444], stage0_57[445], stage0_57[446], stage0_57[447], stage0_57[448], stage0_57[449]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[45],stage1_59[104],stage1_58[147],stage1_57[167]}
   );
   gpc606_5 gpc2250 (
      {stage0_57[450], stage0_57[451], stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[46],stage1_59[105],stage1_58[148],stage1_57[168]}
   );
   gpc606_5 gpc2251 (
      {stage0_57[456], stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[47],stage1_59[106],stage1_58[149],stage1_57[169]}
   );
   gpc606_5 gpc2252 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466], stage0_57[467]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[48],stage1_59[107],stage1_58[150],stage1_57[170]}
   );
   gpc606_5 gpc2253 (
      {stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471], stage0_57[472], stage0_57[473]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[49],stage1_59[108],stage1_58[151],stage1_57[171]}
   );
   gpc606_5 gpc2254 (
      {stage0_57[474], stage0_57[475], stage0_57[476], stage0_57[477], stage0_57[478], stage0_57[479]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[50],stage1_59[109],stage1_58[152],stage1_57[172]}
   );
   gpc606_5 gpc2255 (
      {stage0_57[480], stage0_57[481], stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[51],stage1_59[110],stage1_58[153],stage1_57[173]}
   );
   gpc606_5 gpc2256 (
      {stage0_57[486], stage0_57[487], stage0_57[488], stage0_57[489], stage0_57[490], stage0_57[491]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[52],stage1_59[111],stage1_58[154],stage1_57[174]}
   );
   gpc606_5 gpc2257 (
      {stage0_57[492], stage0_57[493], stage0_57[494], stage0_57[495], stage0_57[496], stage0_57[497]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[53],stage1_59[112],stage1_58[155],stage1_57[175]}
   );
   gpc606_5 gpc2258 (
      {stage0_57[498], stage0_57[499], stage0_57[500], stage0_57[501], stage0_57[502], stage0_57[503]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[54],stage1_59[113],stage1_58[156],stage1_57[176]}
   );
   gpc606_5 gpc2259 (
      {stage0_57[504], stage0_57[505], stage0_57[506], stage0_57[507], stage0_57[508], stage0_57[509]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[55],stage1_59[114],stage1_58[157],stage1_57[177]}
   );
   gpc2135_5 gpc2260 (
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184]},
      {stage0_59[156], stage0_59[157], stage0_59[158]},
      {stage0_60[0]},
      {stage0_61[0], stage0_61[1]},
      {stage1_62[0],stage1_61[26],stage1_60[56],stage1_59[115],stage1_58[158]}
   );
   gpc2135_5 gpc2261 (
      {stage0_58[185], stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189]},
      {stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage0_60[1]},
      {stage0_61[2], stage0_61[3]},
      {stage1_62[1],stage1_61[27],stage1_60[57],stage1_59[116],stage1_58[159]}
   );
   gpc2135_5 gpc2262 (
      {stage0_58[190], stage0_58[191], stage0_58[192], stage0_58[193], stage0_58[194]},
      {stage0_59[162], stage0_59[163], stage0_59[164]},
      {stage0_60[2]},
      {stage0_61[4], stage0_61[5]},
      {stage1_62[2],stage1_61[28],stage1_60[58],stage1_59[117],stage1_58[160]}
   );
   gpc2135_5 gpc2263 (
      {stage0_58[195], stage0_58[196], stage0_58[197], stage0_58[198], stage0_58[199]},
      {stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage0_60[3]},
      {stage0_61[6], stage0_61[7]},
      {stage1_62[3],stage1_61[29],stage1_60[59],stage1_59[118],stage1_58[161]}
   );
   gpc2135_5 gpc2264 (
      {stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203], stage0_58[204]},
      {stage0_59[168], stage0_59[169], stage0_59[170]},
      {stage0_60[4]},
      {stage0_61[8], stage0_61[9]},
      {stage1_62[4],stage1_61[30],stage1_60[60],stage1_59[119],stage1_58[162]}
   );
   gpc2135_5 gpc2265 (
      {stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage0_60[5]},
      {stage0_61[10], stage0_61[11]},
      {stage1_62[5],stage1_61[31],stage1_60[61],stage1_59[120],stage1_58[163]}
   );
   gpc2135_5 gpc2266 (
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214]},
      {stage0_59[174], stage0_59[175], stage0_59[176]},
      {stage0_60[6]},
      {stage0_61[12], stage0_61[13]},
      {stage1_62[6],stage1_61[32],stage1_60[62],stage1_59[121],stage1_58[164]}
   );
   gpc2135_5 gpc2267 (
      {stage0_58[215], stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219]},
      {stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage0_60[7]},
      {stage0_61[14], stage0_61[15]},
      {stage1_62[7],stage1_61[33],stage1_60[63],stage1_59[122],stage1_58[165]}
   );
   gpc2135_5 gpc2268 (
      {stage0_58[220], stage0_58[221], stage0_58[222], stage0_58[223], stage0_58[224]},
      {stage0_59[180], stage0_59[181], stage0_59[182]},
      {stage0_60[8]},
      {stage0_61[16], stage0_61[17]},
      {stage1_62[8],stage1_61[34],stage1_60[64],stage1_59[123],stage1_58[166]}
   );
   gpc2135_5 gpc2269 (
      {stage0_58[225], stage0_58[226], stage0_58[227], stage0_58[228], stage0_58[229]},
      {stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage0_60[9]},
      {stage0_61[18], stage0_61[19]},
      {stage1_62[9],stage1_61[35],stage1_60[65],stage1_59[124],stage1_58[167]}
   );
   gpc2135_5 gpc2270 (
      {stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233], stage0_58[234]},
      {stage0_59[186], stage0_59[187], stage0_59[188]},
      {stage0_60[10]},
      {stage0_61[20], stage0_61[21]},
      {stage1_62[10],stage1_61[36],stage1_60[66],stage1_59[125],stage1_58[168]}
   );
   gpc2135_5 gpc2271 (
      {stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage0_60[11]},
      {stage0_61[22], stage0_61[23]},
      {stage1_62[11],stage1_61[37],stage1_60[67],stage1_59[126],stage1_58[169]}
   );
   gpc2135_5 gpc2272 (
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244]},
      {stage0_59[192], stage0_59[193], stage0_59[194]},
      {stage0_60[12]},
      {stage0_61[24], stage0_61[25]},
      {stage1_62[12],stage1_61[38],stage1_60[68],stage1_59[127],stage1_58[170]}
   );
   gpc2135_5 gpc2273 (
      {stage0_58[245], stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249]},
      {stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage0_60[13]},
      {stage0_61[26], stage0_61[27]},
      {stage1_62[13],stage1_61[39],stage1_60[69],stage1_59[128],stage1_58[171]}
   );
   gpc2135_5 gpc2274 (
      {stage0_58[250], stage0_58[251], stage0_58[252], stage0_58[253], stage0_58[254]},
      {stage0_59[198], stage0_59[199], stage0_59[200]},
      {stage0_60[14]},
      {stage0_61[28], stage0_61[29]},
      {stage1_62[14],stage1_61[40],stage1_60[70],stage1_59[129],stage1_58[172]}
   );
   gpc2135_5 gpc2275 (
      {stage0_58[255], stage0_58[256], stage0_58[257], stage0_58[258], stage0_58[259]},
      {stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage0_60[15]},
      {stage0_61[30], stage0_61[31]},
      {stage1_62[15],stage1_61[41],stage1_60[71],stage1_59[130],stage1_58[173]}
   );
   gpc1163_5 gpc2276 (
      {stage0_58[260], stage0_58[261], stage0_58[262]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage0_60[16]},
      {stage0_61[32]},
      {stage1_62[16],stage1_61[42],stage1_60[72],stage1_59[131],stage1_58[174]}
   );
   gpc1163_5 gpc2277 (
      {stage0_58[263], stage0_58[264], stage0_58[265]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage0_60[17]},
      {stage0_61[33]},
      {stage1_62[17],stage1_61[43],stage1_60[73],stage1_59[132],stage1_58[175]}
   );
   gpc1163_5 gpc2278 (
      {stage0_58[266], stage0_58[267], stage0_58[268]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage0_60[18]},
      {stage0_61[34]},
      {stage1_62[18],stage1_61[44],stage1_60[74],stage1_59[133],stage1_58[176]}
   );
   gpc1163_5 gpc2279 (
      {stage0_58[269], stage0_58[270], stage0_58[271]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage0_60[19]},
      {stage0_61[35]},
      {stage1_62[19],stage1_61[45],stage1_60[75],stage1_59[134],stage1_58[177]}
   );
   gpc1163_5 gpc2280 (
      {stage0_58[272], stage0_58[273], stage0_58[274]},
      {stage0_59[228], stage0_59[229], stage0_59[230], stage0_59[231], stage0_59[232], stage0_59[233]},
      {stage0_60[20]},
      {stage0_61[36]},
      {stage1_62[20],stage1_61[46],stage1_60[76],stage1_59[135],stage1_58[178]}
   );
   gpc1163_5 gpc2281 (
      {stage0_58[275], stage0_58[276], stage0_58[277]},
      {stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238], stage0_59[239]},
      {stage0_60[21]},
      {stage0_61[37]},
      {stage1_62[21],stage1_61[47],stage1_60[77],stage1_59[136],stage1_58[179]}
   );
   gpc1163_5 gpc2282 (
      {stage0_58[278], stage0_58[279], stage0_58[280]},
      {stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[22]},
      {stage0_61[38]},
      {stage1_62[22],stage1_61[48],stage1_60[78],stage1_59[137],stage1_58[180]}
   );
   gpc1163_5 gpc2283 (
      {stage0_58[281], stage0_58[282], stage0_58[283]},
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251]},
      {stage0_60[23]},
      {stage0_61[39]},
      {stage1_62[23],stage1_61[49],stage1_60[79],stage1_59[138],stage1_58[181]}
   );
   gpc1163_5 gpc2284 (
      {stage0_58[284], stage0_58[285], stage0_58[286]},
      {stage0_59[252], stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257]},
      {stage0_60[24]},
      {stage0_61[40]},
      {stage1_62[24],stage1_61[50],stage1_60[80],stage1_59[139],stage1_58[182]}
   );
   gpc1163_5 gpc2285 (
      {stage0_58[287], stage0_58[288], stage0_58[289]},
      {stage0_59[258], stage0_59[259], stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263]},
      {stage0_60[25]},
      {stage0_61[41]},
      {stage1_62[25],stage1_61[51],stage1_60[81],stage1_59[140],stage1_58[183]}
   );
   gpc1163_5 gpc2286 (
      {stage0_58[290], stage0_58[291], stage0_58[292]},
      {stage0_59[264], stage0_59[265], stage0_59[266], stage0_59[267], stage0_59[268], stage0_59[269]},
      {stage0_60[26]},
      {stage0_61[42]},
      {stage1_62[26],stage1_61[52],stage1_60[82],stage1_59[141],stage1_58[184]}
   );
   gpc1163_5 gpc2287 (
      {stage0_58[293], stage0_58[294], stage0_58[295]},
      {stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273], stage0_59[274], stage0_59[275]},
      {stage0_60[27]},
      {stage0_61[43]},
      {stage1_62[27],stage1_61[53],stage1_60[83],stage1_59[142],stage1_58[185]}
   );
   gpc1163_5 gpc2288 (
      {stage0_58[296], stage0_58[297], stage0_58[298]},
      {stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280], stage0_59[281]},
      {stage0_60[28]},
      {stage0_61[44]},
      {stage1_62[28],stage1_61[54],stage1_60[84],stage1_59[143],stage1_58[186]}
   );
   gpc1163_5 gpc2289 (
      {stage0_58[299], stage0_58[300], stage0_58[301]},
      {stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[29]},
      {stage0_61[45]},
      {stage1_62[29],stage1_61[55],stage1_60[85],stage1_59[144],stage1_58[187]}
   );
   gpc1163_5 gpc2290 (
      {stage0_58[302], stage0_58[303], stage0_58[304]},
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293]},
      {stage0_60[30]},
      {stage0_61[46]},
      {stage1_62[30],stage1_61[56],stage1_60[86],stage1_59[145],stage1_58[188]}
   );
   gpc1163_5 gpc2291 (
      {stage0_58[305], stage0_58[306], stage0_58[307]},
      {stage0_59[294], stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299]},
      {stage0_60[31]},
      {stage0_61[47]},
      {stage1_62[31],stage1_61[57],stage1_60[87],stage1_59[146],stage1_58[189]}
   );
   gpc1163_5 gpc2292 (
      {stage0_58[308], stage0_58[309], stage0_58[310]},
      {stage0_59[300], stage0_59[301], stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305]},
      {stage0_60[32]},
      {stage0_61[48]},
      {stage1_62[32],stage1_61[58],stage1_60[88],stage1_59[147],stage1_58[190]}
   );
   gpc1163_5 gpc2293 (
      {stage0_58[311], stage0_58[312], stage0_58[313]},
      {stage0_59[306], stage0_59[307], stage0_59[308], stage0_59[309], stage0_59[310], stage0_59[311]},
      {stage0_60[33]},
      {stage0_61[49]},
      {stage1_62[33],stage1_61[59],stage1_60[89],stage1_59[148],stage1_58[191]}
   );
   gpc1163_5 gpc2294 (
      {stage0_58[314], stage0_58[315], stage0_58[316]},
      {stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315], stage0_59[316], stage0_59[317]},
      {stage0_60[34]},
      {stage0_61[50]},
      {stage1_62[34],stage1_61[60],stage1_60[90],stage1_59[149],stage1_58[192]}
   );
   gpc1163_5 gpc2295 (
      {stage0_58[317], stage0_58[318], stage0_58[319]},
      {stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322], stage0_59[323]},
      {stage0_60[35]},
      {stage0_61[51]},
      {stage1_62[35],stage1_61[61],stage1_60[91],stage1_59[150],stage1_58[193]}
   );
   gpc1163_5 gpc2296 (
      {stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[36]},
      {stage0_61[52]},
      {stage1_62[36],stage1_61[62],stage1_60[92],stage1_59[151],stage1_58[194]}
   );
   gpc606_5 gpc2297 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328]},
      {stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41], stage0_60[42]},
      {stage1_62[37],stage1_61[63],stage1_60[93],stage1_59[152],stage1_58[195]}
   );
   gpc606_5 gpc2298 (
      {stage0_58[329], stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334]},
      {stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47], stage0_60[48]},
      {stage1_62[38],stage1_61[64],stage1_60[94],stage1_59[153],stage1_58[196]}
   );
   gpc606_5 gpc2299 (
      {stage0_58[335], stage0_58[336], stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340]},
      {stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53], stage0_60[54]},
      {stage1_62[39],stage1_61[65],stage1_60[95],stage1_59[154],stage1_58[197]}
   );
   gpc606_5 gpc2300 (
      {stage0_58[341], stage0_58[342], stage0_58[343], stage0_58[344], stage0_58[345], stage0_58[346]},
      {stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59], stage0_60[60]},
      {stage1_62[40],stage1_61[66],stage1_60[96],stage1_59[155],stage1_58[198]}
   );
   gpc606_5 gpc2301 (
      {stage0_58[347], stage0_58[348], stage0_58[349], stage0_58[350], stage0_58[351], stage0_58[352]},
      {stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65], stage0_60[66]},
      {stage1_62[41],stage1_61[67],stage1_60[97],stage1_59[156],stage1_58[199]}
   );
   gpc606_5 gpc2302 (
      {stage0_58[353], stage0_58[354], stage0_58[355], stage0_58[356], stage0_58[357], stage0_58[358]},
      {stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71], stage0_60[72]},
      {stage1_62[42],stage1_61[68],stage1_60[98],stage1_59[157],stage1_58[200]}
   );
   gpc606_5 gpc2303 (
      {stage0_58[359], stage0_58[360], stage0_58[361], stage0_58[362], stage0_58[363], stage0_58[364]},
      {stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77], stage0_60[78]},
      {stage1_62[43],stage1_61[69],stage1_60[99],stage1_59[158],stage1_58[201]}
   );
   gpc606_5 gpc2304 (
      {stage0_58[365], stage0_58[366], stage0_58[367], stage0_58[368], stage0_58[369], stage0_58[370]},
      {stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83], stage0_60[84]},
      {stage1_62[44],stage1_61[70],stage1_60[100],stage1_59[159],stage1_58[202]}
   );
   gpc606_5 gpc2305 (
      {stage0_58[371], stage0_58[372], stage0_58[373], stage0_58[374], stage0_58[375], stage0_58[376]},
      {stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89], stage0_60[90]},
      {stage1_62[45],stage1_61[71],stage1_60[101],stage1_59[160],stage1_58[203]}
   );
   gpc606_5 gpc2306 (
      {stage0_58[377], stage0_58[378], stage0_58[379], stage0_58[380], stage0_58[381], stage0_58[382]},
      {stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95], stage0_60[96]},
      {stage1_62[46],stage1_61[72],stage1_60[102],stage1_59[161],stage1_58[204]}
   );
   gpc606_5 gpc2307 (
      {stage0_58[383], stage0_58[384], stage0_58[385], stage0_58[386], stage0_58[387], stage0_58[388]},
      {stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101], stage0_60[102]},
      {stage1_62[47],stage1_61[73],stage1_60[103],stage1_59[162],stage1_58[205]}
   );
   gpc606_5 gpc2308 (
      {stage0_58[389], stage0_58[390], stage0_58[391], stage0_58[392], stage0_58[393], stage0_58[394]},
      {stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107], stage0_60[108]},
      {stage1_62[48],stage1_61[74],stage1_60[104],stage1_59[163],stage1_58[206]}
   );
   gpc606_5 gpc2309 (
      {stage0_58[395], stage0_58[396], stage0_58[397], stage0_58[398], stage0_58[399], stage0_58[400]},
      {stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113], stage0_60[114]},
      {stage1_62[49],stage1_61[75],stage1_60[105],stage1_59[164],stage1_58[207]}
   );
   gpc606_5 gpc2310 (
      {stage0_58[401], stage0_58[402], stage0_58[403], stage0_58[404], stage0_58[405], stage0_58[406]},
      {stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119], stage0_60[120]},
      {stage1_62[50],stage1_61[76],stage1_60[106],stage1_59[165],stage1_58[208]}
   );
   gpc606_5 gpc2311 (
      {stage0_58[407], stage0_58[408], stage0_58[409], stage0_58[410], stage0_58[411], stage0_58[412]},
      {stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125], stage0_60[126]},
      {stage1_62[51],stage1_61[77],stage1_60[107],stage1_59[166],stage1_58[209]}
   );
   gpc606_5 gpc2312 (
      {stage0_58[413], stage0_58[414], stage0_58[415], stage0_58[416], stage0_58[417], stage0_58[418]},
      {stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131], stage0_60[132]},
      {stage1_62[52],stage1_61[78],stage1_60[108],stage1_59[167],stage1_58[210]}
   );
   gpc606_5 gpc2313 (
      {stage0_58[419], stage0_58[420], stage0_58[421], stage0_58[422], stage0_58[423], stage0_58[424]},
      {stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138]},
      {stage1_62[53],stage1_61[79],stage1_60[109],stage1_59[168],stage1_58[211]}
   );
   gpc606_5 gpc2314 (
      {stage0_58[425], stage0_58[426], stage0_58[427], stage0_58[428], stage0_58[429], stage0_58[430]},
      {stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144]},
      {stage1_62[54],stage1_61[80],stage1_60[110],stage1_59[169],stage1_58[212]}
   );
   gpc606_5 gpc2315 (
      {stage0_58[431], stage0_58[432], stage0_58[433], stage0_58[434], stage0_58[435], stage0_58[436]},
      {stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage1_62[55],stage1_61[81],stage1_60[111],stage1_59[170],stage1_58[213]}
   );
   gpc606_5 gpc2316 (
      {stage0_58[437], stage0_58[438], stage0_58[439], stage0_58[440], stage0_58[441], stage0_58[442]},
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155], stage0_60[156]},
      {stage1_62[56],stage1_61[82],stage1_60[112],stage1_59[171],stage1_58[214]}
   );
   gpc606_5 gpc2317 (
      {stage0_58[443], stage0_58[444], stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448]},
      {stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161], stage0_60[162]},
      {stage1_62[57],stage1_61[83],stage1_60[113],stage1_59[172],stage1_58[215]}
   );
   gpc606_5 gpc2318 (
      {stage0_58[449], stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_60[163], stage0_60[164], stage0_60[165], stage0_60[166], stage0_60[167], stage0_60[168]},
      {stage1_62[58],stage1_61[84],stage1_60[114],stage1_59[173],stage1_58[216]}
   );
   gpc606_5 gpc2319 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459], stage0_58[460]},
      {stage0_60[169], stage0_60[170], stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174]},
      {stage1_62[59],stage1_61[85],stage1_60[115],stage1_59[174],stage1_58[217]}
   );
   gpc606_5 gpc2320 (
      {stage0_58[461], stage0_58[462], stage0_58[463], stage0_58[464], stage0_58[465], stage0_58[466]},
      {stage0_60[175], stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage1_62[60],stage1_61[86],stage1_60[116],stage1_59[175],stage1_58[218]}
   );
   gpc606_5 gpc2321 (
      {stage0_58[467], stage0_58[468], stage0_58[469], stage0_58[470], stage0_58[471], stage0_58[472]},
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185], stage0_60[186]},
      {stage1_62[61],stage1_61[87],stage1_60[117],stage1_59[176],stage1_58[219]}
   );
   gpc615_5 gpc2322 (
      {stage0_58[473], stage0_58[474], stage0_58[475], stage0_58[476], stage0_58[477]},
      {stage0_59[330]},
      {stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190], stage0_60[191], stage0_60[192]},
      {stage1_62[62],stage1_61[88],stage1_60[118],stage1_59[177],stage1_58[220]}
   );
   gpc615_5 gpc2323 (
      {stage0_58[478], stage0_58[479], stage0_58[480], stage0_58[481], stage0_58[482]},
      {stage0_59[331]},
      {stage0_60[193], stage0_60[194], stage0_60[195], stage0_60[196], stage0_60[197], stage0_60[198]},
      {stage1_62[63],stage1_61[89],stage1_60[119],stage1_59[178],stage1_58[221]}
   );
   gpc615_5 gpc2324 (
      {stage0_58[483], stage0_58[484], stage0_58[485], stage0_58[486], stage0_58[487]},
      {stage0_59[332]},
      {stage0_60[199], stage0_60[200], stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204]},
      {stage1_62[64],stage1_61[90],stage1_60[120],stage1_59[179],stage1_58[222]}
   );
   gpc615_5 gpc2325 (
      {stage0_58[488], stage0_58[489], stage0_58[490], stage0_58[491], stage0_58[492]},
      {stage0_59[333]},
      {stage0_60[205], stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage1_62[65],stage1_61[91],stage1_60[121],stage1_59[180],stage1_58[223]}
   );
   gpc606_5 gpc2326 (
      {stage0_59[334], stage0_59[335], stage0_59[336], stage0_59[337], stage0_59[338], stage0_59[339]},
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58]},
      {stage1_63[0],stage1_62[66],stage1_61[92],stage1_60[122],stage1_59[181]}
   );
   gpc606_5 gpc2327 (
      {stage0_59[340], stage0_59[341], stage0_59[342], stage0_59[343], stage0_59[344], stage0_59[345]},
      {stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64]},
      {stage1_63[1],stage1_62[67],stage1_61[93],stage1_60[123],stage1_59[182]}
   );
   gpc606_5 gpc2328 (
      {stage0_59[346], stage0_59[347], stage0_59[348], stage0_59[349], stage0_59[350], stage0_59[351]},
      {stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70]},
      {stage1_63[2],stage1_62[68],stage1_61[94],stage1_60[124],stage1_59[183]}
   );
   gpc606_5 gpc2329 (
      {stage0_59[352], stage0_59[353], stage0_59[354], stage0_59[355], stage0_59[356], stage0_59[357]},
      {stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76]},
      {stage1_63[3],stage1_62[69],stage1_61[95],stage1_60[125],stage1_59[184]}
   );
   gpc606_5 gpc2330 (
      {stage0_59[358], stage0_59[359], stage0_59[360], stage0_59[361], stage0_59[362], stage0_59[363]},
      {stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82]},
      {stage1_63[4],stage1_62[70],stage1_61[96],stage1_60[126],stage1_59[185]}
   );
   gpc606_5 gpc2331 (
      {stage0_59[364], stage0_59[365], stage0_59[366], stage0_59[367], stage0_59[368], stage0_59[369]},
      {stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88]},
      {stage1_63[5],stage1_62[71],stage1_61[97],stage1_60[127],stage1_59[186]}
   );
   gpc606_5 gpc2332 (
      {stage0_59[370], stage0_59[371], stage0_59[372], stage0_59[373], stage0_59[374], stage0_59[375]},
      {stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94]},
      {stage1_63[6],stage1_62[72],stage1_61[98],stage1_60[128],stage1_59[187]}
   );
   gpc606_5 gpc2333 (
      {stage0_59[376], stage0_59[377], stage0_59[378], stage0_59[379], stage0_59[380], stage0_59[381]},
      {stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100]},
      {stage1_63[7],stage1_62[73],stage1_61[99],stage1_60[129],stage1_59[188]}
   );
   gpc606_5 gpc2334 (
      {stage0_59[382], stage0_59[383], stage0_59[384], stage0_59[385], stage0_59[386], stage0_59[387]},
      {stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106]},
      {stage1_63[8],stage1_62[74],stage1_61[100],stage1_60[130],stage1_59[189]}
   );
   gpc606_5 gpc2335 (
      {stage0_59[388], stage0_59[389], stage0_59[390], stage0_59[391], stage0_59[392], stage0_59[393]},
      {stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112]},
      {stage1_63[9],stage1_62[75],stage1_61[101],stage1_60[131],stage1_59[190]}
   );
   gpc606_5 gpc2336 (
      {stage0_59[394], stage0_59[395], stage0_59[396], stage0_59[397], stage0_59[398], stage0_59[399]},
      {stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118]},
      {stage1_63[10],stage1_62[76],stage1_61[102],stage1_60[132],stage1_59[191]}
   );
   gpc606_5 gpc2337 (
      {stage0_59[400], stage0_59[401], stage0_59[402], stage0_59[403], stage0_59[404], stage0_59[405]},
      {stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124]},
      {stage1_63[11],stage1_62[77],stage1_61[103],stage1_60[133],stage1_59[192]}
   );
   gpc606_5 gpc2338 (
      {stage0_59[406], stage0_59[407], stage0_59[408], stage0_59[409], stage0_59[410], stage0_59[411]},
      {stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130]},
      {stage1_63[12],stage1_62[78],stage1_61[104],stage1_60[134],stage1_59[193]}
   );
   gpc606_5 gpc2339 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215], stage0_60[216]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[13],stage1_62[79],stage1_61[105],stage1_60[135]}
   );
   gpc606_5 gpc2340 (
      {stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220], stage0_60[221], stage0_60[222]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[14],stage1_62[80],stage1_61[106],stage1_60[136]}
   );
   gpc606_5 gpc2341 (
      {stage0_60[223], stage0_60[224], stage0_60[225], stage0_60[226], stage0_60[227], stage0_60[228]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[15],stage1_62[81],stage1_61[107],stage1_60[137]}
   );
   gpc606_5 gpc2342 (
      {stage0_60[229], stage0_60[230], stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[16],stage1_62[82],stage1_61[108],stage1_60[138]}
   );
   gpc606_5 gpc2343 (
      {stage0_60[235], stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[17],stage1_62[83],stage1_61[109],stage1_60[139]}
   );
   gpc606_5 gpc2344 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245], stage0_60[246]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[18],stage1_62[84],stage1_61[110],stage1_60[140]}
   );
   gpc606_5 gpc2345 (
      {stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250], stage0_60[251], stage0_60[252]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[19],stage1_62[85],stage1_61[111],stage1_60[141]}
   );
   gpc606_5 gpc2346 (
      {stage0_60[253], stage0_60[254], stage0_60[255], stage0_60[256], stage0_60[257], stage0_60[258]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[20],stage1_62[86],stage1_61[112],stage1_60[142]}
   );
   gpc606_5 gpc2347 (
      {stage0_60[259], stage0_60[260], stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[21],stage1_62[87],stage1_61[113],stage1_60[143]}
   );
   gpc606_5 gpc2348 (
      {stage0_60[265], stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[22],stage1_62[88],stage1_61[114],stage1_60[144]}
   );
   gpc606_5 gpc2349 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275], stage0_60[276]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[23],stage1_62[89],stage1_61[115],stage1_60[145]}
   );
   gpc606_5 gpc2350 (
      {stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280], stage0_60[281], stage0_60[282]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[24],stage1_62[90],stage1_61[116],stage1_60[146]}
   );
   gpc606_5 gpc2351 (
      {stage0_60[283], stage0_60[284], stage0_60[285], stage0_60[286], stage0_60[287], stage0_60[288]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[25],stage1_62[91],stage1_61[117],stage1_60[147]}
   );
   gpc606_5 gpc2352 (
      {stage0_60[289], stage0_60[290], stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[26],stage1_62[92],stage1_61[118],stage1_60[148]}
   );
   gpc606_5 gpc2353 (
      {stage0_60[295], stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[27],stage1_62[93],stage1_61[119],stage1_60[149]}
   );
   gpc606_5 gpc2354 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305], stage0_60[306]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[28],stage1_62[94],stage1_61[120],stage1_60[150]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310], stage0_60[311]},
      {stage0_61[131]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[29],stage1_62[95],stage1_61[121],stage1_60[151]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315], stage0_60[316]},
      {stage0_61[132]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[30],stage1_62[96],stage1_61[122],stage1_60[152]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320], stage0_60[321]},
      {stage0_61[133]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[31],stage1_62[97],stage1_61[123],stage1_60[153]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325], stage0_60[326]},
      {stage0_61[134]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[32],stage1_62[98],stage1_61[124],stage1_60[154]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330], stage0_60[331]},
      {stage0_61[135]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[33],stage1_62[99],stage1_61[125],stage1_60[155]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335], stage0_60[336]},
      {stage0_61[136]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[34],stage1_62[100],stage1_61[126],stage1_60[156]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340], stage0_60[341]},
      {stage0_61[137]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[35],stage1_62[101],stage1_61[127],stage1_60[157]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345], stage0_60[346]},
      {stage0_61[138]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[36],stage1_62[102],stage1_61[128],stage1_60[158]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350], stage0_60[351]},
      {stage0_61[139]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[37],stage1_62[103],stage1_61[129],stage1_60[159]}
   );
   gpc615_5 gpc2364 (
      {stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355], stage0_60[356]},
      {stage0_61[140]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[38],stage1_62[104],stage1_61[130],stage1_60[160]}
   );
   gpc615_5 gpc2365 (
      {stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360], stage0_60[361]},
      {stage0_61[141]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[39],stage1_62[105],stage1_61[131],stage1_60[161]}
   );
   gpc615_5 gpc2366 (
      {stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365], stage0_60[366]},
      {stage0_61[142]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[40],stage1_62[106],stage1_61[132],stage1_60[162]}
   );
   gpc615_5 gpc2367 (
      {stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370], stage0_60[371]},
      {stage0_61[143]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[41],stage1_62[107],stage1_61[133],stage1_60[163]}
   );
   gpc615_5 gpc2368 (
      {stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375], stage0_60[376]},
      {stage0_61[144]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[42],stage1_62[108],stage1_61[134],stage1_60[164]}
   );
   gpc615_5 gpc2369 (
      {stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380], stage0_60[381]},
      {stage0_61[145]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[43],stage1_62[109],stage1_61[135],stage1_60[165]}
   );
   gpc615_5 gpc2370 (
      {stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385], stage0_60[386]},
      {stage0_61[146]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[44],stage1_62[110],stage1_61[136],stage1_60[166]}
   );
   gpc615_5 gpc2371 (
      {stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390], stage0_60[391]},
      {stage0_61[147]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[45],stage1_62[111],stage1_61[137],stage1_60[167]}
   );
   gpc615_5 gpc2372 (
      {stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395], stage0_60[396]},
      {stage0_61[148]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[46],stage1_62[112],stage1_61[138],stage1_60[168]}
   );
   gpc615_5 gpc2373 (
      {stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400], stage0_60[401]},
      {stage0_61[149]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[47],stage1_62[113],stage1_61[139],stage1_60[169]}
   );
   gpc615_5 gpc2374 (
      {stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405], stage0_60[406]},
      {stage0_61[150]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[48],stage1_62[114],stage1_61[140],stage1_60[170]}
   );
   gpc615_5 gpc2375 (
      {stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410], stage0_60[411]},
      {stage0_61[151]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[49],stage1_62[115],stage1_61[141],stage1_60[171]}
   );
   gpc615_5 gpc2376 (
      {stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415], stage0_60[416]},
      {stage0_61[152]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[50],stage1_62[116],stage1_61[142],stage1_60[172]}
   );
   gpc615_5 gpc2377 (
      {stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420], stage0_60[421]},
      {stage0_61[153]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[51],stage1_62[117],stage1_61[143],stage1_60[173]}
   );
   gpc615_5 gpc2378 (
      {stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425], stage0_60[426]},
      {stage0_61[154]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[52],stage1_62[118],stage1_61[144],stage1_60[174]}
   );
   gpc615_5 gpc2379 (
      {stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430], stage0_60[431]},
      {stage0_61[155]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[53],stage1_62[119],stage1_61[145],stage1_60[175]}
   );
   gpc615_5 gpc2380 (
      {stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435], stage0_60[436]},
      {stage0_61[156]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[54],stage1_62[120],stage1_61[146],stage1_60[176]}
   );
   gpc615_5 gpc2381 (
      {stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440], stage0_60[441]},
      {stage0_61[157]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[55],stage1_62[121],stage1_61[147],stage1_60[177]}
   );
   gpc615_5 gpc2382 (
      {stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445], stage0_60[446]},
      {stage0_61[158]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[56],stage1_62[122],stage1_61[148],stage1_60[178]}
   );
   gpc615_5 gpc2383 (
      {stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450], stage0_60[451]},
      {stage0_61[159]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[57],stage1_62[123],stage1_61[149],stage1_60[179]}
   );
   gpc615_5 gpc2384 (
      {stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455], stage0_60[456]},
      {stage0_61[160]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[58],stage1_62[124],stage1_61[150],stage1_60[180]}
   );
   gpc615_5 gpc2385 (
      {stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460], stage0_60[461]},
      {stage0_61[161]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[59],stage1_62[125],stage1_61[151],stage1_60[181]}
   );
   gpc615_5 gpc2386 (
      {stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465], stage0_60[466]},
      {stage0_61[162]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[60],stage1_62[126],stage1_61[152],stage1_60[182]}
   );
   gpc615_5 gpc2387 (
      {stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470], stage0_60[471]},
      {stage0_61[163]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[61],stage1_62[127],stage1_61[153],stage1_60[183]}
   );
   gpc615_5 gpc2388 (
      {stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475], stage0_60[476]},
      {stage0_61[164]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[62],stage1_62[128],stage1_61[154],stage1_60[184]}
   );
   gpc615_5 gpc2389 (
      {stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480], stage0_60[481]},
      {stage0_61[165]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[63],stage1_62[129],stage1_61[155],stage1_60[185]}
   );
   gpc615_5 gpc2390 (
      {stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485], stage0_60[486]},
      {stage0_61[166]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[64],stage1_62[130],stage1_61[156],stage1_60[186]}
   );
   gpc615_5 gpc2391 (
      {stage0_60[487], stage0_60[488], stage0_60[489], stage0_60[490], stage0_60[491]},
      {stage0_61[167]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[65],stage1_62[131],stage1_61[157],stage1_60[187]}
   );
   gpc615_5 gpc2392 (
      {stage0_60[492], stage0_60[493], stage0_60[494], stage0_60[495], stage0_60[496]},
      {stage0_61[168]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[66],stage1_62[132],stage1_61[158],stage1_60[188]}
   );
   gpc615_5 gpc2393 (
      {stage0_60[497], stage0_60[498], stage0_60[499], stage0_60[500], stage0_60[501]},
      {stage0_61[169]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[67],stage1_62[133],stage1_61[159],stage1_60[189]}
   );
   gpc606_5 gpc2394 (
      {stage0_61[170], stage0_61[171], stage0_61[172], stage0_61[173], stage0_61[174], stage0_61[175]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[55],stage1_63[68],stage1_62[134],stage1_61[160]}
   );
   gpc606_5 gpc2395 (
      {stage0_61[176], stage0_61[177], stage0_61[178], stage0_61[179], stage0_61[180], stage0_61[181]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[56],stage1_63[69],stage1_62[135],stage1_61[161]}
   );
   gpc606_5 gpc2396 (
      {stage0_61[182], stage0_61[183], stage0_61[184], stage0_61[185], stage0_61[186], stage0_61[187]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[57],stage1_63[70],stage1_62[136],stage1_61[162]}
   );
   gpc606_5 gpc2397 (
      {stage0_61[188], stage0_61[189], stage0_61[190], stage0_61[191], stage0_61[192], stage0_61[193]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[58],stage1_63[71],stage1_62[137],stage1_61[163]}
   );
   gpc606_5 gpc2398 (
      {stage0_61[194], stage0_61[195], stage0_61[196], stage0_61[197], stage0_61[198], stage0_61[199]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[59],stage1_63[72],stage1_62[138],stage1_61[164]}
   );
   gpc606_5 gpc2399 (
      {stage0_61[200], stage0_61[201], stage0_61[202], stage0_61[203], stage0_61[204], stage0_61[205]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[60],stage1_63[73],stage1_62[139],stage1_61[165]}
   );
   gpc606_5 gpc2400 (
      {stage0_61[206], stage0_61[207], stage0_61[208], stage0_61[209], stage0_61[210], stage0_61[211]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[61],stage1_63[74],stage1_62[140],stage1_61[166]}
   );
   gpc606_5 gpc2401 (
      {stage0_61[212], stage0_61[213], stage0_61[214], stage0_61[215], stage0_61[216], stage0_61[217]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[62],stage1_63[75],stage1_62[141],stage1_61[167]}
   );
   gpc606_5 gpc2402 (
      {stage0_61[218], stage0_61[219], stage0_61[220], stage0_61[221], stage0_61[222], stage0_61[223]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[63],stage1_63[76],stage1_62[142],stage1_61[168]}
   );
   gpc606_5 gpc2403 (
      {stage0_61[224], stage0_61[225], stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[64],stage1_63[77],stage1_62[143],stage1_61[169]}
   );
   gpc606_5 gpc2404 (
      {stage0_61[230], stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[65],stage1_63[78],stage1_62[144],stage1_61[170]}
   );
   gpc606_5 gpc2405 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240], stage0_61[241]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[66],stage1_63[79],stage1_62[145],stage1_61[171]}
   );
   gpc606_5 gpc2406 (
      {stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245], stage0_61[246], stage0_61[247]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[67],stage1_63[80],stage1_62[146],stage1_61[172]}
   );
   gpc606_5 gpc2407 (
      {stage0_61[248], stage0_61[249], stage0_61[250], stage0_61[251], stage0_61[252], stage0_61[253]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[68],stage1_63[81],stage1_62[147],stage1_61[173]}
   );
   gpc606_5 gpc2408 (
      {stage0_61[254], stage0_61[255], stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[69],stage1_63[82],stage1_62[148],stage1_61[174]}
   );
   gpc606_5 gpc2409 (
      {stage0_61[260], stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[70],stage1_63[83],stage1_62[149],stage1_61[175]}
   );
   gpc606_5 gpc2410 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270], stage0_61[271]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[71],stage1_63[84],stage1_62[150],stage1_61[176]}
   );
   gpc606_5 gpc2411 (
      {stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275], stage0_61[276], stage0_61[277]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[72],stage1_63[85],stage1_62[151],stage1_61[177]}
   );
   gpc606_5 gpc2412 (
      {stage0_61[278], stage0_61[279], stage0_61[280], stage0_61[281], stage0_61[282], stage0_61[283]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[73],stage1_63[86],stage1_62[152],stage1_61[178]}
   );
   gpc606_5 gpc2413 (
      {stage0_61[284], stage0_61[285], stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[74],stage1_63[87],stage1_62[153],stage1_61[179]}
   );
   gpc606_5 gpc2414 (
      {stage0_61[290], stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[75],stage1_63[88],stage1_62[154],stage1_61[180]}
   );
   gpc606_5 gpc2415 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300], stage0_61[301]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[76],stage1_63[89],stage1_62[155],stage1_61[181]}
   );
   gpc606_5 gpc2416 (
      {stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305], stage0_61[306], stage0_61[307]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[77],stage1_63[90],stage1_62[156],stage1_61[182]}
   );
   gpc606_5 gpc2417 (
      {stage0_61[308], stage0_61[309], stage0_61[310], stage0_61[311], stage0_61[312], stage0_61[313]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[78],stage1_63[91],stage1_62[157],stage1_61[183]}
   );
   gpc606_5 gpc2418 (
      {stage0_61[314], stage0_61[315], stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[79],stage1_63[92],stage1_62[158],stage1_61[184]}
   );
   gpc606_5 gpc2419 (
      {stage0_61[320], stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[80],stage1_63[93],stage1_62[159],stage1_61[185]}
   );
   gpc606_5 gpc2420 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330], stage0_61[331]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[81],stage1_63[94],stage1_62[160],stage1_61[186]}
   );
   gpc606_5 gpc2421 (
      {stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335], stage0_61[336], stage0_61[337]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[82],stage1_63[95],stage1_62[161],stage1_61[187]}
   );
   gpc606_5 gpc2422 (
      {stage0_61[338], stage0_61[339], stage0_61[340], stage0_61[341], stage0_61[342], stage0_61[343]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[83],stage1_63[96],stage1_62[162],stage1_61[188]}
   );
   gpc606_5 gpc2423 (
      {stage0_61[344], stage0_61[345], stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[84],stage1_63[97],stage1_62[163],stage1_61[189]}
   );
   gpc606_5 gpc2424 (
      {stage0_61[350], stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[85],stage1_63[98],stage1_62[164],stage1_61[190]}
   );
   gpc606_5 gpc2425 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360], stage0_61[361]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[86],stage1_63[99],stage1_62[165],stage1_61[191]}
   );
   gpc606_5 gpc2426 (
      {stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365], stage0_61[366], stage0_61[367]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[87],stage1_63[100],stage1_62[166],stage1_61[192]}
   );
   gpc606_5 gpc2427 (
      {stage0_61[368], stage0_61[369], stage0_61[370], stage0_61[371], stage0_61[372], stage0_61[373]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[88],stage1_63[101],stage1_62[167],stage1_61[193]}
   );
   gpc606_5 gpc2428 (
      {stage0_61[374], stage0_61[375], stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[89],stage1_63[102],stage1_62[168],stage1_61[194]}
   );
   gpc606_5 gpc2429 (
      {stage0_61[380], stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[90],stage1_63[103],stage1_62[169],stage1_61[195]}
   );
   gpc606_5 gpc2430 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390], stage0_61[391]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[91],stage1_63[104],stage1_62[170],stage1_61[196]}
   );
   gpc606_5 gpc2431 (
      {stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395], stage0_61[396], stage0_61[397]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[92],stage1_63[105],stage1_62[171],stage1_61[197]}
   );
   gpc606_5 gpc2432 (
      {stage0_61[398], stage0_61[399], stage0_61[400], stage0_61[401], stage0_61[402], stage0_61[403]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[93],stage1_63[106],stage1_62[172],stage1_61[198]}
   );
   gpc606_5 gpc2433 (
      {stage0_61[404], stage0_61[405], stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[94],stage1_63[107],stage1_62[173],stage1_61[199]}
   );
   gpc606_5 gpc2434 (
      {stage0_61[410], stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[95],stage1_63[108],stage1_62[174],stage1_61[200]}
   );
   gpc606_5 gpc2435 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420], stage0_61[421]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[96],stage1_63[109],stage1_62[175],stage1_61[201]}
   );
   gpc606_5 gpc2436 (
      {stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425], stage0_61[426], stage0_61[427]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[97],stage1_63[110],stage1_62[176],stage1_61[202]}
   );
   gpc606_5 gpc2437 (
      {stage0_61[428], stage0_61[429], stage0_61[430], stage0_61[431], stage0_61[432], stage0_61[433]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[98],stage1_63[111],stage1_62[177],stage1_61[203]}
   );
   gpc606_5 gpc2438 (
      {stage0_61[434], stage0_61[435], stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[99],stage1_63[112],stage1_62[178],stage1_61[204]}
   );
   gpc606_5 gpc2439 (
      {stage0_61[440], stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[100],stage1_63[113],stage1_62[179],stage1_61[205]}
   );
   gpc606_5 gpc2440 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450], stage0_61[451]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[101],stage1_63[114],stage1_62[180],stage1_61[206]}
   );
   gpc606_5 gpc2441 (
      {stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455], stage0_61[456], stage0_61[457]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[102],stage1_63[115],stage1_62[181],stage1_61[207]}
   );
   gpc606_5 gpc2442 (
      {stage0_61[458], stage0_61[459], stage0_61[460], stage0_61[461], stage0_61[462], stage0_61[463]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[103],stage1_63[116],stage1_62[182],stage1_61[208]}
   );
   gpc606_5 gpc2443 (
      {stage0_61[464], stage0_61[465], stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[104],stage1_63[117],stage1_62[183],stage1_61[209]}
   );
   gpc606_5 gpc2444 (
      {stage0_61[470], stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[105],stage1_63[118],stage1_62[184],stage1_61[210]}
   );
   gpc606_5 gpc2445 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480], stage0_61[481]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[106],stage1_63[119],stage1_62[185],stage1_61[211]}
   );
   gpc606_5 gpc2446 (
      {stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485], stage0_61[486], stage0_61[487]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[107],stage1_63[120],stage1_62[186],stage1_61[212]}
   );
   gpc606_5 gpc2447 (
      {stage0_61[488], stage0_61[489], stage0_61[490], stage0_61[491], stage0_61[492], stage0_61[493]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[108],stage1_63[121],stage1_62[187],stage1_61[213]}
   );
   gpc606_5 gpc2448 (
      {stage0_61[494], stage0_61[495], stage0_61[496], stage0_61[497], stage0_61[498], stage0_61[499]},
      {stage0_63[324], stage0_63[325], stage0_63[326], stage0_63[327], stage0_63[328], stage0_63[329]},
      {stage1_65[54],stage1_64[109],stage1_63[122],stage1_62[188],stage1_61[214]}
   );
   gpc606_5 gpc2449 (
      {stage0_61[500], stage0_61[501], stage0_61[502], stage0_61[503], stage0_61[504], stage0_61[505]},
      {stage0_63[330], stage0_63[331], stage0_63[332], stage0_63[333], stage0_63[334], stage0_63[335]},
      {stage1_65[55],stage1_64[110],stage1_63[123],stage1_62[189],stage1_61[215]}
   );
   gpc606_5 gpc2450 (
      {stage0_61[506], stage0_61[507], stage0_61[508], stage0_61[509], stage0_61[510], stage0_61[511]},
      {stage0_63[336], stage0_63[337], stage0_63[338], stage0_63[339], stage0_63[340], stage0_63[341]},
      {stage1_65[56],stage1_64[111],stage1_63[124],stage1_62[190],stage1_61[216]}
   );
   gpc1_1 gpc2451 (
      {stage0_1[481]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2452 (
      {stage0_1[482]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2453 (
      {stage0_1[483]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2454 (
      {stage0_1[484]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2455 (
      {stage0_1[485]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[486]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[487]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[488]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[489]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[490]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[491]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[492]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[493]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[494]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[495]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[496]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[497]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[498]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[499]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[500]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[501]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[502]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[503]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[504]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[505]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[506]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[507]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[508]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[509]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[510]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[511]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2482 (
      {stage0_2[429]},
      {stage1_2[138]}
   );
   gpc1_1 gpc2483 (
      {stage0_2[430]},
      {stage1_2[139]}
   );
   gpc1_1 gpc2484 (
      {stage0_2[431]},
      {stage1_2[140]}
   );
   gpc1_1 gpc2485 (
      {stage0_2[432]},
      {stage1_2[141]}
   );
   gpc1_1 gpc2486 (
      {stage0_2[433]},
      {stage1_2[142]}
   );
   gpc1_1 gpc2487 (
      {stage0_2[434]},
      {stage1_2[143]}
   );
   gpc1_1 gpc2488 (
      {stage0_2[435]},
      {stage1_2[144]}
   );
   gpc1_1 gpc2489 (
      {stage0_2[436]},
      {stage1_2[145]}
   );
   gpc1_1 gpc2490 (
      {stage0_2[437]},
      {stage1_2[146]}
   );
   gpc1_1 gpc2491 (
      {stage0_2[438]},
      {stage1_2[147]}
   );
   gpc1_1 gpc2492 (
      {stage0_2[439]},
      {stage1_2[148]}
   );
   gpc1_1 gpc2493 (
      {stage0_2[440]},
      {stage1_2[149]}
   );
   gpc1_1 gpc2494 (
      {stage0_2[441]},
      {stage1_2[150]}
   );
   gpc1_1 gpc2495 (
      {stage0_2[442]},
      {stage1_2[151]}
   );
   gpc1_1 gpc2496 (
      {stage0_2[443]},
      {stage1_2[152]}
   );
   gpc1_1 gpc2497 (
      {stage0_2[444]},
      {stage1_2[153]}
   );
   gpc1_1 gpc2498 (
      {stage0_2[445]},
      {stage1_2[154]}
   );
   gpc1_1 gpc2499 (
      {stage0_2[446]},
      {stage1_2[155]}
   );
   gpc1_1 gpc2500 (
      {stage0_2[447]},
      {stage1_2[156]}
   );
   gpc1_1 gpc2501 (
      {stage0_2[448]},
      {stage1_2[157]}
   );
   gpc1_1 gpc2502 (
      {stage0_2[449]},
      {stage1_2[158]}
   );
   gpc1_1 gpc2503 (
      {stage0_2[450]},
      {stage1_2[159]}
   );
   gpc1_1 gpc2504 (
      {stage0_2[451]},
      {stage1_2[160]}
   );
   gpc1_1 gpc2505 (
      {stage0_2[452]},
      {stage1_2[161]}
   );
   gpc1_1 gpc2506 (
      {stage0_2[453]},
      {stage1_2[162]}
   );
   gpc1_1 gpc2507 (
      {stage0_2[454]},
      {stage1_2[163]}
   );
   gpc1_1 gpc2508 (
      {stage0_2[455]},
      {stage1_2[164]}
   );
   gpc1_1 gpc2509 (
      {stage0_2[456]},
      {stage1_2[165]}
   );
   gpc1_1 gpc2510 (
      {stage0_2[457]},
      {stage1_2[166]}
   );
   gpc1_1 gpc2511 (
      {stage0_2[458]},
      {stage1_2[167]}
   );
   gpc1_1 gpc2512 (
      {stage0_2[459]},
      {stage1_2[168]}
   );
   gpc1_1 gpc2513 (
      {stage0_2[460]},
      {stage1_2[169]}
   );
   gpc1_1 gpc2514 (
      {stage0_2[461]},
      {stage1_2[170]}
   );
   gpc1_1 gpc2515 (
      {stage0_2[462]},
      {stage1_2[171]}
   );
   gpc1_1 gpc2516 (
      {stage0_2[463]},
      {stage1_2[172]}
   );
   gpc1_1 gpc2517 (
      {stage0_2[464]},
      {stage1_2[173]}
   );
   gpc1_1 gpc2518 (
      {stage0_2[465]},
      {stage1_2[174]}
   );
   gpc1_1 gpc2519 (
      {stage0_2[466]},
      {stage1_2[175]}
   );
   gpc1_1 gpc2520 (
      {stage0_2[467]},
      {stage1_2[176]}
   );
   gpc1_1 gpc2521 (
      {stage0_2[468]},
      {stage1_2[177]}
   );
   gpc1_1 gpc2522 (
      {stage0_2[469]},
      {stage1_2[178]}
   );
   gpc1_1 gpc2523 (
      {stage0_2[470]},
      {stage1_2[179]}
   );
   gpc1_1 gpc2524 (
      {stage0_2[471]},
      {stage1_2[180]}
   );
   gpc1_1 gpc2525 (
      {stage0_2[472]},
      {stage1_2[181]}
   );
   gpc1_1 gpc2526 (
      {stage0_2[473]},
      {stage1_2[182]}
   );
   gpc1_1 gpc2527 (
      {stage0_2[474]},
      {stage1_2[183]}
   );
   gpc1_1 gpc2528 (
      {stage0_2[475]},
      {stage1_2[184]}
   );
   gpc1_1 gpc2529 (
      {stage0_2[476]},
      {stage1_2[185]}
   );
   gpc1_1 gpc2530 (
      {stage0_2[477]},
      {stage1_2[186]}
   );
   gpc1_1 gpc2531 (
      {stage0_2[478]},
      {stage1_2[187]}
   );
   gpc1_1 gpc2532 (
      {stage0_2[479]},
      {stage1_2[188]}
   );
   gpc1_1 gpc2533 (
      {stage0_2[480]},
      {stage1_2[189]}
   );
   gpc1_1 gpc2534 (
      {stage0_2[481]},
      {stage1_2[190]}
   );
   gpc1_1 gpc2535 (
      {stage0_2[482]},
      {stage1_2[191]}
   );
   gpc1_1 gpc2536 (
      {stage0_2[483]},
      {stage1_2[192]}
   );
   gpc1_1 gpc2537 (
      {stage0_2[484]},
      {stage1_2[193]}
   );
   gpc1_1 gpc2538 (
      {stage0_2[485]},
      {stage1_2[194]}
   );
   gpc1_1 gpc2539 (
      {stage0_2[486]},
      {stage1_2[195]}
   );
   gpc1_1 gpc2540 (
      {stage0_2[487]},
      {stage1_2[196]}
   );
   gpc1_1 gpc2541 (
      {stage0_2[488]},
      {stage1_2[197]}
   );
   gpc1_1 gpc2542 (
      {stage0_2[489]},
      {stage1_2[198]}
   );
   gpc1_1 gpc2543 (
      {stage0_2[490]},
      {stage1_2[199]}
   );
   gpc1_1 gpc2544 (
      {stage0_2[491]},
      {stage1_2[200]}
   );
   gpc1_1 gpc2545 (
      {stage0_2[492]},
      {stage1_2[201]}
   );
   gpc1_1 gpc2546 (
      {stage0_2[493]},
      {stage1_2[202]}
   );
   gpc1_1 gpc2547 (
      {stage0_2[494]},
      {stage1_2[203]}
   );
   gpc1_1 gpc2548 (
      {stage0_2[495]},
      {stage1_2[204]}
   );
   gpc1_1 gpc2549 (
      {stage0_2[496]},
      {stage1_2[205]}
   );
   gpc1_1 gpc2550 (
      {stage0_2[497]},
      {stage1_2[206]}
   );
   gpc1_1 gpc2551 (
      {stage0_2[498]},
      {stage1_2[207]}
   );
   gpc1_1 gpc2552 (
      {stage0_2[499]},
      {stage1_2[208]}
   );
   gpc1_1 gpc2553 (
      {stage0_2[500]},
      {stage1_2[209]}
   );
   gpc1_1 gpc2554 (
      {stage0_2[501]},
      {stage1_2[210]}
   );
   gpc1_1 gpc2555 (
      {stage0_2[502]},
      {stage1_2[211]}
   );
   gpc1_1 gpc2556 (
      {stage0_2[503]},
      {stage1_2[212]}
   );
   gpc1_1 gpc2557 (
      {stage0_2[504]},
      {stage1_2[213]}
   );
   gpc1_1 gpc2558 (
      {stage0_2[505]},
      {stage1_2[214]}
   );
   gpc1_1 gpc2559 (
      {stage0_2[506]},
      {stage1_2[215]}
   );
   gpc1_1 gpc2560 (
      {stage0_2[507]},
      {stage1_2[216]}
   );
   gpc1_1 gpc2561 (
      {stage0_2[508]},
      {stage1_2[217]}
   );
   gpc1_1 gpc2562 (
      {stage0_2[509]},
      {stage1_2[218]}
   );
   gpc1_1 gpc2563 (
      {stage0_2[510]},
      {stage1_2[219]}
   );
   gpc1_1 gpc2564 (
      {stage0_2[511]},
      {stage1_2[220]}
   );
   gpc1_1 gpc2565 (
      {stage0_3[372]},
      {stage1_3[182]}
   );
   gpc1_1 gpc2566 (
      {stage0_3[373]},
      {stage1_3[183]}
   );
   gpc1_1 gpc2567 (
      {stage0_3[374]},
      {stage1_3[184]}
   );
   gpc1_1 gpc2568 (
      {stage0_3[375]},
      {stage1_3[185]}
   );
   gpc1_1 gpc2569 (
      {stage0_3[376]},
      {stage1_3[186]}
   );
   gpc1_1 gpc2570 (
      {stage0_3[377]},
      {stage1_3[187]}
   );
   gpc1_1 gpc2571 (
      {stage0_3[378]},
      {stage1_3[188]}
   );
   gpc1_1 gpc2572 (
      {stage0_3[379]},
      {stage1_3[189]}
   );
   gpc1_1 gpc2573 (
      {stage0_3[380]},
      {stage1_3[190]}
   );
   gpc1_1 gpc2574 (
      {stage0_3[381]},
      {stage1_3[191]}
   );
   gpc1_1 gpc2575 (
      {stage0_3[382]},
      {stage1_3[192]}
   );
   gpc1_1 gpc2576 (
      {stage0_3[383]},
      {stage1_3[193]}
   );
   gpc1_1 gpc2577 (
      {stage0_3[384]},
      {stage1_3[194]}
   );
   gpc1_1 gpc2578 (
      {stage0_3[385]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2579 (
      {stage0_3[386]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2580 (
      {stage0_3[387]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2581 (
      {stage0_3[388]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2582 (
      {stage0_3[389]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2583 (
      {stage0_3[390]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2584 (
      {stage0_3[391]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2585 (
      {stage0_3[392]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2586 (
      {stage0_3[393]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2587 (
      {stage0_3[394]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2588 (
      {stage0_3[395]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2589 (
      {stage0_3[396]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2590 (
      {stage0_3[397]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2591 (
      {stage0_3[398]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2592 (
      {stage0_3[399]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2593 (
      {stage0_3[400]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2594 (
      {stage0_3[401]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2595 (
      {stage0_3[402]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2596 (
      {stage0_3[403]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2597 (
      {stage0_3[404]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2598 (
      {stage0_3[405]},
      {stage1_3[215]}
   );
   gpc1_1 gpc2599 (
      {stage0_3[406]},
      {stage1_3[216]}
   );
   gpc1_1 gpc2600 (
      {stage0_3[407]},
      {stage1_3[217]}
   );
   gpc1_1 gpc2601 (
      {stage0_3[408]},
      {stage1_3[218]}
   );
   gpc1_1 gpc2602 (
      {stage0_3[409]},
      {stage1_3[219]}
   );
   gpc1_1 gpc2603 (
      {stage0_3[410]},
      {stage1_3[220]}
   );
   gpc1_1 gpc2604 (
      {stage0_3[411]},
      {stage1_3[221]}
   );
   gpc1_1 gpc2605 (
      {stage0_3[412]},
      {stage1_3[222]}
   );
   gpc1_1 gpc2606 (
      {stage0_3[413]},
      {stage1_3[223]}
   );
   gpc1_1 gpc2607 (
      {stage0_3[414]},
      {stage1_3[224]}
   );
   gpc1_1 gpc2608 (
      {stage0_3[415]},
      {stage1_3[225]}
   );
   gpc1_1 gpc2609 (
      {stage0_3[416]},
      {stage1_3[226]}
   );
   gpc1_1 gpc2610 (
      {stage0_3[417]},
      {stage1_3[227]}
   );
   gpc1_1 gpc2611 (
      {stage0_3[418]},
      {stage1_3[228]}
   );
   gpc1_1 gpc2612 (
      {stage0_3[419]},
      {stage1_3[229]}
   );
   gpc1_1 gpc2613 (
      {stage0_3[420]},
      {stage1_3[230]}
   );
   gpc1_1 gpc2614 (
      {stage0_3[421]},
      {stage1_3[231]}
   );
   gpc1_1 gpc2615 (
      {stage0_3[422]},
      {stage1_3[232]}
   );
   gpc1_1 gpc2616 (
      {stage0_3[423]},
      {stage1_3[233]}
   );
   gpc1_1 gpc2617 (
      {stage0_3[424]},
      {stage1_3[234]}
   );
   gpc1_1 gpc2618 (
      {stage0_3[425]},
      {stage1_3[235]}
   );
   gpc1_1 gpc2619 (
      {stage0_3[426]},
      {stage1_3[236]}
   );
   gpc1_1 gpc2620 (
      {stage0_3[427]},
      {stage1_3[237]}
   );
   gpc1_1 gpc2621 (
      {stage0_3[428]},
      {stage1_3[238]}
   );
   gpc1_1 gpc2622 (
      {stage0_3[429]},
      {stage1_3[239]}
   );
   gpc1_1 gpc2623 (
      {stage0_3[430]},
      {stage1_3[240]}
   );
   gpc1_1 gpc2624 (
      {stage0_3[431]},
      {stage1_3[241]}
   );
   gpc1_1 gpc2625 (
      {stage0_3[432]},
      {stage1_3[242]}
   );
   gpc1_1 gpc2626 (
      {stage0_3[433]},
      {stage1_3[243]}
   );
   gpc1_1 gpc2627 (
      {stage0_3[434]},
      {stage1_3[244]}
   );
   gpc1_1 gpc2628 (
      {stage0_3[435]},
      {stage1_3[245]}
   );
   gpc1_1 gpc2629 (
      {stage0_3[436]},
      {stage1_3[246]}
   );
   gpc1_1 gpc2630 (
      {stage0_3[437]},
      {stage1_3[247]}
   );
   gpc1_1 gpc2631 (
      {stage0_3[438]},
      {stage1_3[248]}
   );
   gpc1_1 gpc2632 (
      {stage0_3[439]},
      {stage1_3[249]}
   );
   gpc1_1 gpc2633 (
      {stage0_3[440]},
      {stage1_3[250]}
   );
   gpc1_1 gpc2634 (
      {stage0_3[441]},
      {stage1_3[251]}
   );
   gpc1_1 gpc2635 (
      {stage0_3[442]},
      {stage1_3[252]}
   );
   gpc1_1 gpc2636 (
      {stage0_3[443]},
      {stage1_3[253]}
   );
   gpc1_1 gpc2637 (
      {stage0_3[444]},
      {stage1_3[254]}
   );
   gpc1_1 gpc2638 (
      {stage0_3[445]},
      {stage1_3[255]}
   );
   gpc1_1 gpc2639 (
      {stage0_3[446]},
      {stage1_3[256]}
   );
   gpc1_1 gpc2640 (
      {stage0_3[447]},
      {stage1_3[257]}
   );
   gpc1_1 gpc2641 (
      {stage0_3[448]},
      {stage1_3[258]}
   );
   gpc1_1 gpc2642 (
      {stage0_3[449]},
      {stage1_3[259]}
   );
   gpc1_1 gpc2643 (
      {stage0_3[450]},
      {stage1_3[260]}
   );
   gpc1_1 gpc2644 (
      {stage0_3[451]},
      {stage1_3[261]}
   );
   gpc1_1 gpc2645 (
      {stage0_3[452]},
      {stage1_3[262]}
   );
   gpc1_1 gpc2646 (
      {stage0_3[453]},
      {stage1_3[263]}
   );
   gpc1_1 gpc2647 (
      {stage0_3[454]},
      {stage1_3[264]}
   );
   gpc1_1 gpc2648 (
      {stage0_3[455]},
      {stage1_3[265]}
   );
   gpc1_1 gpc2649 (
      {stage0_3[456]},
      {stage1_3[266]}
   );
   gpc1_1 gpc2650 (
      {stage0_3[457]},
      {stage1_3[267]}
   );
   gpc1_1 gpc2651 (
      {stage0_3[458]},
      {stage1_3[268]}
   );
   gpc1_1 gpc2652 (
      {stage0_3[459]},
      {stage1_3[269]}
   );
   gpc1_1 gpc2653 (
      {stage0_3[460]},
      {stage1_3[270]}
   );
   gpc1_1 gpc2654 (
      {stage0_3[461]},
      {stage1_3[271]}
   );
   gpc1_1 gpc2655 (
      {stage0_3[462]},
      {stage1_3[272]}
   );
   gpc1_1 gpc2656 (
      {stage0_3[463]},
      {stage1_3[273]}
   );
   gpc1_1 gpc2657 (
      {stage0_3[464]},
      {stage1_3[274]}
   );
   gpc1_1 gpc2658 (
      {stage0_3[465]},
      {stage1_3[275]}
   );
   gpc1_1 gpc2659 (
      {stage0_3[466]},
      {stage1_3[276]}
   );
   gpc1_1 gpc2660 (
      {stage0_3[467]},
      {stage1_3[277]}
   );
   gpc1_1 gpc2661 (
      {stage0_3[468]},
      {stage1_3[278]}
   );
   gpc1_1 gpc2662 (
      {stage0_3[469]},
      {stage1_3[279]}
   );
   gpc1_1 gpc2663 (
      {stage0_3[470]},
      {stage1_3[280]}
   );
   gpc1_1 gpc2664 (
      {stage0_3[471]},
      {stage1_3[281]}
   );
   gpc1_1 gpc2665 (
      {stage0_3[472]},
      {stage1_3[282]}
   );
   gpc1_1 gpc2666 (
      {stage0_3[473]},
      {stage1_3[283]}
   );
   gpc1_1 gpc2667 (
      {stage0_3[474]},
      {stage1_3[284]}
   );
   gpc1_1 gpc2668 (
      {stage0_3[475]},
      {stage1_3[285]}
   );
   gpc1_1 gpc2669 (
      {stage0_3[476]},
      {stage1_3[286]}
   );
   gpc1_1 gpc2670 (
      {stage0_3[477]},
      {stage1_3[287]}
   );
   gpc1_1 gpc2671 (
      {stage0_3[478]},
      {stage1_3[288]}
   );
   gpc1_1 gpc2672 (
      {stage0_3[479]},
      {stage1_3[289]}
   );
   gpc1_1 gpc2673 (
      {stage0_3[480]},
      {stage1_3[290]}
   );
   gpc1_1 gpc2674 (
      {stage0_3[481]},
      {stage1_3[291]}
   );
   gpc1_1 gpc2675 (
      {stage0_3[482]},
      {stage1_3[292]}
   );
   gpc1_1 gpc2676 (
      {stage0_3[483]},
      {stage1_3[293]}
   );
   gpc1_1 gpc2677 (
      {stage0_3[484]},
      {stage1_3[294]}
   );
   gpc1_1 gpc2678 (
      {stage0_3[485]},
      {stage1_3[295]}
   );
   gpc1_1 gpc2679 (
      {stage0_3[486]},
      {stage1_3[296]}
   );
   gpc1_1 gpc2680 (
      {stage0_3[487]},
      {stage1_3[297]}
   );
   gpc1_1 gpc2681 (
      {stage0_3[488]},
      {stage1_3[298]}
   );
   gpc1_1 gpc2682 (
      {stage0_3[489]},
      {stage1_3[299]}
   );
   gpc1_1 gpc2683 (
      {stage0_3[490]},
      {stage1_3[300]}
   );
   gpc1_1 gpc2684 (
      {stage0_3[491]},
      {stage1_3[301]}
   );
   gpc1_1 gpc2685 (
      {stage0_3[492]},
      {stage1_3[302]}
   );
   gpc1_1 gpc2686 (
      {stage0_3[493]},
      {stage1_3[303]}
   );
   gpc1_1 gpc2687 (
      {stage0_3[494]},
      {stage1_3[304]}
   );
   gpc1_1 gpc2688 (
      {stage0_3[495]},
      {stage1_3[305]}
   );
   gpc1_1 gpc2689 (
      {stage0_3[496]},
      {stage1_3[306]}
   );
   gpc1_1 gpc2690 (
      {stage0_3[497]},
      {stage1_3[307]}
   );
   gpc1_1 gpc2691 (
      {stage0_3[498]},
      {stage1_3[308]}
   );
   gpc1_1 gpc2692 (
      {stage0_3[499]},
      {stage1_3[309]}
   );
   gpc1_1 gpc2693 (
      {stage0_3[500]},
      {stage1_3[310]}
   );
   gpc1_1 gpc2694 (
      {stage0_3[501]},
      {stage1_3[311]}
   );
   gpc1_1 gpc2695 (
      {stage0_3[502]},
      {stage1_3[312]}
   );
   gpc1_1 gpc2696 (
      {stage0_3[503]},
      {stage1_3[313]}
   );
   gpc1_1 gpc2697 (
      {stage0_3[504]},
      {stage1_3[314]}
   );
   gpc1_1 gpc2698 (
      {stage0_3[505]},
      {stage1_3[315]}
   );
   gpc1_1 gpc2699 (
      {stage0_3[506]},
      {stage1_3[316]}
   );
   gpc1_1 gpc2700 (
      {stage0_3[507]},
      {stage1_3[317]}
   );
   gpc1_1 gpc2701 (
      {stage0_3[508]},
      {stage1_3[318]}
   );
   gpc1_1 gpc2702 (
      {stage0_3[509]},
      {stage1_3[319]}
   );
   gpc1_1 gpc2703 (
      {stage0_3[510]},
      {stage1_3[320]}
   );
   gpc1_1 gpc2704 (
      {stage0_3[511]},
      {stage1_3[321]}
   );
   gpc1_1 gpc2705 (
      {stage0_5[468]},
      {stage1_5[173]}
   );
   gpc1_1 gpc2706 (
      {stage0_5[469]},
      {stage1_5[174]}
   );
   gpc1_1 gpc2707 (
      {stage0_5[470]},
      {stage1_5[175]}
   );
   gpc1_1 gpc2708 (
      {stage0_5[471]},
      {stage1_5[176]}
   );
   gpc1_1 gpc2709 (
      {stage0_5[472]},
      {stage1_5[177]}
   );
   gpc1_1 gpc2710 (
      {stage0_5[473]},
      {stage1_5[178]}
   );
   gpc1_1 gpc2711 (
      {stage0_5[474]},
      {stage1_5[179]}
   );
   gpc1_1 gpc2712 (
      {stage0_5[475]},
      {stage1_5[180]}
   );
   gpc1_1 gpc2713 (
      {stage0_5[476]},
      {stage1_5[181]}
   );
   gpc1_1 gpc2714 (
      {stage0_5[477]},
      {stage1_5[182]}
   );
   gpc1_1 gpc2715 (
      {stage0_5[478]},
      {stage1_5[183]}
   );
   gpc1_1 gpc2716 (
      {stage0_5[479]},
      {stage1_5[184]}
   );
   gpc1_1 gpc2717 (
      {stage0_5[480]},
      {stage1_5[185]}
   );
   gpc1_1 gpc2718 (
      {stage0_5[481]},
      {stage1_5[186]}
   );
   gpc1_1 gpc2719 (
      {stage0_5[482]},
      {stage1_5[187]}
   );
   gpc1_1 gpc2720 (
      {stage0_5[483]},
      {stage1_5[188]}
   );
   gpc1_1 gpc2721 (
      {stage0_5[484]},
      {stage1_5[189]}
   );
   gpc1_1 gpc2722 (
      {stage0_5[485]},
      {stage1_5[190]}
   );
   gpc1_1 gpc2723 (
      {stage0_5[486]},
      {stage1_5[191]}
   );
   gpc1_1 gpc2724 (
      {stage0_5[487]},
      {stage1_5[192]}
   );
   gpc1_1 gpc2725 (
      {stage0_5[488]},
      {stage1_5[193]}
   );
   gpc1_1 gpc2726 (
      {stage0_5[489]},
      {stage1_5[194]}
   );
   gpc1_1 gpc2727 (
      {stage0_5[490]},
      {stage1_5[195]}
   );
   gpc1_1 gpc2728 (
      {stage0_5[491]},
      {stage1_5[196]}
   );
   gpc1_1 gpc2729 (
      {stage0_5[492]},
      {stage1_5[197]}
   );
   gpc1_1 gpc2730 (
      {stage0_5[493]},
      {stage1_5[198]}
   );
   gpc1_1 gpc2731 (
      {stage0_5[494]},
      {stage1_5[199]}
   );
   gpc1_1 gpc2732 (
      {stage0_5[495]},
      {stage1_5[200]}
   );
   gpc1_1 gpc2733 (
      {stage0_5[496]},
      {stage1_5[201]}
   );
   gpc1_1 gpc2734 (
      {stage0_5[497]},
      {stage1_5[202]}
   );
   gpc1_1 gpc2735 (
      {stage0_5[498]},
      {stage1_5[203]}
   );
   gpc1_1 gpc2736 (
      {stage0_5[499]},
      {stage1_5[204]}
   );
   gpc1_1 gpc2737 (
      {stage0_5[500]},
      {stage1_5[205]}
   );
   gpc1_1 gpc2738 (
      {stage0_5[501]},
      {stage1_5[206]}
   );
   gpc1_1 gpc2739 (
      {stage0_5[502]},
      {stage1_5[207]}
   );
   gpc1_1 gpc2740 (
      {stage0_5[503]},
      {stage1_5[208]}
   );
   gpc1_1 gpc2741 (
      {stage0_5[504]},
      {stage1_5[209]}
   );
   gpc1_1 gpc2742 (
      {stage0_5[505]},
      {stage1_5[210]}
   );
   gpc1_1 gpc2743 (
      {stage0_5[506]},
      {stage1_5[211]}
   );
   gpc1_1 gpc2744 (
      {stage0_5[507]},
      {stage1_5[212]}
   );
   gpc1_1 gpc2745 (
      {stage0_5[508]},
      {stage1_5[213]}
   );
   gpc1_1 gpc2746 (
      {stage0_5[509]},
      {stage1_5[214]}
   );
   gpc1_1 gpc2747 (
      {stage0_5[510]},
      {stage1_5[215]}
   );
   gpc1_1 gpc2748 (
      {stage0_5[511]},
      {stage1_5[216]}
   );
   gpc1_1 gpc2749 (
      {stage0_6[493]},
      {stage1_6[161]}
   );
   gpc1_1 gpc2750 (
      {stage0_6[494]},
      {stage1_6[162]}
   );
   gpc1_1 gpc2751 (
      {stage0_6[495]},
      {stage1_6[163]}
   );
   gpc1_1 gpc2752 (
      {stage0_6[496]},
      {stage1_6[164]}
   );
   gpc1_1 gpc2753 (
      {stage0_6[497]},
      {stage1_6[165]}
   );
   gpc1_1 gpc2754 (
      {stage0_6[498]},
      {stage1_6[166]}
   );
   gpc1_1 gpc2755 (
      {stage0_6[499]},
      {stage1_6[167]}
   );
   gpc1_1 gpc2756 (
      {stage0_6[500]},
      {stage1_6[168]}
   );
   gpc1_1 gpc2757 (
      {stage0_6[501]},
      {stage1_6[169]}
   );
   gpc1_1 gpc2758 (
      {stage0_6[502]},
      {stage1_6[170]}
   );
   gpc1_1 gpc2759 (
      {stage0_6[503]},
      {stage1_6[171]}
   );
   gpc1_1 gpc2760 (
      {stage0_6[504]},
      {stage1_6[172]}
   );
   gpc1_1 gpc2761 (
      {stage0_6[505]},
      {stage1_6[173]}
   );
   gpc1_1 gpc2762 (
      {stage0_6[506]},
      {stage1_6[174]}
   );
   gpc1_1 gpc2763 (
      {stage0_6[507]},
      {stage1_6[175]}
   );
   gpc1_1 gpc2764 (
      {stage0_6[508]},
      {stage1_6[176]}
   );
   gpc1_1 gpc2765 (
      {stage0_6[509]},
      {stage1_6[177]}
   );
   gpc1_1 gpc2766 (
      {stage0_6[510]},
      {stage1_6[178]}
   );
   gpc1_1 gpc2767 (
      {stage0_6[511]},
      {stage1_6[179]}
   );
   gpc1_1 gpc2768 (
      {stage0_7[364]},
      {stage1_7[192]}
   );
   gpc1_1 gpc2769 (
      {stage0_7[365]},
      {stage1_7[193]}
   );
   gpc1_1 gpc2770 (
      {stage0_7[366]},
      {stage1_7[194]}
   );
   gpc1_1 gpc2771 (
      {stage0_7[367]},
      {stage1_7[195]}
   );
   gpc1_1 gpc2772 (
      {stage0_7[368]},
      {stage1_7[196]}
   );
   gpc1_1 gpc2773 (
      {stage0_7[369]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2774 (
      {stage0_7[370]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2775 (
      {stage0_7[371]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2776 (
      {stage0_7[372]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2777 (
      {stage0_7[373]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2778 (
      {stage0_7[374]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2779 (
      {stage0_7[375]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2780 (
      {stage0_7[376]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2781 (
      {stage0_7[377]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2782 (
      {stage0_7[378]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2783 (
      {stage0_7[379]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2784 (
      {stage0_7[380]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2785 (
      {stage0_7[381]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2786 (
      {stage0_7[382]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2787 (
      {stage0_7[383]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2788 (
      {stage0_7[384]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2789 (
      {stage0_7[385]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2790 (
      {stage0_7[386]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2791 (
      {stage0_7[387]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2792 (
      {stage0_7[388]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2793 (
      {stage0_7[389]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2794 (
      {stage0_7[390]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2795 (
      {stage0_7[391]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2796 (
      {stage0_7[392]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2797 (
      {stage0_7[393]},
      {stage1_7[221]}
   );
   gpc1_1 gpc2798 (
      {stage0_7[394]},
      {stage1_7[222]}
   );
   gpc1_1 gpc2799 (
      {stage0_7[395]},
      {stage1_7[223]}
   );
   gpc1_1 gpc2800 (
      {stage0_7[396]},
      {stage1_7[224]}
   );
   gpc1_1 gpc2801 (
      {stage0_7[397]},
      {stage1_7[225]}
   );
   gpc1_1 gpc2802 (
      {stage0_7[398]},
      {stage1_7[226]}
   );
   gpc1_1 gpc2803 (
      {stage0_7[399]},
      {stage1_7[227]}
   );
   gpc1_1 gpc2804 (
      {stage0_7[400]},
      {stage1_7[228]}
   );
   gpc1_1 gpc2805 (
      {stage0_7[401]},
      {stage1_7[229]}
   );
   gpc1_1 gpc2806 (
      {stage0_7[402]},
      {stage1_7[230]}
   );
   gpc1_1 gpc2807 (
      {stage0_7[403]},
      {stage1_7[231]}
   );
   gpc1_1 gpc2808 (
      {stage0_7[404]},
      {stage1_7[232]}
   );
   gpc1_1 gpc2809 (
      {stage0_7[405]},
      {stage1_7[233]}
   );
   gpc1_1 gpc2810 (
      {stage0_7[406]},
      {stage1_7[234]}
   );
   gpc1_1 gpc2811 (
      {stage0_7[407]},
      {stage1_7[235]}
   );
   gpc1_1 gpc2812 (
      {stage0_7[408]},
      {stage1_7[236]}
   );
   gpc1_1 gpc2813 (
      {stage0_7[409]},
      {stage1_7[237]}
   );
   gpc1_1 gpc2814 (
      {stage0_7[410]},
      {stage1_7[238]}
   );
   gpc1_1 gpc2815 (
      {stage0_7[411]},
      {stage1_7[239]}
   );
   gpc1_1 gpc2816 (
      {stage0_7[412]},
      {stage1_7[240]}
   );
   gpc1_1 gpc2817 (
      {stage0_7[413]},
      {stage1_7[241]}
   );
   gpc1_1 gpc2818 (
      {stage0_7[414]},
      {stage1_7[242]}
   );
   gpc1_1 gpc2819 (
      {stage0_7[415]},
      {stage1_7[243]}
   );
   gpc1_1 gpc2820 (
      {stage0_7[416]},
      {stage1_7[244]}
   );
   gpc1_1 gpc2821 (
      {stage0_7[417]},
      {stage1_7[245]}
   );
   gpc1_1 gpc2822 (
      {stage0_7[418]},
      {stage1_7[246]}
   );
   gpc1_1 gpc2823 (
      {stage0_7[419]},
      {stage1_7[247]}
   );
   gpc1_1 gpc2824 (
      {stage0_7[420]},
      {stage1_7[248]}
   );
   gpc1_1 gpc2825 (
      {stage0_7[421]},
      {stage1_7[249]}
   );
   gpc1_1 gpc2826 (
      {stage0_7[422]},
      {stage1_7[250]}
   );
   gpc1_1 gpc2827 (
      {stage0_7[423]},
      {stage1_7[251]}
   );
   gpc1_1 gpc2828 (
      {stage0_7[424]},
      {stage1_7[252]}
   );
   gpc1_1 gpc2829 (
      {stage0_7[425]},
      {stage1_7[253]}
   );
   gpc1_1 gpc2830 (
      {stage0_7[426]},
      {stage1_7[254]}
   );
   gpc1_1 gpc2831 (
      {stage0_7[427]},
      {stage1_7[255]}
   );
   gpc1_1 gpc2832 (
      {stage0_7[428]},
      {stage1_7[256]}
   );
   gpc1_1 gpc2833 (
      {stage0_7[429]},
      {stage1_7[257]}
   );
   gpc1_1 gpc2834 (
      {stage0_7[430]},
      {stage1_7[258]}
   );
   gpc1_1 gpc2835 (
      {stage0_7[431]},
      {stage1_7[259]}
   );
   gpc1_1 gpc2836 (
      {stage0_7[432]},
      {stage1_7[260]}
   );
   gpc1_1 gpc2837 (
      {stage0_7[433]},
      {stage1_7[261]}
   );
   gpc1_1 gpc2838 (
      {stage0_7[434]},
      {stage1_7[262]}
   );
   gpc1_1 gpc2839 (
      {stage0_7[435]},
      {stage1_7[263]}
   );
   gpc1_1 gpc2840 (
      {stage0_7[436]},
      {stage1_7[264]}
   );
   gpc1_1 gpc2841 (
      {stage0_7[437]},
      {stage1_7[265]}
   );
   gpc1_1 gpc2842 (
      {stage0_7[438]},
      {stage1_7[266]}
   );
   gpc1_1 gpc2843 (
      {stage0_7[439]},
      {stage1_7[267]}
   );
   gpc1_1 gpc2844 (
      {stage0_7[440]},
      {stage1_7[268]}
   );
   gpc1_1 gpc2845 (
      {stage0_7[441]},
      {stage1_7[269]}
   );
   gpc1_1 gpc2846 (
      {stage0_7[442]},
      {stage1_7[270]}
   );
   gpc1_1 gpc2847 (
      {stage0_7[443]},
      {stage1_7[271]}
   );
   gpc1_1 gpc2848 (
      {stage0_7[444]},
      {stage1_7[272]}
   );
   gpc1_1 gpc2849 (
      {stage0_7[445]},
      {stage1_7[273]}
   );
   gpc1_1 gpc2850 (
      {stage0_7[446]},
      {stage1_7[274]}
   );
   gpc1_1 gpc2851 (
      {stage0_7[447]},
      {stage1_7[275]}
   );
   gpc1_1 gpc2852 (
      {stage0_7[448]},
      {stage1_7[276]}
   );
   gpc1_1 gpc2853 (
      {stage0_7[449]},
      {stage1_7[277]}
   );
   gpc1_1 gpc2854 (
      {stage0_7[450]},
      {stage1_7[278]}
   );
   gpc1_1 gpc2855 (
      {stage0_7[451]},
      {stage1_7[279]}
   );
   gpc1_1 gpc2856 (
      {stage0_7[452]},
      {stage1_7[280]}
   );
   gpc1_1 gpc2857 (
      {stage0_7[453]},
      {stage1_7[281]}
   );
   gpc1_1 gpc2858 (
      {stage0_7[454]},
      {stage1_7[282]}
   );
   gpc1_1 gpc2859 (
      {stage0_7[455]},
      {stage1_7[283]}
   );
   gpc1_1 gpc2860 (
      {stage0_7[456]},
      {stage1_7[284]}
   );
   gpc1_1 gpc2861 (
      {stage0_7[457]},
      {stage1_7[285]}
   );
   gpc1_1 gpc2862 (
      {stage0_7[458]},
      {stage1_7[286]}
   );
   gpc1_1 gpc2863 (
      {stage0_7[459]},
      {stage1_7[287]}
   );
   gpc1_1 gpc2864 (
      {stage0_7[460]},
      {stage1_7[288]}
   );
   gpc1_1 gpc2865 (
      {stage0_7[461]},
      {stage1_7[289]}
   );
   gpc1_1 gpc2866 (
      {stage0_7[462]},
      {stage1_7[290]}
   );
   gpc1_1 gpc2867 (
      {stage0_7[463]},
      {stage1_7[291]}
   );
   gpc1_1 gpc2868 (
      {stage0_7[464]},
      {stage1_7[292]}
   );
   gpc1_1 gpc2869 (
      {stage0_7[465]},
      {stage1_7[293]}
   );
   gpc1_1 gpc2870 (
      {stage0_7[466]},
      {stage1_7[294]}
   );
   gpc1_1 gpc2871 (
      {stage0_7[467]},
      {stage1_7[295]}
   );
   gpc1_1 gpc2872 (
      {stage0_7[468]},
      {stage1_7[296]}
   );
   gpc1_1 gpc2873 (
      {stage0_7[469]},
      {stage1_7[297]}
   );
   gpc1_1 gpc2874 (
      {stage0_7[470]},
      {stage1_7[298]}
   );
   gpc1_1 gpc2875 (
      {stage0_7[471]},
      {stage1_7[299]}
   );
   gpc1_1 gpc2876 (
      {stage0_7[472]},
      {stage1_7[300]}
   );
   gpc1_1 gpc2877 (
      {stage0_7[473]},
      {stage1_7[301]}
   );
   gpc1_1 gpc2878 (
      {stage0_7[474]},
      {stage1_7[302]}
   );
   gpc1_1 gpc2879 (
      {stage0_7[475]},
      {stage1_7[303]}
   );
   gpc1_1 gpc2880 (
      {stage0_7[476]},
      {stage1_7[304]}
   );
   gpc1_1 gpc2881 (
      {stage0_7[477]},
      {stage1_7[305]}
   );
   gpc1_1 gpc2882 (
      {stage0_7[478]},
      {stage1_7[306]}
   );
   gpc1_1 gpc2883 (
      {stage0_7[479]},
      {stage1_7[307]}
   );
   gpc1_1 gpc2884 (
      {stage0_7[480]},
      {stage1_7[308]}
   );
   gpc1_1 gpc2885 (
      {stage0_7[481]},
      {stage1_7[309]}
   );
   gpc1_1 gpc2886 (
      {stage0_7[482]},
      {stage1_7[310]}
   );
   gpc1_1 gpc2887 (
      {stage0_7[483]},
      {stage1_7[311]}
   );
   gpc1_1 gpc2888 (
      {stage0_7[484]},
      {stage1_7[312]}
   );
   gpc1_1 gpc2889 (
      {stage0_7[485]},
      {stage1_7[313]}
   );
   gpc1_1 gpc2890 (
      {stage0_7[486]},
      {stage1_7[314]}
   );
   gpc1_1 gpc2891 (
      {stage0_7[487]},
      {stage1_7[315]}
   );
   gpc1_1 gpc2892 (
      {stage0_7[488]},
      {stage1_7[316]}
   );
   gpc1_1 gpc2893 (
      {stage0_7[489]},
      {stage1_7[317]}
   );
   gpc1_1 gpc2894 (
      {stage0_7[490]},
      {stage1_7[318]}
   );
   gpc1_1 gpc2895 (
      {stage0_7[491]},
      {stage1_7[319]}
   );
   gpc1_1 gpc2896 (
      {stage0_7[492]},
      {stage1_7[320]}
   );
   gpc1_1 gpc2897 (
      {stage0_7[493]},
      {stage1_7[321]}
   );
   gpc1_1 gpc2898 (
      {stage0_7[494]},
      {stage1_7[322]}
   );
   gpc1_1 gpc2899 (
      {stage0_7[495]},
      {stage1_7[323]}
   );
   gpc1_1 gpc2900 (
      {stage0_7[496]},
      {stage1_7[324]}
   );
   gpc1_1 gpc2901 (
      {stage0_7[497]},
      {stage1_7[325]}
   );
   gpc1_1 gpc2902 (
      {stage0_7[498]},
      {stage1_7[326]}
   );
   gpc1_1 gpc2903 (
      {stage0_7[499]},
      {stage1_7[327]}
   );
   gpc1_1 gpc2904 (
      {stage0_7[500]},
      {stage1_7[328]}
   );
   gpc1_1 gpc2905 (
      {stage0_7[501]},
      {stage1_7[329]}
   );
   gpc1_1 gpc2906 (
      {stage0_7[502]},
      {stage1_7[330]}
   );
   gpc1_1 gpc2907 (
      {stage0_7[503]},
      {stage1_7[331]}
   );
   gpc1_1 gpc2908 (
      {stage0_7[504]},
      {stage1_7[332]}
   );
   gpc1_1 gpc2909 (
      {stage0_7[505]},
      {stage1_7[333]}
   );
   gpc1_1 gpc2910 (
      {stage0_7[506]},
      {stage1_7[334]}
   );
   gpc1_1 gpc2911 (
      {stage0_7[507]},
      {stage1_7[335]}
   );
   gpc1_1 gpc2912 (
      {stage0_7[508]},
      {stage1_7[336]}
   );
   gpc1_1 gpc2913 (
      {stage0_7[509]},
      {stage1_7[337]}
   );
   gpc1_1 gpc2914 (
      {stage0_7[510]},
      {stage1_7[338]}
   );
   gpc1_1 gpc2915 (
      {stage0_7[511]},
      {stage1_7[339]}
   );
   gpc1_1 gpc2916 (
      {stage0_8[493]},
      {stage1_8[220]}
   );
   gpc1_1 gpc2917 (
      {stage0_8[494]},
      {stage1_8[221]}
   );
   gpc1_1 gpc2918 (
      {stage0_8[495]},
      {stage1_8[222]}
   );
   gpc1_1 gpc2919 (
      {stage0_8[496]},
      {stage1_8[223]}
   );
   gpc1_1 gpc2920 (
      {stage0_8[497]},
      {stage1_8[224]}
   );
   gpc1_1 gpc2921 (
      {stage0_8[498]},
      {stage1_8[225]}
   );
   gpc1_1 gpc2922 (
      {stage0_8[499]},
      {stage1_8[226]}
   );
   gpc1_1 gpc2923 (
      {stage0_8[500]},
      {stage1_8[227]}
   );
   gpc1_1 gpc2924 (
      {stage0_8[501]},
      {stage1_8[228]}
   );
   gpc1_1 gpc2925 (
      {stage0_8[502]},
      {stage1_8[229]}
   );
   gpc1_1 gpc2926 (
      {stage0_8[503]},
      {stage1_8[230]}
   );
   gpc1_1 gpc2927 (
      {stage0_8[504]},
      {stage1_8[231]}
   );
   gpc1_1 gpc2928 (
      {stage0_8[505]},
      {stage1_8[232]}
   );
   gpc1_1 gpc2929 (
      {stage0_8[506]},
      {stage1_8[233]}
   );
   gpc1_1 gpc2930 (
      {stage0_8[507]},
      {stage1_8[234]}
   );
   gpc1_1 gpc2931 (
      {stage0_8[508]},
      {stage1_8[235]}
   );
   gpc1_1 gpc2932 (
      {stage0_8[509]},
      {stage1_8[236]}
   );
   gpc1_1 gpc2933 (
      {stage0_8[510]},
      {stage1_8[237]}
   );
   gpc1_1 gpc2934 (
      {stage0_8[511]},
      {stage1_8[238]}
   );
   gpc1_1 gpc2935 (
      {stage0_9[312]},
      {stage1_9[163]}
   );
   gpc1_1 gpc2936 (
      {stage0_9[313]},
      {stage1_9[164]}
   );
   gpc1_1 gpc2937 (
      {stage0_9[314]},
      {stage1_9[165]}
   );
   gpc1_1 gpc2938 (
      {stage0_9[315]},
      {stage1_9[166]}
   );
   gpc1_1 gpc2939 (
      {stage0_9[316]},
      {stage1_9[167]}
   );
   gpc1_1 gpc2940 (
      {stage0_9[317]},
      {stage1_9[168]}
   );
   gpc1_1 gpc2941 (
      {stage0_9[318]},
      {stage1_9[169]}
   );
   gpc1_1 gpc2942 (
      {stage0_9[319]},
      {stage1_9[170]}
   );
   gpc1_1 gpc2943 (
      {stage0_9[320]},
      {stage1_9[171]}
   );
   gpc1_1 gpc2944 (
      {stage0_9[321]},
      {stage1_9[172]}
   );
   gpc1_1 gpc2945 (
      {stage0_9[322]},
      {stage1_9[173]}
   );
   gpc1_1 gpc2946 (
      {stage0_9[323]},
      {stage1_9[174]}
   );
   gpc1_1 gpc2947 (
      {stage0_9[324]},
      {stage1_9[175]}
   );
   gpc1_1 gpc2948 (
      {stage0_9[325]},
      {stage1_9[176]}
   );
   gpc1_1 gpc2949 (
      {stage0_9[326]},
      {stage1_9[177]}
   );
   gpc1_1 gpc2950 (
      {stage0_9[327]},
      {stage1_9[178]}
   );
   gpc1_1 gpc2951 (
      {stage0_9[328]},
      {stage1_9[179]}
   );
   gpc1_1 gpc2952 (
      {stage0_9[329]},
      {stage1_9[180]}
   );
   gpc1_1 gpc2953 (
      {stage0_9[330]},
      {stage1_9[181]}
   );
   gpc1_1 gpc2954 (
      {stage0_9[331]},
      {stage1_9[182]}
   );
   gpc1_1 gpc2955 (
      {stage0_9[332]},
      {stage1_9[183]}
   );
   gpc1_1 gpc2956 (
      {stage0_9[333]},
      {stage1_9[184]}
   );
   gpc1_1 gpc2957 (
      {stage0_9[334]},
      {stage1_9[185]}
   );
   gpc1_1 gpc2958 (
      {stage0_9[335]},
      {stage1_9[186]}
   );
   gpc1_1 gpc2959 (
      {stage0_9[336]},
      {stage1_9[187]}
   );
   gpc1_1 gpc2960 (
      {stage0_9[337]},
      {stage1_9[188]}
   );
   gpc1_1 gpc2961 (
      {stage0_9[338]},
      {stage1_9[189]}
   );
   gpc1_1 gpc2962 (
      {stage0_9[339]},
      {stage1_9[190]}
   );
   gpc1_1 gpc2963 (
      {stage0_9[340]},
      {stage1_9[191]}
   );
   gpc1_1 gpc2964 (
      {stage0_9[341]},
      {stage1_9[192]}
   );
   gpc1_1 gpc2965 (
      {stage0_9[342]},
      {stage1_9[193]}
   );
   gpc1_1 gpc2966 (
      {stage0_9[343]},
      {stage1_9[194]}
   );
   gpc1_1 gpc2967 (
      {stage0_9[344]},
      {stage1_9[195]}
   );
   gpc1_1 gpc2968 (
      {stage0_9[345]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2969 (
      {stage0_9[346]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2970 (
      {stage0_9[347]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2971 (
      {stage0_9[348]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2972 (
      {stage0_9[349]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2973 (
      {stage0_9[350]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2974 (
      {stage0_9[351]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2975 (
      {stage0_9[352]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2976 (
      {stage0_9[353]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2977 (
      {stage0_9[354]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2978 (
      {stage0_9[355]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2979 (
      {stage0_9[356]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2980 (
      {stage0_9[357]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2981 (
      {stage0_9[358]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2982 (
      {stage0_9[359]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2983 (
      {stage0_9[360]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2984 (
      {stage0_9[361]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2985 (
      {stage0_9[362]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2986 (
      {stage0_9[363]},
      {stage1_9[214]}
   );
   gpc1_1 gpc2987 (
      {stage0_9[364]},
      {stage1_9[215]}
   );
   gpc1_1 gpc2988 (
      {stage0_9[365]},
      {stage1_9[216]}
   );
   gpc1_1 gpc2989 (
      {stage0_9[366]},
      {stage1_9[217]}
   );
   gpc1_1 gpc2990 (
      {stage0_9[367]},
      {stage1_9[218]}
   );
   gpc1_1 gpc2991 (
      {stage0_9[368]},
      {stage1_9[219]}
   );
   gpc1_1 gpc2992 (
      {stage0_9[369]},
      {stage1_9[220]}
   );
   gpc1_1 gpc2993 (
      {stage0_9[370]},
      {stage1_9[221]}
   );
   gpc1_1 gpc2994 (
      {stage0_9[371]},
      {stage1_9[222]}
   );
   gpc1_1 gpc2995 (
      {stage0_9[372]},
      {stage1_9[223]}
   );
   gpc1_1 gpc2996 (
      {stage0_9[373]},
      {stage1_9[224]}
   );
   gpc1_1 gpc2997 (
      {stage0_9[374]},
      {stage1_9[225]}
   );
   gpc1_1 gpc2998 (
      {stage0_9[375]},
      {stage1_9[226]}
   );
   gpc1_1 gpc2999 (
      {stage0_9[376]},
      {stage1_9[227]}
   );
   gpc1_1 gpc3000 (
      {stage0_9[377]},
      {stage1_9[228]}
   );
   gpc1_1 gpc3001 (
      {stage0_9[378]},
      {stage1_9[229]}
   );
   gpc1_1 gpc3002 (
      {stage0_9[379]},
      {stage1_9[230]}
   );
   gpc1_1 gpc3003 (
      {stage0_9[380]},
      {stage1_9[231]}
   );
   gpc1_1 gpc3004 (
      {stage0_9[381]},
      {stage1_9[232]}
   );
   gpc1_1 gpc3005 (
      {stage0_9[382]},
      {stage1_9[233]}
   );
   gpc1_1 gpc3006 (
      {stage0_9[383]},
      {stage1_9[234]}
   );
   gpc1_1 gpc3007 (
      {stage0_9[384]},
      {stage1_9[235]}
   );
   gpc1_1 gpc3008 (
      {stage0_9[385]},
      {stage1_9[236]}
   );
   gpc1_1 gpc3009 (
      {stage0_9[386]},
      {stage1_9[237]}
   );
   gpc1_1 gpc3010 (
      {stage0_9[387]},
      {stage1_9[238]}
   );
   gpc1_1 gpc3011 (
      {stage0_9[388]},
      {stage1_9[239]}
   );
   gpc1_1 gpc3012 (
      {stage0_9[389]},
      {stage1_9[240]}
   );
   gpc1_1 gpc3013 (
      {stage0_9[390]},
      {stage1_9[241]}
   );
   gpc1_1 gpc3014 (
      {stage0_9[391]},
      {stage1_9[242]}
   );
   gpc1_1 gpc3015 (
      {stage0_9[392]},
      {stage1_9[243]}
   );
   gpc1_1 gpc3016 (
      {stage0_9[393]},
      {stage1_9[244]}
   );
   gpc1_1 gpc3017 (
      {stage0_9[394]},
      {stage1_9[245]}
   );
   gpc1_1 gpc3018 (
      {stage0_9[395]},
      {stage1_9[246]}
   );
   gpc1_1 gpc3019 (
      {stage0_9[396]},
      {stage1_9[247]}
   );
   gpc1_1 gpc3020 (
      {stage0_9[397]},
      {stage1_9[248]}
   );
   gpc1_1 gpc3021 (
      {stage0_9[398]},
      {stage1_9[249]}
   );
   gpc1_1 gpc3022 (
      {stage0_9[399]},
      {stage1_9[250]}
   );
   gpc1_1 gpc3023 (
      {stage0_9[400]},
      {stage1_9[251]}
   );
   gpc1_1 gpc3024 (
      {stage0_9[401]},
      {stage1_9[252]}
   );
   gpc1_1 gpc3025 (
      {stage0_9[402]},
      {stage1_9[253]}
   );
   gpc1_1 gpc3026 (
      {stage0_9[403]},
      {stage1_9[254]}
   );
   gpc1_1 gpc3027 (
      {stage0_9[404]},
      {stage1_9[255]}
   );
   gpc1_1 gpc3028 (
      {stage0_9[405]},
      {stage1_9[256]}
   );
   gpc1_1 gpc3029 (
      {stage0_9[406]},
      {stage1_9[257]}
   );
   gpc1_1 gpc3030 (
      {stage0_9[407]},
      {stage1_9[258]}
   );
   gpc1_1 gpc3031 (
      {stage0_9[408]},
      {stage1_9[259]}
   );
   gpc1_1 gpc3032 (
      {stage0_9[409]},
      {stage1_9[260]}
   );
   gpc1_1 gpc3033 (
      {stage0_9[410]},
      {stage1_9[261]}
   );
   gpc1_1 gpc3034 (
      {stage0_9[411]},
      {stage1_9[262]}
   );
   gpc1_1 gpc3035 (
      {stage0_9[412]},
      {stage1_9[263]}
   );
   gpc1_1 gpc3036 (
      {stage0_9[413]},
      {stage1_9[264]}
   );
   gpc1_1 gpc3037 (
      {stage0_9[414]},
      {stage1_9[265]}
   );
   gpc1_1 gpc3038 (
      {stage0_9[415]},
      {stage1_9[266]}
   );
   gpc1_1 gpc3039 (
      {stage0_9[416]},
      {stage1_9[267]}
   );
   gpc1_1 gpc3040 (
      {stage0_9[417]},
      {stage1_9[268]}
   );
   gpc1_1 gpc3041 (
      {stage0_9[418]},
      {stage1_9[269]}
   );
   gpc1_1 gpc3042 (
      {stage0_9[419]},
      {stage1_9[270]}
   );
   gpc1_1 gpc3043 (
      {stage0_9[420]},
      {stage1_9[271]}
   );
   gpc1_1 gpc3044 (
      {stage0_9[421]},
      {stage1_9[272]}
   );
   gpc1_1 gpc3045 (
      {stage0_9[422]},
      {stage1_9[273]}
   );
   gpc1_1 gpc3046 (
      {stage0_9[423]},
      {stage1_9[274]}
   );
   gpc1_1 gpc3047 (
      {stage0_9[424]},
      {stage1_9[275]}
   );
   gpc1_1 gpc3048 (
      {stage0_9[425]},
      {stage1_9[276]}
   );
   gpc1_1 gpc3049 (
      {stage0_9[426]},
      {stage1_9[277]}
   );
   gpc1_1 gpc3050 (
      {stage0_9[427]},
      {stage1_9[278]}
   );
   gpc1_1 gpc3051 (
      {stage0_9[428]},
      {stage1_9[279]}
   );
   gpc1_1 gpc3052 (
      {stage0_9[429]},
      {stage1_9[280]}
   );
   gpc1_1 gpc3053 (
      {stage0_9[430]},
      {stage1_9[281]}
   );
   gpc1_1 gpc3054 (
      {stage0_9[431]},
      {stage1_9[282]}
   );
   gpc1_1 gpc3055 (
      {stage0_9[432]},
      {stage1_9[283]}
   );
   gpc1_1 gpc3056 (
      {stage0_9[433]},
      {stage1_9[284]}
   );
   gpc1_1 gpc3057 (
      {stage0_9[434]},
      {stage1_9[285]}
   );
   gpc1_1 gpc3058 (
      {stage0_9[435]},
      {stage1_9[286]}
   );
   gpc1_1 gpc3059 (
      {stage0_9[436]},
      {stage1_9[287]}
   );
   gpc1_1 gpc3060 (
      {stage0_9[437]},
      {stage1_9[288]}
   );
   gpc1_1 gpc3061 (
      {stage0_9[438]},
      {stage1_9[289]}
   );
   gpc1_1 gpc3062 (
      {stage0_9[439]},
      {stage1_9[290]}
   );
   gpc1_1 gpc3063 (
      {stage0_9[440]},
      {stage1_9[291]}
   );
   gpc1_1 gpc3064 (
      {stage0_9[441]},
      {stage1_9[292]}
   );
   gpc1_1 gpc3065 (
      {stage0_9[442]},
      {stage1_9[293]}
   );
   gpc1_1 gpc3066 (
      {stage0_9[443]},
      {stage1_9[294]}
   );
   gpc1_1 gpc3067 (
      {stage0_9[444]},
      {stage1_9[295]}
   );
   gpc1_1 gpc3068 (
      {stage0_9[445]},
      {stage1_9[296]}
   );
   gpc1_1 gpc3069 (
      {stage0_9[446]},
      {stage1_9[297]}
   );
   gpc1_1 gpc3070 (
      {stage0_9[447]},
      {stage1_9[298]}
   );
   gpc1_1 gpc3071 (
      {stage0_9[448]},
      {stage1_9[299]}
   );
   gpc1_1 gpc3072 (
      {stage0_9[449]},
      {stage1_9[300]}
   );
   gpc1_1 gpc3073 (
      {stage0_9[450]},
      {stage1_9[301]}
   );
   gpc1_1 gpc3074 (
      {stage0_9[451]},
      {stage1_9[302]}
   );
   gpc1_1 gpc3075 (
      {stage0_9[452]},
      {stage1_9[303]}
   );
   gpc1_1 gpc3076 (
      {stage0_9[453]},
      {stage1_9[304]}
   );
   gpc1_1 gpc3077 (
      {stage0_9[454]},
      {stage1_9[305]}
   );
   gpc1_1 gpc3078 (
      {stage0_9[455]},
      {stage1_9[306]}
   );
   gpc1_1 gpc3079 (
      {stage0_9[456]},
      {stage1_9[307]}
   );
   gpc1_1 gpc3080 (
      {stage0_9[457]},
      {stage1_9[308]}
   );
   gpc1_1 gpc3081 (
      {stage0_9[458]},
      {stage1_9[309]}
   );
   gpc1_1 gpc3082 (
      {stage0_9[459]},
      {stage1_9[310]}
   );
   gpc1_1 gpc3083 (
      {stage0_9[460]},
      {stage1_9[311]}
   );
   gpc1_1 gpc3084 (
      {stage0_9[461]},
      {stage1_9[312]}
   );
   gpc1_1 gpc3085 (
      {stage0_9[462]},
      {stage1_9[313]}
   );
   gpc1_1 gpc3086 (
      {stage0_9[463]},
      {stage1_9[314]}
   );
   gpc1_1 gpc3087 (
      {stage0_9[464]},
      {stage1_9[315]}
   );
   gpc1_1 gpc3088 (
      {stage0_9[465]},
      {stage1_9[316]}
   );
   gpc1_1 gpc3089 (
      {stage0_9[466]},
      {stage1_9[317]}
   );
   gpc1_1 gpc3090 (
      {stage0_9[467]},
      {stage1_9[318]}
   );
   gpc1_1 gpc3091 (
      {stage0_9[468]},
      {stage1_9[319]}
   );
   gpc1_1 gpc3092 (
      {stage0_9[469]},
      {stage1_9[320]}
   );
   gpc1_1 gpc3093 (
      {stage0_9[470]},
      {stage1_9[321]}
   );
   gpc1_1 gpc3094 (
      {stage0_9[471]},
      {stage1_9[322]}
   );
   gpc1_1 gpc3095 (
      {stage0_9[472]},
      {stage1_9[323]}
   );
   gpc1_1 gpc3096 (
      {stage0_9[473]},
      {stage1_9[324]}
   );
   gpc1_1 gpc3097 (
      {stage0_9[474]},
      {stage1_9[325]}
   );
   gpc1_1 gpc3098 (
      {stage0_9[475]},
      {stage1_9[326]}
   );
   gpc1_1 gpc3099 (
      {stage0_9[476]},
      {stage1_9[327]}
   );
   gpc1_1 gpc3100 (
      {stage0_9[477]},
      {stage1_9[328]}
   );
   gpc1_1 gpc3101 (
      {stage0_9[478]},
      {stage1_9[329]}
   );
   gpc1_1 gpc3102 (
      {stage0_9[479]},
      {stage1_9[330]}
   );
   gpc1_1 gpc3103 (
      {stage0_9[480]},
      {stage1_9[331]}
   );
   gpc1_1 gpc3104 (
      {stage0_9[481]},
      {stage1_9[332]}
   );
   gpc1_1 gpc3105 (
      {stage0_9[482]},
      {stage1_9[333]}
   );
   gpc1_1 gpc3106 (
      {stage0_9[483]},
      {stage1_9[334]}
   );
   gpc1_1 gpc3107 (
      {stage0_9[484]},
      {stage1_9[335]}
   );
   gpc1_1 gpc3108 (
      {stage0_9[485]},
      {stage1_9[336]}
   );
   gpc1_1 gpc3109 (
      {stage0_9[486]},
      {stage1_9[337]}
   );
   gpc1_1 gpc3110 (
      {stage0_9[487]},
      {stage1_9[338]}
   );
   gpc1_1 gpc3111 (
      {stage0_9[488]},
      {stage1_9[339]}
   );
   gpc1_1 gpc3112 (
      {stage0_9[489]},
      {stage1_9[340]}
   );
   gpc1_1 gpc3113 (
      {stage0_9[490]},
      {stage1_9[341]}
   );
   gpc1_1 gpc3114 (
      {stage0_9[491]},
      {stage1_9[342]}
   );
   gpc1_1 gpc3115 (
      {stage0_9[492]},
      {stage1_9[343]}
   );
   gpc1_1 gpc3116 (
      {stage0_9[493]},
      {stage1_9[344]}
   );
   gpc1_1 gpc3117 (
      {stage0_9[494]},
      {stage1_9[345]}
   );
   gpc1_1 gpc3118 (
      {stage0_9[495]},
      {stage1_9[346]}
   );
   gpc1_1 gpc3119 (
      {stage0_9[496]},
      {stage1_9[347]}
   );
   gpc1_1 gpc3120 (
      {stage0_9[497]},
      {stage1_9[348]}
   );
   gpc1_1 gpc3121 (
      {stage0_9[498]},
      {stage1_9[349]}
   );
   gpc1_1 gpc3122 (
      {stage0_9[499]},
      {stage1_9[350]}
   );
   gpc1_1 gpc3123 (
      {stage0_9[500]},
      {stage1_9[351]}
   );
   gpc1_1 gpc3124 (
      {stage0_9[501]},
      {stage1_9[352]}
   );
   gpc1_1 gpc3125 (
      {stage0_9[502]},
      {stage1_9[353]}
   );
   gpc1_1 gpc3126 (
      {stage0_9[503]},
      {stage1_9[354]}
   );
   gpc1_1 gpc3127 (
      {stage0_9[504]},
      {stage1_9[355]}
   );
   gpc1_1 gpc3128 (
      {stage0_9[505]},
      {stage1_9[356]}
   );
   gpc1_1 gpc3129 (
      {stage0_9[506]},
      {stage1_9[357]}
   );
   gpc1_1 gpc3130 (
      {stage0_9[507]},
      {stage1_9[358]}
   );
   gpc1_1 gpc3131 (
      {stage0_9[508]},
      {stage1_9[359]}
   );
   gpc1_1 gpc3132 (
      {stage0_9[509]},
      {stage1_9[360]}
   );
   gpc1_1 gpc3133 (
      {stage0_9[510]},
      {stage1_9[361]}
   );
   gpc1_1 gpc3134 (
      {stage0_9[511]},
      {stage1_9[362]}
   );
   gpc1_1 gpc3135 (
      {stage0_10[502]},
      {stage1_10[143]}
   );
   gpc1_1 gpc3136 (
      {stage0_10[503]},
      {stage1_10[144]}
   );
   gpc1_1 gpc3137 (
      {stage0_10[504]},
      {stage1_10[145]}
   );
   gpc1_1 gpc3138 (
      {stage0_10[505]},
      {stage1_10[146]}
   );
   gpc1_1 gpc3139 (
      {stage0_10[506]},
      {stage1_10[147]}
   );
   gpc1_1 gpc3140 (
      {stage0_10[507]},
      {stage1_10[148]}
   );
   gpc1_1 gpc3141 (
      {stage0_10[508]},
      {stage1_10[149]}
   );
   gpc1_1 gpc3142 (
      {stage0_10[509]},
      {stage1_10[150]}
   );
   gpc1_1 gpc3143 (
      {stage0_10[510]},
      {stage1_10[151]}
   );
   gpc1_1 gpc3144 (
      {stage0_10[511]},
      {stage1_10[152]}
   );
   gpc1_1 gpc3145 (
      {stage0_11[380]},
      {stage1_11[186]}
   );
   gpc1_1 gpc3146 (
      {stage0_11[381]},
      {stage1_11[187]}
   );
   gpc1_1 gpc3147 (
      {stage0_11[382]},
      {stage1_11[188]}
   );
   gpc1_1 gpc3148 (
      {stage0_11[383]},
      {stage1_11[189]}
   );
   gpc1_1 gpc3149 (
      {stage0_11[384]},
      {stage1_11[190]}
   );
   gpc1_1 gpc3150 (
      {stage0_11[385]},
      {stage1_11[191]}
   );
   gpc1_1 gpc3151 (
      {stage0_11[386]},
      {stage1_11[192]}
   );
   gpc1_1 gpc3152 (
      {stage0_11[387]},
      {stage1_11[193]}
   );
   gpc1_1 gpc3153 (
      {stage0_11[388]},
      {stage1_11[194]}
   );
   gpc1_1 gpc3154 (
      {stage0_11[389]},
      {stage1_11[195]}
   );
   gpc1_1 gpc3155 (
      {stage0_11[390]},
      {stage1_11[196]}
   );
   gpc1_1 gpc3156 (
      {stage0_11[391]},
      {stage1_11[197]}
   );
   gpc1_1 gpc3157 (
      {stage0_11[392]},
      {stage1_11[198]}
   );
   gpc1_1 gpc3158 (
      {stage0_11[393]},
      {stage1_11[199]}
   );
   gpc1_1 gpc3159 (
      {stage0_11[394]},
      {stage1_11[200]}
   );
   gpc1_1 gpc3160 (
      {stage0_11[395]},
      {stage1_11[201]}
   );
   gpc1_1 gpc3161 (
      {stage0_11[396]},
      {stage1_11[202]}
   );
   gpc1_1 gpc3162 (
      {stage0_11[397]},
      {stage1_11[203]}
   );
   gpc1_1 gpc3163 (
      {stage0_11[398]},
      {stage1_11[204]}
   );
   gpc1_1 gpc3164 (
      {stage0_11[399]},
      {stage1_11[205]}
   );
   gpc1_1 gpc3165 (
      {stage0_11[400]},
      {stage1_11[206]}
   );
   gpc1_1 gpc3166 (
      {stage0_11[401]},
      {stage1_11[207]}
   );
   gpc1_1 gpc3167 (
      {stage0_11[402]},
      {stage1_11[208]}
   );
   gpc1_1 gpc3168 (
      {stage0_11[403]},
      {stage1_11[209]}
   );
   gpc1_1 gpc3169 (
      {stage0_11[404]},
      {stage1_11[210]}
   );
   gpc1_1 gpc3170 (
      {stage0_11[405]},
      {stage1_11[211]}
   );
   gpc1_1 gpc3171 (
      {stage0_11[406]},
      {stage1_11[212]}
   );
   gpc1_1 gpc3172 (
      {stage0_11[407]},
      {stage1_11[213]}
   );
   gpc1_1 gpc3173 (
      {stage0_11[408]},
      {stage1_11[214]}
   );
   gpc1_1 gpc3174 (
      {stage0_11[409]},
      {stage1_11[215]}
   );
   gpc1_1 gpc3175 (
      {stage0_11[410]},
      {stage1_11[216]}
   );
   gpc1_1 gpc3176 (
      {stage0_11[411]},
      {stage1_11[217]}
   );
   gpc1_1 gpc3177 (
      {stage0_11[412]},
      {stage1_11[218]}
   );
   gpc1_1 gpc3178 (
      {stage0_11[413]},
      {stage1_11[219]}
   );
   gpc1_1 gpc3179 (
      {stage0_11[414]},
      {stage1_11[220]}
   );
   gpc1_1 gpc3180 (
      {stage0_11[415]},
      {stage1_11[221]}
   );
   gpc1_1 gpc3181 (
      {stage0_11[416]},
      {stage1_11[222]}
   );
   gpc1_1 gpc3182 (
      {stage0_11[417]},
      {stage1_11[223]}
   );
   gpc1_1 gpc3183 (
      {stage0_11[418]},
      {stage1_11[224]}
   );
   gpc1_1 gpc3184 (
      {stage0_11[419]},
      {stage1_11[225]}
   );
   gpc1_1 gpc3185 (
      {stage0_11[420]},
      {stage1_11[226]}
   );
   gpc1_1 gpc3186 (
      {stage0_11[421]},
      {stage1_11[227]}
   );
   gpc1_1 gpc3187 (
      {stage0_11[422]},
      {stage1_11[228]}
   );
   gpc1_1 gpc3188 (
      {stage0_11[423]},
      {stage1_11[229]}
   );
   gpc1_1 gpc3189 (
      {stage0_11[424]},
      {stage1_11[230]}
   );
   gpc1_1 gpc3190 (
      {stage0_11[425]},
      {stage1_11[231]}
   );
   gpc1_1 gpc3191 (
      {stage0_11[426]},
      {stage1_11[232]}
   );
   gpc1_1 gpc3192 (
      {stage0_11[427]},
      {stage1_11[233]}
   );
   gpc1_1 gpc3193 (
      {stage0_11[428]},
      {stage1_11[234]}
   );
   gpc1_1 gpc3194 (
      {stage0_11[429]},
      {stage1_11[235]}
   );
   gpc1_1 gpc3195 (
      {stage0_11[430]},
      {stage1_11[236]}
   );
   gpc1_1 gpc3196 (
      {stage0_11[431]},
      {stage1_11[237]}
   );
   gpc1_1 gpc3197 (
      {stage0_11[432]},
      {stage1_11[238]}
   );
   gpc1_1 gpc3198 (
      {stage0_11[433]},
      {stage1_11[239]}
   );
   gpc1_1 gpc3199 (
      {stage0_11[434]},
      {stage1_11[240]}
   );
   gpc1_1 gpc3200 (
      {stage0_11[435]},
      {stage1_11[241]}
   );
   gpc1_1 gpc3201 (
      {stage0_11[436]},
      {stage1_11[242]}
   );
   gpc1_1 gpc3202 (
      {stage0_11[437]},
      {stage1_11[243]}
   );
   gpc1_1 gpc3203 (
      {stage0_11[438]},
      {stage1_11[244]}
   );
   gpc1_1 gpc3204 (
      {stage0_11[439]},
      {stage1_11[245]}
   );
   gpc1_1 gpc3205 (
      {stage0_11[440]},
      {stage1_11[246]}
   );
   gpc1_1 gpc3206 (
      {stage0_11[441]},
      {stage1_11[247]}
   );
   gpc1_1 gpc3207 (
      {stage0_11[442]},
      {stage1_11[248]}
   );
   gpc1_1 gpc3208 (
      {stage0_11[443]},
      {stage1_11[249]}
   );
   gpc1_1 gpc3209 (
      {stage0_11[444]},
      {stage1_11[250]}
   );
   gpc1_1 gpc3210 (
      {stage0_11[445]},
      {stage1_11[251]}
   );
   gpc1_1 gpc3211 (
      {stage0_11[446]},
      {stage1_11[252]}
   );
   gpc1_1 gpc3212 (
      {stage0_11[447]},
      {stage1_11[253]}
   );
   gpc1_1 gpc3213 (
      {stage0_11[448]},
      {stage1_11[254]}
   );
   gpc1_1 gpc3214 (
      {stage0_11[449]},
      {stage1_11[255]}
   );
   gpc1_1 gpc3215 (
      {stage0_11[450]},
      {stage1_11[256]}
   );
   gpc1_1 gpc3216 (
      {stage0_11[451]},
      {stage1_11[257]}
   );
   gpc1_1 gpc3217 (
      {stage0_11[452]},
      {stage1_11[258]}
   );
   gpc1_1 gpc3218 (
      {stage0_11[453]},
      {stage1_11[259]}
   );
   gpc1_1 gpc3219 (
      {stage0_11[454]},
      {stage1_11[260]}
   );
   gpc1_1 gpc3220 (
      {stage0_11[455]},
      {stage1_11[261]}
   );
   gpc1_1 gpc3221 (
      {stage0_11[456]},
      {stage1_11[262]}
   );
   gpc1_1 gpc3222 (
      {stage0_11[457]},
      {stage1_11[263]}
   );
   gpc1_1 gpc3223 (
      {stage0_11[458]},
      {stage1_11[264]}
   );
   gpc1_1 gpc3224 (
      {stage0_11[459]},
      {stage1_11[265]}
   );
   gpc1_1 gpc3225 (
      {stage0_11[460]},
      {stage1_11[266]}
   );
   gpc1_1 gpc3226 (
      {stage0_11[461]},
      {stage1_11[267]}
   );
   gpc1_1 gpc3227 (
      {stage0_11[462]},
      {stage1_11[268]}
   );
   gpc1_1 gpc3228 (
      {stage0_11[463]},
      {stage1_11[269]}
   );
   gpc1_1 gpc3229 (
      {stage0_11[464]},
      {stage1_11[270]}
   );
   gpc1_1 gpc3230 (
      {stage0_11[465]},
      {stage1_11[271]}
   );
   gpc1_1 gpc3231 (
      {stage0_11[466]},
      {stage1_11[272]}
   );
   gpc1_1 gpc3232 (
      {stage0_11[467]},
      {stage1_11[273]}
   );
   gpc1_1 gpc3233 (
      {stage0_11[468]},
      {stage1_11[274]}
   );
   gpc1_1 gpc3234 (
      {stage0_11[469]},
      {stage1_11[275]}
   );
   gpc1_1 gpc3235 (
      {stage0_11[470]},
      {stage1_11[276]}
   );
   gpc1_1 gpc3236 (
      {stage0_11[471]},
      {stage1_11[277]}
   );
   gpc1_1 gpc3237 (
      {stage0_11[472]},
      {stage1_11[278]}
   );
   gpc1_1 gpc3238 (
      {stage0_11[473]},
      {stage1_11[279]}
   );
   gpc1_1 gpc3239 (
      {stage0_11[474]},
      {stage1_11[280]}
   );
   gpc1_1 gpc3240 (
      {stage0_11[475]},
      {stage1_11[281]}
   );
   gpc1_1 gpc3241 (
      {stage0_11[476]},
      {stage1_11[282]}
   );
   gpc1_1 gpc3242 (
      {stage0_11[477]},
      {stage1_11[283]}
   );
   gpc1_1 gpc3243 (
      {stage0_11[478]},
      {stage1_11[284]}
   );
   gpc1_1 gpc3244 (
      {stage0_11[479]},
      {stage1_11[285]}
   );
   gpc1_1 gpc3245 (
      {stage0_11[480]},
      {stage1_11[286]}
   );
   gpc1_1 gpc3246 (
      {stage0_11[481]},
      {stage1_11[287]}
   );
   gpc1_1 gpc3247 (
      {stage0_11[482]},
      {stage1_11[288]}
   );
   gpc1_1 gpc3248 (
      {stage0_11[483]},
      {stage1_11[289]}
   );
   gpc1_1 gpc3249 (
      {stage0_11[484]},
      {stage1_11[290]}
   );
   gpc1_1 gpc3250 (
      {stage0_11[485]},
      {stage1_11[291]}
   );
   gpc1_1 gpc3251 (
      {stage0_11[486]},
      {stage1_11[292]}
   );
   gpc1_1 gpc3252 (
      {stage0_11[487]},
      {stage1_11[293]}
   );
   gpc1_1 gpc3253 (
      {stage0_11[488]},
      {stage1_11[294]}
   );
   gpc1_1 gpc3254 (
      {stage0_11[489]},
      {stage1_11[295]}
   );
   gpc1_1 gpc3255 (
      {stage0_11[490]},
      {stage1_11[296]}
   );
   gpc1_1 gpc3256 (
      {stage0_11[491]},
      {stage1_11[297]}
   );
   gpc1_1 gpc3257 (
      {stage0_11[492]},
      {stage1_11[298]}
   );
   gpc1_1 gpc3258 (
      {stage0_11[493]},
      {stage1_11[299]}
   );
   gpc1_1 gpc3259 (
      {stage0_11[494]},
      {stage1_11[300]}
   );
   gpc1_1 gpc3260 (
      {stage0_11[495]},
      {stage1_11[301]}
   );
   gpc1_1 gpc3261 (
      {stage0_11[496]},
      {stage1_11[302]}
   );
   gpc1_1 gpc3262 (
      {stage0_11[497]},
      {stage1_11[303]}
   );
   gpc1_1 gpc3263 (
      {stage0_11[498]},
      {stage1_11[304]}
   );
   gpc1_1 gpc3264 (
      {stage0_11[499]},
      {stage1_11[305]}
   );
   gpc1_1 gpc3265 (
      {stage0_11[500]},
      {stage1_11[306]}
   );
   gpc1_1 gpc3266 (
      {stage0_11[501]},
      {stage1_11[307]}
   );
   gpc1_1 gpc3267 (
      {stage0_11[502]},
      {stage1_11[308]}
   );
   gpc1_1 gpc3268 (
      {stage0_11[503]},
      {stage1_11[309]}
   );
   gpc1_1 gpc3269 (
      {stage0_11[504]},
      {stage1_11[310]}
   );
   gpc1_1 gpc3270 (
      {stage0_11[505]},
      {stage1_11[311]}
   );
   gpc1_1 gpc3271 (
      {stage0_11[506]},
      {stage1_11[312]}
   );
   gpc1_1 gpc3272 (
      {stage0_11[507]},
      {stage1_11[313]}
   );
   gpc1_1 gpc3273 (
      {stage0_11[508]},
      {stage1_11[314]}
   );
   gpc1_1 gpc3274 (
      {stage0_11[509]},
      {stage1_11[315]}
   );
   gpc1_1 gpc3275 (
      {stage0_11[510]},
      {stage1_11[316]}
   );
   gpc1_1 gpc3276 (
      {stage0_11[511]},
      {stage1_11[317]}
   );
   gpc1_1 gpc3277 (
      {stage0_14[429]},
      {stage1_14[173]}
   );
   gpc1_1 gpc3278 (
      {stage0_14[430]},
      {stage1_14[174]}
   );
   gpc1_1 gpc3279 (
      {stage0_14[431]},
      {stage1_14[175]}
   );
   gpc1_1 gpc3280 (
      {stage0_14[432]},
      {stage1_14[176]}
   );
   gpc1_1 gpc3281 (
      {stage0_14[433]},
      {stage1_14[177]}
   );
   gpc1_1 gpc3282 (
      {stage0_14[434]},
      {stage1_14[178]}
   );
   gpc1_1 gpc3283 (
      {stage0_14[435]},
      {stage1_14[179]}
   );
   gpc1_1 gpc3284 (
      {stage0_14[436]},
      {stage1_14[180]}
   );
   gpc1_1 gpc3285 (
      {stage0_14[437]},
      {stage1_14[181]}
   );
   gpc1_1 gpc3286 (
      {stage0_14[438]},
      {stage1_14[182]}
   );
   gpc1_1 gpc3287 (
      {stage0_14[439]},
      {stage1_14[183]}
   );
   gpc1_1 gpc3288 (
      {stage0_14[440]},
      {stage1_14[184]}
   );
   gpc1_1 gpc3289 (
      {stage0_14[441]},
      {stage1_14[185]}
   );
   gpc1_1 gpc3290 (
      {stage0_14[442]},
      {stage1_14[186]}
   );
   gpc1_1 gpc3291 (
      {stage0_14[443]},
      {stage1_14[187]}
   );
   gpc1_1 gpc3292 (
      {stage0_14[444]},
      {stage1_14[188]}
   );
   gpc1_1 gpc3293 (
      {stage0_14[445]},
      {stage1_14[189]}
   );
   gpc1_1 gpc3294 (
      {stage0_14[446]},
      {stage1_14[190]}
   );
   gpc1_1 gpc3295 (
      {stage0_14[447]},
      {stage1_14[191]}
   );
   gpc1_1 gpc3296 (
      {stage0_14[448]},
      {stage1_14[192]}
   );
   gpc1_1 gpc3297 (
      {stage0_14[449]},
      {stage1_14[193]}
   );
   gpc1_1 gpc3298 (
      {stage0_14[450]},
      {stage1_14[194]}
   );
   gpc1_1 gpc3299 (
      {stage0_14[451]},
      {stage1_14[195]}
   );
   gpc1_1 gpc3300 (
      {stage0_14[452]},
      {stage1_14[196]}
   );
   gpc1_1 gpc3301 (
      {stage0_14[453]},
      {stage1_14[197]}
   );
   gpc1_1 gpc3302 (
      {stage0_14[454]},
      {stage1_14[198]}
   );
   gpc1_1 gpc3303 (
      {stage0_14[455]},
      {stage1_14[199]}
   );
   gpc1_1 gpc3304 (
      {stage0_14[456]},
      {stage1_14[200]}
   );
   gpc1_1 gpc3305 (
      {stage0_14[457]},
      {stage1_14[201]}
   );
   gpc1_1 gpc3306 (
      {stage0_14[458]},
      {stage1_14[202]}
   );
   gpc1_1 gpc3307 (
      {stage0_14[459]},
      {stage1_14[203]}
   );
   gpc1_1 gpc3308 (
      {stage0_14[460]},
      {stage1_14[204]}
   );
   gpc1_1 gpc3309 (
      {stage0_14[461]},
      {stage1_14[205]}
   );
   gpc1_1 gpc3310 (
      {stage0_14[462]},
      {stage1_14[206]}
   );
   gpc1_1 gpc3311 (
      {stage0_14[463]},
      {stage1_14[207]}
   );
   gpc1_1 gpc3312 (
      {stage0_14[464]},
      {stage1_14[208]}
   );
   gpc1_1 gpc3313 (
      {stage0_14[465]},
      {stage1_14[209]}
   );
   gpc1_1 gpc3314 (
      {stage0_14[466]},
      {stage1_14[210]}
   );
   gpc1_1 gpc3315 (
      {stage0_14[467]},
      {stage1_14[211]}
   );
   gpc1_1 gpc3316 (
      {stage0_14[468]},
      {stage1_14[212]}
   );
   gpc1_1 gpc3317 (
      {stage0_14[469]},
      {stage1_14[213]}
   );
   gpc1_1 gpc3318 (
      {stage0_14[470]},
      {stage1_14[214]}
   );
   gpc1_1 gpc3319 (
      {stage0_14[471]},
      {stage1_14[215]}
   );
   gpc1_1 gpc3320 (
      {stage0_14[472]},
      {stage1_14[216]}
   );
   gpc1_1 gpc3321 (
      {stage0_14[473]},
      {stage1_14[217]}
   );
   gpc1_1 gpc3322 (
      {stage0_14[474]},
      {stage1_14[218]}
   );
   gpc1_1 gpc3323 (
      {stage0_14[475]},
      {stage1_14[219]}
   );
   gpc1_1 gpc3324 (
      {stage0_14[476]},
      {stage1_14[220]}
   );
   gpc1_1 gpc3325 (
      {stage0_14[477]},
      {stage1_14[221]}
   );
   gpc1_1 gpc3326 (
      {stage0_14[478]},
      {stage1_14[222]}
   );
   gpc1_1 gpc3327 (
      {stage0_14[479]},
      {stage1_14[223]}
   );
   gpc1_1 gpc3328 (
      {stage0_14[480]},
      {stage1_14[224]}
   );
   gpc1_1 gpc3329 (
      {stage0_14[481]},
      {stage1_14[225]}
   );
   gpc1_1 gpc3330 (
      {stage0_14[482]},
      {stage1_14[226]}
   );
   gpc1_1 gpc3331 (
      {stage0_14[483]},
      {stage1_14[227]}
   );
   gpc1_1 gpc3332 (
      {stage0_14[484]},
      {stage1_14[228]}
   );
   gpc1_1 gpc3333 (
      {stage0_14[485]},
      {stage1_14[229]}
   );
   gpc1_1 gpc3334 (
      {stage0_14[486]},
      {stage1_14[230]}
   );
   gpc1_1 gpc3335 (
      {stage0_14[487]},
      {stage1_14[231]}
   );
   gpc1_1 gpc3336 (
      {stage0_14[488]},
      {stage1_14[232]}
   );
   gpc1_1 gpc3337 (
      {stage0_14[489]},
      {stage1_14[233]}
   );
   gpc1_1 gpc3338 (
      {stage0_14[490]},
      {stage1_14[234]}
   );
   gpc1_1 gpc3339 (
      {stage0_14[491]},
      {stage1_14[235]}
   );
   gpc1_1 gpc3340 (
      {stage0_14[492]},
      {stage1_14[236]}
   );
   gpc1_1 gpc3341 (
      {stage0_14[493]},
      {stage1_14[237]}
   );
   gpc1_1 gpc3342 (
      {stage0_14[494]},
      {stage1_14[238]}
   );
   gpc1_1 gpc3343 (
      {stage0_14[495]},
      {stage1_14[239]}
   );
   gpc1_1 gpc3344 (
      {stage0_14[496]},
      {stage1_14[240]}
   );
   gpc1_1 gpc3345 (
      {stage0_14[497]},
      {stage1_14[241]}
   );
   gpc1_1 gpc3346 (
      {stage0_14[498]},
      {stage1_14[242]}
   );
   gpc1_1 gpc3347 (
      {stage0_14[499]},
      {stage1_14[243]}
   );
   gpc1_1 gpc3348 (
      {stage0_14[500]},
      {stage1_14[244]}
   );
   gpc1_1 gpc3349 (
      {stage0_14[501]},
      {stage1_14[245]}
   );
   gpc1_1 gpc3350 (
      {stage0_14[502]},
      {stage1_14[246]}
   );
   gpc1_1 gpc3351 (
      {stage0_14[503]},
      {stage1_14[247]}
   );
   gpc1_1 gpc3352 (
      {stage0_14[504]},
      {stage1_14[248]}
   );
   gpc1_1 gpc3353 (
      {stage0_14[505]},
      {stage1_14[249]}
   );
   gpc1_1 gpc3354 (
      {stage0_14[506]},
      {stage1_14[250]}
   );
   gpc1_1 gpc3355 (
      {stage0_14[507]},
      {stage1_14[251]}
   );
   gpc1_1 gpc3356 (
      {stage0_14[508]},
      {stage1_14[252]}
   );
   gpc1_1 gpc3357 (
      {stage0_14[509]},
      {stage1_14[253]}
   );
   gpc1_1 gpc3358 (
      {stage0_14[510]},
      {stage1_14[254]}
   );
   gpc1_1 gpc3359 (
      {stage0_14[511]},
      {stage1_14[255]}
   );
   gpc1_1 gpc3360 (
      {stage0_15[457]},
      {stage1_15[203]}
   );
   gpc1_1 gpc3361 (
      {stage0_15[458]},
      {stage1_15[204]}
   );
   gpc1_1 gpc3362 (
      {stage0_15[459]},
      {stage1_15[205]}
   );
   gpc1_1 gpc3363 (
      {stage0_15[460]},
      {stage1_15[206]}
   );
   gpc1_1 gpc3364 (
      {stage0_15[461]},
      {stage1_15[207]}
   );
   gpc1_1 gpc3365 (
      {stage0_15[462]},
      {stage1_15[208]}
   );
   gpc1_1 gpc3366 (
      {stage0_15[463]},
      {stage1_15[209]}
   );
   gpc1_1 gpc3367 (
      {stage0_15[464]},
      {stage1_15[210]}
   );
   gpc1_1 gpc3368 (
      {stage0_15[465]},
      {stage1_15[211]}
   );
   gpc1_1 gpc3369 (
      {stage0_15[466]},
      {stage1_15[212]}
   );
   gpc1_1 gpc3370 (
      {stage0_15[467]},
      {stage1_15[213]}
   );
   gpc1_1 gpc3371 (
      {stage0_15[468]},
      {stage1_15[214]}
   );
   gpc1_1 gpc3372 (
      {stage0_15[469]},
      {stage1_15[215]}
   );
   gpc1_1 gpc3373 (
      {stage0_15[470]},
      {stage1_15[216]}
   );
   gpc1_1 gpc3374 (
      {stage0_15[471]},
      {stage1_15[217]}
   );
   gpc1_1 gpc3375 (
      {stage0_15[472]},
      {stage1_15[218]}
   );
   gpc1_1 gpc3376 (
      {stage0_15[473]},
      {stage1_15[219]}
   );
   gpc1_1 gpc3377 (
      {stage0_15[474]},
      {stage1_15[220]}
   );
   gpc1_1 gpc3378 (
      {stage0_15[475]},
      {stage1_15[221]}
   );
   gpc1_1 gpc3379 (
      {stage0_15[476]},
      {stage1_15[222]}
   );
   gpc1_1 gpc3380 (
      {stage0_15[477]},
      {stage1_15[223]}
   );
   gpc1_1 gpc3381 (
      {stage0_15[478]},
      {stage1_15[224]}
   );
   gpc1_1 gpc3382 (
      {stage0_15[479]},
      {stage1_15[225]}
   );
   gpc1_1 gpc3383 (
      {stage0_15[480]},
      {stage1_15[226]}
   );
   gpc1_1 gpc3384 (
      {stage0_15[481]},
      {stage1_15[227]}
   );
   gpc1_1 gpc3385 (
      {stage0_15[482]},
      {stage1_15[228]}
   );
   gpc1_1 gpc3386 (
      {stage0_15[483]},
      {stage1_15[229]}
   );
   gpc1_1 gpc3387 (
      {stage0_15[484]},
      {stage1_15[230]}
   );
   gpc1_1 gpc3388 (
      {stage0_15[485]},
      {stage1_15[231]}
   );
   gpc1_1 gpc3389 (
      {stage0_15[486]},
      {stage1_15[232]}
   );
   gpc1_1 gpc3390 (
      {stage0_15[487]},
      {stage1_15[233]}
   );
   gpc1_1 gpc3391 (
      {stage0_15[488]},
      {stage1_15[234]}
   );
   gpc1_1 gpc3392 (
      {stage0_15[489]},
      {stage1_15[235]}
   );
   gpc1_1 gpc3393 (
      {stage0_15[490]},
      {stage1_15[236]}
   );
   gpc1_1 gpc3394 (
      {stage0_15[491]},
      {stage1_15[237]}
   );
   gpc1_1 gpc3395 (
      {stage0_15[492]},
      {stage1_15[238]}
   );
   gpc1_1 gpc3396 (
      {stage0_15[493]},
      {stage1_15[239]}
   );
   gpc1_1 gpc3397 (
      {stage0_15[494]},
      {stage1_15[240]}
   );
   gpc1_1 gpc3398 (
      {stage0_15[495]},
      {stage1_15[241]}
   );
   gpc1_1 gpc3399 (
      {stage0_15[496]},
      {stage1_15[242]}
   );
   gpc1_1 gpc3400 (
      {stage0_15[497]},
      {stage1_15[243]}
   );
   gpc1_1 gpc3401 (
      {stage0_15[498]},
      {stage1_15[244]}
   );
   gpc1_1 gpc3402 (
      {stage0_15[499]},
      {stage1_15[245]}
   );
   gpc1_1 gpc3403 (
      {stage0_15[500]},
      {stage1_15[246]}
   );
   gpc1_1 gpc3404 (
      {stage0_15[501]},
      {stage1_15[247]}
   );
   gpc1_1 gpc3405 (
      {stage0_15[502]},
      {stage1_15[248]}
   );
   gpc1_1 gpc3406 (
      {stage0_15[503]},
      {stage1_15[249]}
   );
   gpc1_1 gpc3407 (
      {stage0_15[504]},
      {stage1_15[250]}
   );
   gpc1_1 gpc3408 (
      {stage0_15[505]},
      {stage1_15[251]}
   );
   gpc1_1 gpc3409 (
      {stage0_15[506]},
      {stage1_15[252]}
   );
   gpc1_1 gpc3410 (
      {stage0_15[507]},
      {stage1_15[253]}
   );
   gpc1_1 gpc3411 (
      {stage0_15[508]},
      {stage1_15[254]}
   );
   gpc1_1 gpc3412 (
      {stage0_15[509]},
      {stage1_15[255]}
   );
   gpc1_1 gpc3413 (
      {stage0_15[510]},
      {stage1_15[256]}
   );
   gpc1_1 gpc3414 (
      {stage0_15[511]},
      {stage1_15[257]}
   );
   gpc1_1 gpc3415 (
      {stage0_17[492]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3416 (
      {stage0_17[493]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3417 (
      {stage0_17[494]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3418 (
      {stage0_17[495]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3419 (
      {stage0_17[496]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3420 (
      {stage0_17[497]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3421 (
      {stage0_17[498]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3422 (
      {stage0_17[499]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3423 (
      {stage0_17[500]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3424 (
      {stage0_17[501]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3425 (
      {stage0_17[502]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3426 (
      {stage0_17[503]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3427 (
      {stage0_17[504]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3428 (
      {stage0_17[505]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3429 (
      {stage0_17[506]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3430 (
      {stage0_17[507]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3431 (
      {stage0_17[508]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3432 (
      {stage0_17[509]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3433 (
      {stage0_17[510]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3434 (
      {stage0_17[511]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3435 (
      {stage0_18[434]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3436 (
      {stage0_18[435]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3437 (
      {stage0_18[436]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3438 (
      {stage0_18[437]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3439 (
      {stage0_18[438]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3440 (
      {stage0_18[439]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3441 (
      {stage0_18[440]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3442 (
      {stage0_18[441]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3443 (
      {stage0_18[442]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3444 (
      {stage0_18[443]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3445 (
      {stage0_18[444]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3446 (
      {stage0_18[445]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3447 (
      {stage0_18[446]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3448 (
      {stage0_18[447]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3449 (
      {stage0_18[448]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3450 (
      {stage0_18[449]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3451 (
      {stage0_18[450]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3452 (
      {stage0_18[451]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3453 (
      {stage0_18[452]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3454 (
      {stage0_18[453]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3455 (
      {stage0_18[454]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3456 (
      {stage0_18[455]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3457 (
      {stage0_18[456]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3458 (
      {stage0_18[457]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3459 (
      {stage0_18[458]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3460 (
      {stage0_18[459]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3461 (
      {stage0_18[460]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3462 (
      {stage0_18[461]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3463 (
      {stage0_18[462]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3464 (
      {stage0_18[463]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3465 (
      {stage0_18[464]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3466 (
      {stage0_18[465]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3467 (
      {stage0_18[466]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3468 (
      {stage0_18[467]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3469 (
      {stage0_18[468]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3470 (
      {stage0_18[469]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3471 (
      {stage0_18[470]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3472 (
      {stage0_18[471]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3473 (
      {stage0_18[472]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3474 (
      {stage0_18[473]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3475 (
      {stage0_18[474]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3476 (
      {stage0_18[475]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3477 (
      {stage0_18[476]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3478 (
      {stage0_18[477]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3479 (
      {stage0_18[478]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3480 (
      {stage0_18[479]},
      {stage1_18[209]}
   );
   gpc1_1 gpc3481 (
      {stage0_18[480]},
      {stage1_18[210]}
   );
   gpc1_1 gpc3482 (
      {stage0_18[481]},
      {stage1_18[211]}
   );
   gpc1_1 gpc3483 (
      {stage0_18[482]},
      {stage1_18[212]}
   );
   gpc1_1 gpc3484 (
      {stage0_18[483]},
      {stage1_18[213]}
   );
   gpc1_1 gpc3485 (
      {stage0_18[484]},
      {stage1_18[214]}
   );
   gpc1_1 gpc3486 (
      {stage0_18[485]},
      {stage1_18[215]}
   );
   gpc1_1 gpc3487 (
      {stage0_18[486]},
      {stage1_18[216]}
   );
   gpc1_1 gpc3488 (
      {stage0_18[487]},
      {stage1_18[217]}
   );
   gpc1_1 gpc3489 (
      {stage0_18[488]},
      {stage1_18[218]}
   );
   gpc1_1 gpc3490 (
      {stage0_18[489]},
      {stage1_18[219]}
   );
   gpc1_1 gpc3491 (
      {stage0_18[490]},
      {stage1_18[220]}
   );
   gpc1_1 gpc3492 (
      {stage0_18[491]},
      {stage1_18[221]}
   );
   gpc1_1 gpc3493 (
      {stage0_18[492]},
      {stage1_18[222]}
   );
   gpc1_1 gpc3494 (
      {stage0_18[493]},
      {stage1_18[223]}
   );
   gpc1_1 gpc3495 (
      {stage0_18[494]},
      {stage1_18[224]}
   );
   gpc1_1 gpc3496 (
      {stage0_18[495]},
      {stage1_18[225]}
   );
   gpc1_1 gpc3497 (
      {stage0_18[496]},
      {stage1_18[226]}
   );
   gpc1_1 gpc3498 (
      {stage0_18[497]},
      {stage1_18[227]}
   );
   gpc1_1 gpc3499 (
      {stage0_18[498]},
      {stage1_18[228]}
   );
   gpc1_1 gpc3500 (
      {stage0_18[499]},
      {stage1_18[229]}
   );
   gpc1_1 gpc3501 (
      {stage0_18[500]},
      {stage1_18[230]}
   );
   gpc1_1 gpc3502 (
      {stage0_18[501]},
      {stage1_18[231]}
   );
   gpc1_1 gpc3503 (
      {stage0_18[502]},
      {stage1_18[232]}
   );
   gpc1_1 gpc3504 (
      {stage0_18[503]},
      {stage1_18[233]}
   );
   gpc1_1 gpc3505 (
      {stage0_18[504]},
      {stage1_18[234]}
   );
   gpc1_1 gpc3506 (
      {stage0_18[505]},
      {stage1_18[235]}
   );
   gpc1_1 gpc3507 (
      {stage0_18[506]},
      {stage1_18[236]}
   );
   gpc1_1 gpc3508 (
      {stage0_18[507]},
      {stage1_18[237]}
   );
   gpc1_1 gpc3509 (
      {stage0_18[508]},
      {stage1_18[238]}
   );
   gpc1_1 gpc3510 (
      {stage0_18[509]},
      {stage1_18[239]}
   );
   gpc1_1 gpc3511 (
      {stage0_18[510]},
      {stage1_18[240]}
   );
   gpc1_1 gpc3512 (
      {stage0_18[511]},
      {stage1_18[241]}
   );
   gpc1_1 gpc3513 (
      {stage0_19[502]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3514 (
      {stage0_19[503]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3515 (
      {stage0_19[504]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3516 (
      {stage0_19[505]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3517 (
      {stage0_19[506]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3518 (
      {stage0_19[507]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3519 (
      {stage0_19[508]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3520 (
      {stage0_19[509]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3521 (
      {stage0_19[510]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3522 (
      {stage0_19[511]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3523 (
      {stage0_20[504]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3524 (
      {stage0_20[505]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3525 (
      {stage0_20[506]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3526 (
      {stage0_20[507]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3527 (
      {stage0_20[508]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3528 (
      {stage0_20[509]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3529 (
      {stage0_20[510]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3530 (
      {stage0_20[511]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3531 (
      {stage0_21[504]},
      {stage1_21[197]}
   );
   gpc1_1 gpc3532 (
      {stage0_21[505]},
      {stage1_21[198]}
   );
   gpc1_1 gpc3533 (
      {stage0_21[506]},
      {stage1_21[199]}
   );
   gpc1_1 gpc3534 (
      {stage0_21[507]},
      {stage1_21[200]}
   );
   gpc1_1 gpc3535 (
      {stage0_21[508]},
      {stage1_21[201]}
   );
   gpc1_1 gpc3536 (
      {stage0_21[509]},
      {stage1_21[202]}
   );
   gpc1_1 gpc3537 (
      {stage0_21[510]},
      {stage1_21[203]}
   );
   gpc1_1 gpc3538 (
      {stage0_21[511]},
      {stage1_21[204]}
   );
   gpc1_1 gpc3539 (
      {stage0_22[481]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3540 (
      {stage0_22[482]},
      {stage1_22[171]}
   );
   gpc1_1 gpc3541 (
      {stage0_22[483]},
      {stage1_22[172]}
   );
   gpc1_1 gpc3542 (
      {stage0_22[484]},
      {stage1_22[173]}
   );
   gpc1_1 gpc3543 (
      {stage0_22[485]},
      {stage1_22[174]}
   );
   gpc1_1 gpc3544 (
      {stage0_22[486]},
      {stage1_22[175]}
   );
   gpc1_1 gpc3545 (
      {stage0_22[487]},
      {stage1_22[176]}
   );
   gpc1_1 gpc3546 (
      {stage0_22[488]},
      {stage1_22[177]}
   );
   gpc1_1 gpc3547 (
      {stage0_22[489]},
      {stage1_22[178]}
   );
   gpc1_1 gpc3548 (
      {stage0_22[490]},
      {stage1_22[179]}
   );
   gpc1_1 gpc3549 (
      {stage0_22[491]},
      {stage1_22[180]}
   );
   gpc1_1 gpc3550 (
      {stage0_22[492]},
      {stage1_22[181]}
   );
   gpc1_1 gpc3551 (
      {stage0_22[493]},
      {stage1_22[182]}
   );
   gpc1_1 gpc3552 (
      {stage0_22[494]},
      {stage1_22[183]}
   );
   gpc1_1 gpc3553 (
      {stage0_22[495]},
      {stage1_22[184]}
   );
   gpc1_1 gpc3554 (
      {stage0_22[496]},
      {stage1_22[185]}
   );
   gpc1_1 gpc3555 (
      {stage0_22[497]},
      {stage1_22[186]}
   );
   gpc1_1 gpc3556 (
      {stage0_22[498]},
      {stage1_22[187]}
   );
   gpc1_1 gpc3557 (
      {stage0_22[499]},
      {stage1_22[188]}
   );
   gpc1_1 gpc3558 (
      {stage0_22[500]},
      {stage1_22[189]}
   );
   gpc1_1 gpc3559 (
      {stage0_22[501]},
      {stage1_22[190]}
   );
   gpc1_1 gpc3560 (
      {stage0_22[502]},
      {stage1_22[191]}
   );
   gpc1_1 gpc3561 (
      {stage0_22[503]},
      {stage1_22[192]}
   );
   gpc1_1 gpc3562 (
      {stage0_22[504]},
      {stage1_22[193]}
   );
   gpc1_1 gpc3563 (
      {stage0_22[505]},
      {stage1_22[194]}
   );
   gpc1_1 gpc3564 (
      {stage0_22[506]},
      {stage1_22[195]}
   );
   gpc1_1 gpc3565 (
      {stage0_22[507]},
      {stage1_22[196]}
   );
   gpc1_1 gpc3566 (
      {stage0_22[508]},
      {stage1_22[197]}
   );
   gpc1_1 gpc3567 (
      {stage0_22[509]},
      {stage1_22[198]}
   );
   gpc1_1 gpc3568 (
      {stage0_22[510]},
      {stage1_22[199]}
   );
   gpc1_1 gpc3569 (
      {stage0_22[511]},
      {stage1_22[200]}
   );
   gpc1_1 gpc3570 (
      {stage0_23[418]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3571 (
      {stage0_23[419]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3572 (
      {stage0_23[420]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3573 (
      {stage0_23[421]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3574 (
      {stage0_23[422]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3575 (
      {stage0_23[423]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3576 (
      {stage0_23[424]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3577 (
      {stage0_23[425]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3578 (
      {stage0_23[426]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3579 (
      {stage0_23[427]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3580 (
      {stage0_23[428]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3581 (
      {stage0_23[429]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3582 (
      {stage0_23[430]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3583 (
      {stage0_23[431]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3584 (
      {stage0_23[432]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3585 (
      {stage0_23[433]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3586 (
      {stage0_23[434]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3587 (
      {stage0_23[435]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3588 (
      {stage0_23[436]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3589 (
      {stage0_23[437]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3590 (
      {stage0_23[438]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3591 (
      {stage0_23[439]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3592 (
      {stage0_23[440]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3593 (
      {stage0_23[441]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3594 (
      {stage0_23[442]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3595 (
      {stage0_23[443]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3596 (
      {stage0_23[444]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3597 (
      {stage0_23[445]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3598 (
      {stage0_23[446]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3599 (
      {stage0_23[447]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3600 (
      {stage0_23[448]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3601 (
      {stage0_23[449]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3602 (
      {stage0_23[450]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3603 (
      {stage0_23[451]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3604 (
      {stage0_23[452]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3605 (
      {stage0_23[453]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3606 (
      {stage0_23[454]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3607 (
      {stage0_23[455]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3608 (
      {stage0_23[456]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3609 (
      {stage0_23[457]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3610 (
      {stage0_23[458]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3611 (
      {stage0_23[459]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3612 (
      {stage0_23[460]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3613 (
      {stage0_23[461]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3614 (
      {stage0_23[462]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3615 (
      {stage0_23[463]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3616 (
      {stage0_23[464]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3617 (
      {stage0_23[465]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3618 (
      {stage0_23[466]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3619 (
      {stage0_23[467]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3620 (
      {stage0_23[468]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3621 (
      {stage0_23[469]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3622 (
      {stage0_23[470]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3623 (
      {stage0_23[471]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3624 (
      {stage0_23[472]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3625 (
      {stage0_23[473]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3626 (
      {stage0_23[474]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3627 (
      {stage0_23[475]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3628 (
      {stage0_23[476]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3629 (
      {stage0_23[477]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3630 (
      {stage0_23[478]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3631 (
      {stage0_23[479]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3632 (
      {stage0_23[480]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3633 (
      {stage0_23[481]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3634 (
      {stage0_23[482]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3635 (
      {stage0_23[483]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3636 (
      {stage0_23[484]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3637 (
      {stage0_23[485]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3638 (
      {stage0_23[486]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3639 (
      {stage0_23[487]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3640 (
      {stage0_23[488]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3641 (
      {stage0_23[489]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3642 (
      {stage0_23[490]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3643 (
      {stage0_23[491]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3644 (
      {stage0_23[492]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3645 (
      {stage0_23[493]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3646 (
      {stage0_23[494]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3647 (
      {stage0_23[495]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3648 (
      {stage0_23[496]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3649 (
      {stage0_23[497]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3650 (
      {stage0_23[498]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3651 (
      {stage0_23[499]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3652 (
      {stage0_23[500]},
      {stage1_23[287]}
   );
   gpc1_1 gpc3653 (
      {stage0_23[501]},
      {stage1_23[288]}
   );
   gpc1_1 gpc3654 (
      {stage0_23[502]},
      {stage1_23[289]}
   );
   gpc1_1 gpc3655 (
      {stage0_23[503]},
      {stage1_23[290]}
   );
   gpc1_1 gpc3656 (
      {stage0_23[504]},
      {stage1_23[291]}
   );
   gpc1_1 gpc3657 (
      {stage0_23[505]},
      {stage1_23[292]}
   );
   gpc1_1 gpc3658 (
      {stage0_23[506]},
      {stage1_23[293]}
   );
   gpc1_1 gpc3659 (
      {stage0_23[507]},
      {stage1_23[294]}
   );
   gpc1_1 gpc3660 (
      {stage0_23[508]},
      {stage1_23[295]}
   );
   gpc1_1 gpc3661 (
      {stage0_23[509]},
      {stage1_23[296]}
   );
   gpc1_1 gpc3662 (
      {stage0_23[510]},
      {stage1_23[297]}
   );
   gpc1_1 gpc3663 (
      {stage0_23[511]},
      {stage1_23[298]}
   );
   gpc1_1 gpc3664 (
      {stage0_24[499]},
      {stage1_24[222]}
   );
   gpc1_1 gpc3665 (
      {stage0_24[500]},
      {stage1_24[223]}
   );
   gpc1_1 gpc3666 (
      {stage0_24[501]},
      {stage1_24[224]}
   );
   gpc1_1 gpc3667 (
      {stage0_24[502]},
      {stage1_24[225]}
   );
   gpc1_1 gpc3668 (
      {stage0_24[503]},
      {stage1_24[226]}
   );
   gpc1_1 gpc3669 (
      {stage0_24[504]},
      {stage1_24[227]}
   );
   gpc1_1 gpc3670 (
      {stage0_24[505]},
      {stage1_24[228]}
   );
   gpc1_1 gpc3671 (
      {stage0_24[506]},
      {stage1_24[229]}
   );
   gpc1_1 gpc3672 (
      {stage0_24[507]},
      {stage1_24[230]}
   );
   gpc1_1 gpc3673 (
      {stage0_24[508]},
      {stage1_24[231]}
   );
   gpc1_1 gpc3674 (
      {stage0_24[509]},
      {stage1_24[232]}
   );
   gpc1_1 gpc3675 (
      {stage0_24[510]},
      {stage1_24[233]}
   );
   gpc1_1 gpc3676 (
      {stage0_24[511]},
      {stage1_24[234]}
   );
   gpc1_1 gpc3677 (
      {stage0_25[506]},
      {stage1_25[205]}
   );
   gpc1_1 gpc3678 (
      {stage0_25[507]},
      {stage1_25[206]}
   );
   gpc1_1 gpc3679 (
      {stage0_25[508]},
      {stage1_25[207]}
   );
   gpc1_1 gpc3680 (
      {stage0_25[509]},
      {stage1_25[208]}
   );
   gpc1_1 gpc3681 (
      {stage0_25[510]},
      {stage1_25[209]}
   );
   gpc1_1 gpc3682 (
      {stage0_25[511]},
      {stage1_25[210]}
   );
   gpc1_1 gpc3683 (
      {stage0_26[503]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3684 (
      {stage0_26[504]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3685 (
      {stage0_26[505]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3686 (
      {stage0_26[506]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3687 (
      {stage0_26[507]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3688 (
      {stage0_26[508]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3689 (
      {stage0_26[509]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3690 (
      {stage0_26[510]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3691 (
      {stage0_26[511]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3692 (
      {stage0_27[503]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3693 (
      {stage0_27[504]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3694 (
      {stage0_27[505]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3695 (
      {stage0_27[506]},
      {stage1_27[206]}
   );
   gpc1_1 gpc3696 (
      {stage0_27[507]},
      {stage1_27[207]}
   );
   gpc1_1 gpc3697 (
      {stage0_27[508]},
      {stage1_27[208]}
   );
   gpc1_1 gpc3698 (
      {stage0_27[509]},
      {stage1_27[209]}
   );
   gpc1_1 gpc3699 (
      {stage0_27[510]},
      {stage1_27[210]}
   );
   gpc1_1 gpc3700 (
      {stage0_27[511]},
      {stage1_27[211]}
   );
   gpc1_1 gpc3701 (
      {stage0_28[500]},
      {stage1_28[237]}
   );
   gpc1_1 gpc3702 (
      {stage0_28[501]},
      {stage1_28[238]}
   );
   gpc1_1 gpc3703 (
      {stage0_28[502]},
      {stage1_28[239]}
   );
   gpc1_1 gpc3704 (
      {stage0_28[503]},
      {stage1_28[240]}
   );
   gpc1_1 gpc3705 (
      {stage0_28[504]},
      {stage1_28[241]}
   );
   gpc1_1 gpc3706 (
      {stage0_28[505]},
      {stage1_28[242]}
   );
   gpc1_1 gpc3707 (
      {stage0_28[506]},
      {stage1_28[243]}
   );
   gpc1_1 gpc3708 (
      {stage0_28[507]},
      {stage1_28[244]}
   );
   gpc1_1 gpc3709 (
      {stage0_28[508]},
      {stage1_28[245]}
   );
   gpc1_1 gpc3710 (
      {stage0_28[509]},
      {stage1_28[246]}
   );
   gpc1_1 gpc3711 (
      {stage0_28[510]},
      {stage1_28[247]}
   );
   gpc1_1 gpc3712 (
      {stage0_28[511]},
      {stage1_28[248]}
   );
   gpc1_1 gpc3713 (
      {stage0_29[510]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3714 (
      {stage0_29[511]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3715 (
      {stage0_30[443]},
      {stage1_30[164]}
   );
   gpc1_1 gpc3716 (
      {stage0_30[444]},
      {stage1_30[165]}
   );
   gpc1_1 gpc3717 (
      {stage0_30[445]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3718 (
      {stage0_30[446]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3719 (
      {stage0_30[447]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3720 (
      {stage0_30[448]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3721 (
      {stage0_30[449]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3722 (
      {stage0_30[450]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3723 (
      {stage0_30[451]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3724 (
      {stage0_30[452]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3725 (
      {stage0_30[453]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3726 (
      {stage0_30[454]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3727 (
      {stage0_30[455]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3728 (
      {stage0_30[456]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3729 (
      {stage0_30[457]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3730 (
      {stage0_30[458]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3731 (
      {stage0_30[459]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3732 (
      {stage0_30[460]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3733 (
      {stage0_30[461]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3734 (
      {stage0_30[462]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3735 (
      {stage0_30[463]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3736 (
      {stage0_30[464]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3737 (
      {stage0_30[465]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3738 (
      {stage0_30[466]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3739 (
      {stage0_30[467]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3740 (
      {stage0_30[468]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3741 (
      {stage0_30[469]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3742 (
      {stage0_30[470]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3743 (
      {stage0_30[471]},
      {stage1_30[192]}
   );
   gpc1_1 gpc3744 (
      {stage0_30[472]},
      {stage1_30[193]}
   );
   gpc1_1 gpc3745 (
      {stage0_30[473]},
      {stage1_30[194]}
   );
   gpc1_1 gpc3746 (
      {stage0_30[474]},
      {stage1_30[195]}
   );
   gpc1_1 gpc3747 (
      {stage0_30[475]},
      {stage1_30[196]}
   );
   gpc1_1 gpc3748 (
      {stage0_30[476]},
      {stage1_30[197]}
   );
   gpc1_1 gpc3749 (
      {stage0_30[477]},
      {stage1_30[198]}
   );
   gpc1_1 gpc3750 (
      {stage0_30[478]},
      {stage1_30[199]}
   );
   gpc1_1 gpc3751 (
      {stage0_30[479]},
      {stage1_30[200]}
   );
   gpc1_1 gpc3752 (
      {stage0_30[480]},
      {stage1_30[201]}
   );
   gpc1_1 gpc3753 (
      {stage0_30[481]},
      {stage1_30[202]}
   );
   gpc1_1 gpc3754 (
      {stage0_30[482]},
      {stage1_30[203]}
   );
   gpc1_1 gpc3755 (
      {stage0_30[483]},
      {stage1_30[204]}
   );
   gpc1_1 gpc3756 (
      {stage0_30[484]},
      {stage1_30[205]}
   );
   gpc1_1 gpc3757 (
      {stage0_30[485]},
      {stage1_30[206]}
   );
   gpc1_1 gpc3758 (
      {stage0_30[486]},
      {stage1_30[207]}
   );
   gpc1_1 gpc3759 (
      {stage0_30[487]},
      {stage1_30[208]}
   );
   gpc1_1 gpc3760 (
      {stage0_30[488]},
      {stage1_30[209]}
   );
   gpc1_1 gpc3761 (
      {stage0_30[489]},
      {stage1_30[210]}
   );
   gpc1_1 gpc3762 (
      {stage0_30[490]},
      {stage1_30[211]}
   );
   gpc1_1 gpc3763 (
      {stage0_30[491]},
      {stage1_30[212]}
   );
   gpc1_1 gpc3764 (
      {stage0_30[492]},
      {stage1_30[213]}
   );
   gpc1_1 gpc3765 (
      {stage0_30[493]},
      {stage1_30[214]}
   );
   gpc1_1 gpc3766 (
      {stage0_30[494]},
      {stage1_30[215]}
   );
   gpc1_1 gpc3767 (
      {stage0_30[495]},
      {stage1_30[216]}
   );
   gpc1_1 gpc3768 (
      {stage0_30[496]},
      {stage1_30[217]}
   );
   gpc1_1 gpc3769 (
      {stage0_30[497]},
      {stage1_30[218]}
   );
   gpc1_1 gpc3770 (
      {stage0_30[498]},
      {stage1_30[219]}
   );
   gpc1_1 gpc3771 (
      {stage0_30[499]},
      {stage1_30[220]}
   );
   gpc1_1 gpc3772 (
      {stage0_30[500]},
      {stage1_30[221]}
   );
   gpc1_1 gpc3773 (
      {stage0_30[501]},
      {stage1_30[222]}
   );
   gpc1_1 gpc3774 (
      {stage0_30[502]},
      {stage1_30[223]}
   );
   gpc1_1 gpc3775 (
      {stage0_30[503]},
      {stage1_30[224]}
   );
   gpc1_1 gpc3776 (
      {stage0_30[504]},
      {stage1_30[225]}
   );
   gpc1_1 gpc3777 (
      {stage0_30[505]},
      {stage1_30[226]}
   );
   gpc1_1 gpc3778 (
      {stage0_30[506]},
      {stage1_30[227]}
   );
   gpc1_1 gpc3779 (
      {stage0_30[507]},
      {stage1_30[228]}
   );
   gpc1_1 gpc3780 (
      {stage0_30[508]},
      {stage1_30[229]}
   );
   gpc1_1 gpc3781 (
      {stage0_30[509]},
      {stage1_30[230]}
   );
   gpc1_1 gpc3782 (
      {stage0_30[510]},
      {stage1_30[231]}
   );
   gpc1_1 gpc3783 (
      {stage0_30[511]},
      {stage1_30[232]}
   );
   gpc1_1 gpc3784 (
      {stage0_31[494]},
      {stage1_31[194]}
   );
   gpc1_1 gpc3785 (
      {stage0_31[495]},
      {stage1_31[195]}
   );
   gpc1_1 gpc3786 (
      {stage0_31[496]},
      {stage1_31[196]}
   );
   gpc1_1 gpc3787 (
      {stage0_31[497]},
      {stage1_31[197]}
   );
   gpc1_1 gpc3788 (
      {stage0_31[498]},
      {stage1_31[198]}
   );
   gpc1_1 gpc3789 (
      {stage0_31[499]},
      {stage1_31[199]}
   );
   gpc1_1 gpc3790 (
      {stage0_31[500]},
      {stage1_31[200]}
   );
   gpc1_1 gpc3791 (
      {stage0_31[501]},
      {stage1_31[201]}
   );
   gpc1_1 gpc3792 (
      {stage0_31[502]},
      {stage1_31[202]}
   );
   gpc1_1 gpc3793 (
      {stage0_31[503]},
      {stage1_31[203]}
   );
   gpc1_1 gpc3794 (
      {stage0_31[504]},
      {stage1_31[204]}
   );
   gpc1_1 gpc3795 (
      {stage0_31[505]},
      {stage1_31[205]}
   );
   gpc1_1 gpc3796 (
      {stage0_31[506]},
      {stage1_31[206]}
   );
   gpc1_1 gpc3797 (
      {stage0_31[507]},
      {stage1_31[207]}
   );
   gpc1_1 gpc3798 (
      {stage0_31[508]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3799 (
      {stage0_31[509]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3800 (
      {stage0_31[510]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3801 (
      {stage0_31[511]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3802 (
      {stage0_32[303]},
      {stage1_32[206]}
   );
   gpc1_1 gpc3803 (
      {stage0_32[304]},
      {stage1_32[207]}
   );
   gpc1_1 gpc3804 (
      {stage0_32[305]},
      {stage1_32[208]}
   );
   gpc1_1 gpc3805 (
      {stage0_32[306]},
      {stage1_32[209]}
   );
   gpc1_1 gpc3806 (
      {stage0_32[307]},
      {stage1_32[210]}
   );
   gpc1_1 gpc3807 (
      {stage0_32[308]},
      {stage1_32[211]}
   );
   gpc1_1 gpc3808 (
      {stage0_32[309]},
      {stage1_32[212]}
   );
   gpc1_1 gpc3809 (
      {stage0_32[310]},
      {stage1_32[213]}
   );
   gpc1_1 gpc3810 (
      {stage0_32[311]},
      {stage1_32[214]}
   );
   gpc1_1 gpc3811 (
      {stage0_32[312]},
      {stage1_32[215]}
   );
   gpc1_1 gpc3812 (
      {stage0_32[313]},
      {stage1_32[216]}
   );
   gpc1_1 gpc3813 (
      {stage0_32[314]},
      {stage1_32[217]}
   );
   gpc1_1 gpc3814 (
      {stage0_32[315]},
      {stage1_32[218]}
   );
   gpc1_1 gpc3815 (
      {stage0_32[316]},
      {stage1_32[219]}
   );
   gpc1_1 gpc3816 (
      {stage0_32[317]},
      {stage1_32[220]}
   );
   gpc1_1 gpc3817 (
      {stage0_32[318]},
      {stage1_32[221]}
   );
   gpc1_1 gpc3818 (
      {stage0_32[319]},
      {stage1_32[222]}
   );
   gpc1_1 gpc3819 (
      {stage0_32[320]},
      {stage1_32[223]}
   );
   gpc1_1 gpc3820 (
      {stage0_32[321]},
      {stage1_32[224]}
   );
   gpc1_1 gpc3821 (
      {stage0_32[322]},
      {stage1_32[225]}
   );
   gpc1_1 gpc3822 (
      {stage0_32[323]},
      {stage1_32[226]}
   );
   gpc1_1 gpc3823 (
      {stage0_32[324]},
      {stage1_32[227]}
   );
   gpc1_1 gpc3824 (
      {stage0_32[325]},
      {stage1_32[228]}
   );
   gpc1_1 gpc3825 (
      {stage0_32[326]},
      {stage1_32[229]}
   );
   gpc1_1 gpc3826 (
      {stage0_32[327]},
      {stage1_32[230]}
   );
   gpc1_1 gpc3827 (
      {stage0_32[328]},
      {stage1_32[231]}
   );
   gpc1_1 gpc3828 (
      {stage0_32[329]},
      {stage1_32[232]}
   );
   gpc1_1 gpc3829 (
      {stage0_32[330]},
      {stage1_32[233]}
   );
   gpc1_1 gpc3830 (
      {stage0_32[331]},
      {stage1_32[234]}
   );
   gpc1_1 gpc3831 (
      {stage0_32[332]},
      {stage1_32[235]}
   );
   gpc1_1 gpc3832 (
      {stage0_32[333]},
      {stage1_32[236]}
   );
   gpc1_1 gpc3833 (
      {stage0_32[334]},
      {stage1_32[237]}
   );
   gpc1_1 gpc3834 (
      {stage0_32[335]},
      {stage1_32[238]}
   );
   gpc1_1 gpc3835 (
      {stage0_32[336]},
      {stage1_32[239]}
   );
   gpc1_1 gpc3836 (
      {stage0_32[337]},
      {stage1_32[240]}
   );
   gpc1_1 gpc3837 (
      {stage0_32[338]},
      {stage1_32[241]}
   );
   gpc1_1 gpc3838 (
      {stage0_32[339]},
      {stage1_32[242]}
   );
   gpc1_1 gpc3839 (
      {stage0_32[340]},
      {stage1_32[243]}
   );
   gpc1_1 gpc3840 (
      {stage0_32[341]},
      {stage1_32[244]}
   );
   gpc1_1 gpc3841 (
      {stage0_32[342]},
      {stage1_32[245]}
   );
   gpc1_1 gpc3842 (
      {stage0_32[343]},
      {stage1_32[246]}
   );
   gpc1_1 gpc3843 (
      {stage0_32[344]},
      {stage1_32[247]}
   );
   gpc1_1 gpc3844 (
      {stage0_32[345]},
      {stage1_32[248]}
   );
   gpc1_1 gpc3845 (
      {stage0_32[346]},
      {stage1_32[249]}
   );
   gpc1_1 gpc3846 (
      {stage0_32[347]},
      {stage1_32[250]}
   );
   gpc1_1 gpc3847 (
      {stage0_32[348]},
      {stage1_32[251]}
   );
   gpc1_1 gpc3848 (
      {stage0_32[349]},
      {stage1_32[252]}
   );
   gpc1_1 gpc3849 (
      {stage0_32[350]},
      {stage1_32[253]}
   );
   gpc1_1 gpc3850 (
      {stage0_32[351]},
      {stage1_32[254]}
   );
   gpc1_1 gpc3851 (
      {stage0_32[352]},
      {stage1_32[255]}
   );
   gpc1_1 gpc3852 (
      {stage0_32[353]},
      {stage1_32[256]}
   );
   gpc1_1 gpc3853 (
      {stage0_32[354]},
      {stage1_32[257]}
   );
   gpc1_1 gpc3854 (
      {stage0_32[355]},
      {stage1_32[258]}
   );
   gpc1_1 gpc3855 (
      {stage0_32[356]},
      {stage1_32[259]}
   );
   gpc1_1 gpc3856 (
      {stage0_32[357]},
      {stage1_32[260]}
   );
   gpc1_1 gpc3857 (
      {stage0_32[358]},
      {stage1_32[261]}
   );
   gpc1_1 gpc3858 (
      {stage0_32[359]},
      {stage1_32[262]}
   );
   gpc1_1 gpc3859 (
      {stage0_32[360]},
      {stage1_32[263]}
   );
   gpc1_1 gpc3860 (
      {stage0_32[361]},
      {stage1_32[264]}
   );
   gpc1_1 gpc3861 (
      {stage0_32[362]},
      {stage1_32[265]}
   );
   gpc1_1 gpc3862 (
      {stage0_32[363]},
      {stage1_32[266]}
   );
   gpc1_1 gpc3863 (
      {stage0_32[364]},
      {stage1_32[267]}
   );
   gpc1_1 gpc3864 (
      {stage0_32[365]},
      {stage1_32[268]}
   );
   gpc1_1 gpc3865 (
      {stage0_32[366]},
      {stage1_32[269]}
   );
   gpc1_1 gpc3866 (
      {stage0_32[367]},
      {stage1_32[270]}
   );
   gpc1_1 gpc3867 (
      {stage0_32[368]},
      {stage1_32[271]}
   );
   gpc1_1 gpc3868 (
      {stage0_32[369]},
      {stage1_32[272]}
   );
   gpc1_1 gpc3869 (
      {stage0_32[370]},
      {stage1_32[273]}
   );
   gpc1_1 gpc3870 (
      {stage0_32[371]},
      {stage1_32[274]}
   );
   gpc1_1 gpc3871 (
      {stage0_32[372]},
      {stage1_32[275]}
   );
   gpc1_1 gpc3872 (
      {stage0_32[373]},
      {stage1_32[276]}
   );
   gpc1_1 gpc3873 (
      {stage0_32[374]},
      {stage1_32[277]}
   );
   gpc1_1 gpc3874 (
      {stage0_32[375]},
      {stage1_32[278]}
   );
   gpc1_1 gpc3875 (
      {stage0_32[376]},
      {stage1_32[279]}
   );
   gpc1_1 gpc3876 (
      {stage0_32[377]},
      {stage1_32[280]}
   );
   gpc1_1 gpc3877 (
      {stage0_32[378]},
      {stage1_32[281]}
   );
   gpc1_1 gpc3878 (
      {stage0_32[379]},
      {stage1_32[282]}
   );
   gpc1_1 gpc3879 (
      {stage0_32[380]},
      {stage1_32[283]}
   );
   gpc1_1 gpc3880 (
      {stage0_32[381]},
      {stage1_32[284]}
   );
   gpc1_1 gpc3881 (
      {stage0_32[382]},
      {stage1_32[285]}
   );
   gpc1_1 gpc3882 (
      {stage0_32[383]},
      {stage1_32[286]}
   );
   gpc1_1 gpc3883 (
      {stage0_32[384]},
      {stage1_32[287]}
   );
   gpc1_1 gpc3884 (
      {stage0_32[385]},
      {stage1_32[288]}
   );
   gpc1_1 gpc3885 (
      {stage0_32[386]},
      {stage1_32[289]}
   );
   gpc1_1 gpc3886 (
      {stage0_32[387]},
      {stage1_32[290]}
   );
   gpc1_1 gpc3887 (
      {stage0_32[388]},
      {stage1_32[291]}
   );
   gpc1_1 gpc3888 (
      {stage0_32[389]},
      {stage1_32[292]}
   );
   gpc1_1 gpc3889 (
      {stage0_32[390]},
      {stage1_32[293]}
   );
   gpc1_1 gpc3890 (
      {stage0_32[391]},
      {stage1_32[294]}
   );
   gpc1_1 gpc3891 (
      {stage0_32[392]},
      {stage1_32[295]}
   );
   gpc1_1 gpc3892 (
      {stage0_32[393]},
      {stage1_32[296]}
   );
   gpc1_1 gpc3893 (
      {stage0_32[394]},
      {stage1_32[297]}
   );
   gpc1_1 gpc3894 (
      {stage0_32[395]},
      {stage1_32[298]}
   );
   gpc1_1 gpc3895 (
      {stage0_32[396]},
      {stage1_32[299]}
   );
   gpc1_1 gpc3896 (
      {stage0_32[397]},
      {stage1_32[300]}
   );
   gpc1_1 gpc3897 (
      {stage0_32[398]},
      {stage1_32[301]}
   );
   gpc1_1 gpc3898 (
      {stage0_32[399]},
      {stage1_32[302]}
   );
   gpc1_1 gpc3899 (
      {stage0_32[400]},
      {stage1_32[303]}
   );
   gpc1_1 gpc3900 (
      {stage0_32[401]},
      {stage1_32[304]}
   );
   gpc1_1 gpc3901 (
      {stage0_32[402]},
      {stage1_32[305]}
   );
   gpc1_1 gpc3902 (
      {stage0_32[403]},
      {stage1_32[306]}
   );
   gpc1_1 gpc3903 (
      {stage0_32[404]},
      {stage1_32[307]}
   );
   gpc1_1 gpc3904 (
      {stage0_32[405]},
      {stage1_32[308]}
   );
   gpc1_1 gpc3905 (
      {stage0_32[406]},
      {stage1_32[309]}
   );
   gpc1_1 gpc3906 (
      {stage0_32[407]},
      {stage1_32[310]}
   );
   gpc1_1 gpc3907 (
      {stage0_32[408]},
      {stage1_32[311]}
   );
   gpc1_1 gpc3908 (
      {stage0_32[409]},
      {stage1_32[312]}
   );
   gpc1_1 gpc3909 (
      {stage0_32[410]},
      {stage1_32[313]}
   );
   gpc1_1 gpc3910 (
      {stage0_32[411]},
      {stage1_32[314]}
   );
   gpc1_1 gpc3911 (
      {stage0_32[412]},
      {stage1_32[315]}
   );
   gpc1_1 gpc3912 (
      {stage0_32[413]},
      {stage1_32[316]}
   );
   gpc1_1 gpc3913 (
      {stage0_32[414]},
      {stage1_32[317]}
   );
   gpc1_1 gpc3914 (
      {stage0_32[415]},
      {stage1_32[318]}
   );
   gpc1_1 gpc3915 (
      {stage0_32[416]},
      {stage1_32[319]}
   );
   gpc1_1 gpc3916 (
      {stage0_32[417]},
      {stage1_32[320]}
   );
   gpc1_1 gpc3917 (
      {stage0_32[418]},
      {stage1_32[321]}
   );
   gpc1_1 gpc3918 (
      {stage0_32[419]},
      {stage1_32[322]}
   );
   gpc1_1 gpc3919 (
      {stage0_32[420]},
      {stage1_32[323]}
   );
   gpc1_1 gpc3920 (
      {stage0_32[421]},
      {stage1_32[324]}
   );
   gpc1_1 gpc3921 (
      {stage0_32[422]},
      {stage1_32[325]}
   );
   gpc1_1 gpc3922 (
      {stage0_32[423]},
      {stage1_32[326]}
   );
   gpc1_1 gpc3923 (
      {stage0_32[424]},
      {stage1_32[327]}
   );
   gpc1_1 gpc3924 (
      {stage0_32[425]},
      {stage1_32[328]}
   );
   gpc1_1 gpc3925 (
      {stage0_32[426]},
      {stage1_32[329]}
   );
   gpc1_1 gpc3926 (
      {stage0_32[427]},
      {stage1_32[330]}
   );
   gpc1_1 gpc3927 (
      {stage0_32[428]},
      {stage1_32[331]}
   );
   gpc1_1 gpc3928 (
      {stage0_32[429]},
      {stage1_32[332]}
   );
   gpc1_1 gpc3929 (
      {stage0_32[430]},
      {stage1_32[333]}
   );
   gpc1_1 gpc3930 (
      {stage0_32[431]},
      {stage1_32[334]}
   );
   gpc1_1 gpc3931 (
      {stage0_32[432]},
      {stage1_32[335]}
   );
   gpc1_1 gpc3932 (
      {stage0_32[433]},
      {stage1_32[336]}
   );
   gpc1_1 gpc3933 (
      {stage0_32[434]},
      {stage1_32[337]}
   );
   gpc1_1 gpc3934 (
      {stage0_32[435]},
      {stage1_32[338]}
   );
   gpc1_1 gpc3935 (
      {stage0_32[436]},
      {stage1_32[339]}
   );
   gpc1_1 gpc3936 (
      {stage0_32[437]},
      {stage1_32[340]}
   );
   gpc1_1 gpc3937 (
      {stage0_32[438]},
      {stage1_32[341]}
   );
   gpc1_1 gpc3938 (
      {stage0_32[439]},
      {stage1_32[342]}
   );
   gpc1_1 gpc3939 (
      {stage0_32[440]},
      {stage1_32[343]}
   );
   gpc1_1 gpc3940 (
      {stage0_32[441]},
      {stage1_32[344]}
   );
   gpc1_1 gpc3941 (
      {stage0_32[442]},
      {stage1_32[345]}
   );
   gpc1_1 gpc3942 (
      {stage0_32[443]},
      {stage1_32[346]}
   );
   gpc1_1 gpc3943 (
      {stage0_32[444]},
      {stage1_32[347]}
   );
   gpc1_1 gpc3944 (
      {stage0_32[445]},
      {stage1_32[348]}
   );
   gpc1_1 gpc3945 (
      {stage0_32[446]},
      {stage1_32[349]}
   );
   gpc1_1 gpc3946 (
      {stage0_32[447]},
      {stage1_32[350]}
   );
   gpc1_1 gpc3947 (
      {stage0_32[448]},
      {stage1_32[351]}
   );
   gpc1_1 gpc3948 (
      {stage0_32[449]},
      {stage1_32[352]}
   );
   gpc1_1 gpc3949 (
      {stage0_32[450]},
      {stage1_32[353]}
   );
   gpc1_1 gpc3950 (
      {stage0_32[451]},
      {stage1_32[354]}
   );
   gpc1_1 gpc3951 (
      {stage0_32[452]},
      {stage1_32[355]}
   );
   gpc1_1 gpc3952 (
      {stage0_32[453]},
      {stage1_32[356]}
   );
   gpc1_1 gpc3953 (
      {stage0_32[454]},
      {stage1_32[357]}
   );
   gpc1_1 gpc3954 (
      {stage0_32[455]},
      {stage1_32[358]}
   );
   gpc1_1 gpc3955 (
      {stage0_32[456]},
      {stage1_32[359]}
   );
   gpc1_1 gpc3956 (
      {stage0_32[457]},
      {stage1_32[360]}
   );
   gpc1_1 gpc3957 (
      {stage0_32[458]},
      {stage1_32[361]}
   );
   gpc1_1 gpc3958 (
      {stage0_32[459]},
      {stage1_32[362]}
   );
   gpc1_1 gpc3959 (
      {stage0_32[460]},
      {stage1_32[363]}
   );
   gpc1_1 gpc3960 (
      {stage0_32[461]},
      {stage1_32[364]}
   );
   gpc1_1 gpc3961 (
      {stage0_32[462]},
      {stage1_32[365]}
   );
   gpc1_1 gpc3962 (
      {stage0_32[463]},
      {stage1_32[366]}
   );
   gpc1_1 gpc3963 (
      {stage0_32[464]},
      {stage1_32[367]}
   );
   gpc1_1 gpc3964 (
      {stage0_32[465]},
      {stage1_32[368]}
   );
   gpc1_1 gpc3965 (
      {stage0_32[466]},
      {stage1_32[369]}
   );
   gpc1_1 gpc3966 (
      {stage0_32[467]},
      {stage1_32[370]}
   );
   gpc1_1 gpc3967 (
      {stage0_32[468]},
      {stage1_32[371]}
   );
   gpc1_1 gpc3968 (
      {stage0_32[469]},
      {stage1_32[372]}
   );
   gpc1_1 gpc3969 (
      {stage0_32[470]},
      {stage1_32[373]}
   );
   gpc1_1 gpc3970 (
      {stage0_32[471]},
      {stage1_32[374]}
   );
   gpc1_1 gpc3971 (
      {stage0_32[472]},
      {stage1_32[375]}
   );
   gpc1_1 gpc3972 (
      {stage0_32[473]},
      {stage1_32[376]}
   );
   gpc1_1 gpc3973 (
      {stage0_32[474]},
      {stage1_32[377]}
   );
   gpc1_1 gpc3974 (
      {stage0_32[475]},
      {stage1_32[378]}
   );
   gpc1_1 gpc3975 (
      {stage0_32[476]},
      {stage1_32[379]}
   );
   gpc1_1 gpc3976 (
      {stage0_32[477]},
      {stage1_32[380]}
   );
   gpc1_1 gpc3977 (
      {stage0_32[478]},
      {stage1_32[381]}
   );
   gpc1_1 gpc3978 (
      {stage0_32[479]},
      {stage1_32[382]}
   );
   gpc1_1 gpc3979 (
      {stage0_32[480]},
      {stage1_32[383]}
   );
   gpc1_1 gpc3980 (
      {stage0_32[481]},
      {stage1_32[384]}
   );
   gpc1_1 gpc3981 (
      {stage0_32[482]},
      {stage1_32[385]}
   );
   gpc1_1 gpc3982 (
      {stage0_32[483]},
      {stage1_32[386]}
   );
   gpc1_1 gpc3983 (
      {stage0_32[484]},
      {stage1_32[387]}
   );
   gpc1_1 gpc3984 (
      {stage0_32[485]},
      {stage1_32[388]}
   );
   gpc1_1 gpc3985 (
      {stage0_32[486]},
      {stage1_32[389]}
   );
   gpc1_1 gpc3986 (
      {stage0_32[487]},
      {stage1_32[390]}
   );
   gpc1_1 gpc3987 (
      {stage0_32[488]},
      {stage1_32[391]}
   );
   gpc1_1 gpc3988 (
      {stage0_32[489]},
      {stage1_32[392]}
   );
   gpc1_1 gpc3989 (
      {stage0_32[490]},
      {stage1_32[393]}
   );
   gpc1_1 gpc3990 (
      {stage0_32[491]},
      {stage1_32[394]}
   );
   gpc1_1 gpc3991 (
      {stage0_32[492]},
      {stage1_32[395]}
   );
   gpc1_1 gpc3992 (
      {stage0_32[493]},
      {stage1_32[396]}
   );
   gpc1_1 gpc3993 (
      {stage0_32[494]},
      {stage1_32[397]}
   );
   gpc1_1 gpc3994 (
      {stage0_32[495]},
      {stage1_32[398]}
   );
   gpc1_1 gpc3995 (
      {stage0_32[496]},
      {stage1_32[399]}
   );
   gpc1_1 gpc3996 (
      {stage0_32[497]},
      {stage1_32[400]}
   );
   gpc1_1 gpc3997 (
      {stage0_32[498]},
      {stage1_32[401]}
   );
   gpc1_1 gpc3998 (
      {stage0_32[499]},
      {stage1_32[402]}
   );
   gpc1_1 gpc3999 (
      {stage0_32[500]},
      {stage1_32[403]}
   );
   gpc1_1 gpc4000 (
      {stage0_32[501]},
      {stage1_32[404]}
   );
   gpc1_1 gpc4001 (
      {stage0_32[502]},
      {stage1_32[405]}
   );
   gpc1_1 gpc4002 (
      {stage0_32[503]},
      {stage1_32[406]}
   );
   gpc1_1 gpc4003 (
      {stage0_32[504]},
      {stage1_32[407]}
   );
   gpc1_1 gpc4004 (
      {stage0_32[505]},
      {stage1_32[408]}
   );
   gpc1_1 gpc4005 (
      {stage0_32[506]},
      {stage1_32[409]}
   );
   gpc1_1 gpc4006 (
      {stage0_32[507]},
      {stage1_32[410]}
   );
   gpc1_1 gpc4007 (
      {stage0_32[508]},
      {stage1_32[411]}
   );
   gpc1_1 gpc4008 (
      {stage0_32[509]},
      {stage1_32[412]}
   );
   gpc1_1 gpc4009 (
      {stage0_32[510]},
      {stage1_32[413]}
   );
   gpc1_1 gpc4010 (
      {stage0_32[511]},
      {stage1_32[414]}
   );
   gpc1_1 gpc4011 (
      {stage0_33[491]},
      {stage1_33[189]}
   );
   gpc1_1 gpc4012 (
      {stage0_33[492]},
      {stage1_33[190]}
   );
   gpc1_1 gpc4013 (
      {stage0_33[493]},
      {stage1_33[191]}
   );
   gpc1_1 gpc4014 (
      {stage0_33[494]},
      {stage1_33[192]}
   );
   gpc1_1 gpc4015 (
      {stage0_33[495]},
      {stage1_33[193]}
   );
   gpc1_1 gpc4016 (
      {stage0_33[496]},
      {stage1_33[194]}
   );
   gpc1_1 gpc4017 (
      {stage0_33[497]},
      {stage1_33[195]}
   );
   gpc1_1 gpc4018 (
      {stage0_33[498]},
      {stage1_33[196]}
   );
   gpc1_1 gpc4019 (
      {stage0_33[499]},
      {stage1_33[197]}
   );
   gpc1_1 gpc4020 (
      {stage0_33[500]},
      {stage1_33[198]}
   );
   gpc1_1 gpc4021 (
      {stage0_33[501]},
      {stage1_33[199]}
   );
   gpc1_1 gpc4022 (
      {stage0_33[502]},
      {stage1_33[200]}
   );
   gpc1_1 gpc4023 (
      {stage0_33[503]},
      {stage1_33[201]}
   );
   gpc1_1 gpc4024 (
      {stage0_33[504]},
      {stage1_33[202]}
   );
   gpc1_1 gpc4025 (
      {stage0_33[505]},
      {stage1_33[203]}
   );
   gpc1_1 gpc4026 (
      {stage0_33[506]},
      {stage1_33[204]}
   );
   gpc1_1 gpc4027 (
      {stage0_33[507]},
      {stage1_33[205]}
   );
   gpc1_1 gpc4028 (
      {stage0_33[508]},
      {stage1_33[206]}
   );
   gpc1_1 gpc4029 (
      {stage0_33[509]},
      {stage1_33[207]}
   );
   gpc1_1 gpc4030 (
      {stage0_33[510]},
      {stage1_33[208]}
   );
   gpc1_1 gpc4031 (
      {stage0_33[511]},
      {stage1_33[209]}
   );
   gpc1_1 gpc4032 (
      {stage0_34[396]},
      {stage1_34[152]}
   );
   gpc1_1 gpc4033 (
      {stage0_34[397]},
      {stage1_34[153]}
   );
   gpc1_1 gpc4034 (
      {stage0_34[398]},
      {stage1_34[154]}
   );
   gpc1_1 gpc4035 (
      {stage0_34[399]},
      {stage1_34[155]}
   );
   gpc1_1 gpc4036 (
      {stage0_34[400]},
      {stage1_34[156]}
   );
   gpc1_1 gpc4037 (
      {stage0_34[401]},
      {stage1_34[157]}
   );
   gpc1_1 gpc4038 (
      {stage0_34[402]},
      {stage1_34[158]}
   );
   gpc1_1 gpc4039 (
      {stage0_34[403]},
      {stage1_34[159]}
   );
   gpc1_1 gpc4040 (
      {stage0_34[404]},
      {stage1_34[160]}
   );
   gpc1_1 gpc4041 (
      {stage0_34[405]},
      {stage1_34[161]}
   );
   gpc1_1 gpc4042 (
      {stage0_34[406]},
      {stage1_34[162]}
   );
   gpc1_1 gpc4043 (
      {stage0_34[407]},
      {stage1_34[163]}
   );
   gpc1_1 gpc4044 (
      {stage0_34[408]},
      {stage1_34[164]}
   );
   gpc1_1 gpc4045 (
      {stage0_34[409]},
      {stage1_34[165]}
   );
   gpc1_1 gpc4046 (
      {stage0_34[410]},
      {stage1_34[166]}
   );
   gpc1_1 gpc4047 (
      {stage0_34[411]},
      {stage1_34[167]}
   );
   gpc1_1 gpc4048 (
      {stage0_34[412]},
      {stage1_34[168]}
   );
   gpc1_1 gpc4049 (
      {stage0_34[413]},
      {stage1_34[169]}
   );
   gpc1_1 gpc4050 (
      {stage0_34[414]},
      {stage1_34[170]}
   );
   gpc1_1 gpc4051 (
      {stage0_34[415]},
      {stage1_34[171]}
   );
   gpc1_1 gpc4052 (
      {stage0_34[416]},
      {stage1_34[172]}
   );
   gpc1_1 gpc4053 (
      {stage0_34[417]},
      {stage1_34[173]}
   );
   gpc1_1 gpc4054 (
      {stage0_34[418]},
      {stage1_34[174]}
   );
   gpc1_1 gpc4055 (
      {stage0_34[419]},
      {stage1_34[175]}
   );
   gpc1_1 gpc4056 (
      {stage0_34[420]},
      {stage1_34[176]}
   );
   gpc1_1 gpc4057 (
      {stage0_34[421]},
      {stage1_34[177]}
   );
   gpc1_1 gpc4058 (
      {stage0_34[422]},
      {stage1_34[178]}
   );
   gpc1_1 gpc4059 (
      {stage0_34[423]},
      {stage1_34[179]}
   );
   gpc1_1 gpc4060 (
      {stage0_34[424]},
      {stage1_34[180]}
   );
   gpc1_1 gpc4061 (
      {stage0_34[425]},
      {stage1_34[181]}
   );
   gpc1_1 gpc4062 (
      {stage0_34[426]},
      {stage1_34[182]}
   );
   gpc1_1 gpc4063 (
      {stage0_34[427]},
      {stage1_34[183]}
   );
   gpc1_1 gpc4064 (
      {stage0_34[428]},
      {stage1_34[184]}
   );
   gpc1_1 gpc4065 (
      {stage0_34[429]},
      {stage1_34[185]}
   );
   gpc1_1 gpc4066 (
      {stage0_34[430]},
      {stage1_34[186]}
   );
   gpc1_1 gpc4067 (
      {stage0_34[431]},
      {stage1_34[187]}
   );
   gpc1_1 gpc4068 (
      {stage0_34[432]},
      {stage1_34[188]}
   );
   gpc1_1 gpc4069 (
      {stage0_34[433]},
      {stage1_34[189]}
   );
   gpc1_1 gpc4070 (
      {stage0_34[434]},
      {stage1_34[190]}
   );
   gpc1_1 gpc4071 (
      {stage0_34[435]},
      {stage1_34[191]}
   );
   gpc1_1 gpc4072 (
      {stage0_34[436]},
      {stage1_34[192]}
   );
   gpc1_1 gpc4073 (
      {stage0_34[437]},
      {stage1_34[193]}
   );
   gpc1_1 gpc4074 (
      {stage0_34[438]},
      {stage1_34[194]}
   );
   gpc1_1 gpc4075 (
      {stage0_34[439]},
      {stage1_34[195]}
   );
   gpc1_1 gpc4076 (
      {stage0_34[440]},
      {stage1_34[196]}
   );
   gpc1_1 gpc4077 (
      {stage0_34[441]},
      {stage1_34[197]}
   );
   gpc1_1 gpc4078 (
      {stage0_34[442]},
      {stage1_34[198]}
   );
   gpc1_1 gpc4079 (
      {stage0_34[443]},
      {stage1_34[199]}
   );
   gpc1_1 gpc4080 (
      {stage0_34[444]},
      {stage1_34[200]}
   );
   gpc1_1 gpc4081 (
      {stage0_34[445]},
      {stage1_34[201]}
   );
   gpc1_1 gpc4082 (
      {stage0_34[446]},
      {stage1_34[202]}
   );
   gpc1_1 gpc4083 (
      {stage0_34[447]},
      {stage1_34[203]}
   );
   gpc1_1 gpc4084 (
      {stage0_34[448]},
      {stage1_34[204]}
   );
   gpc1_1 gpc4085 (
      {stage0_34[449]},
      {stage1_34[205]}
   );
   gpc1_1 gpc4086 (
      {stage0_34[450]},
      {stage1_34[206]}
   );
   gpc1_1 gpc4087 (
      {stage0_34[451]},
      {stage1_34[207]}
   );
   gpc1_1 gpc4088 (
      {stage0_34[452]},
      {stage1_34[208]}
   );
   gpc1_1 gpc4089 (
      {stage0_34[453]},
      {stage1_34[209]}
   );
   gpc1_1 gpc4090 (
      {stage0_34[454]},
      {stage1_34[210]}
   );
   gpc1_1 gpc4091 (
      {stage0_34[455]},
      {stage1_34[211]}
   );
   gpc1_1 gpc4092 (
      {stage0_34[456]},
      {stage1_34[212]}
   );
   gpc1_1 gpc4093 (
      {stage0_34[457]},
      {stage1_34[213]}
   );
   gpc1_1 gpc4094 (
      {stage0_34[458]},
      {stage1_34[214]}
   );
   gpc1_1 gpc4095 (
      {stage0_34[459]},
      {stage1_34[215]}
   );
   gpc1_1 gpc4096 (
      {stage0_34[460]},
      {stage1_34[216]}
   );
   gpc1_1 gpc4097 (
      {stage0_34[461]},
      {stage1_34[217]}
   );
   gpc1_1 gpc4098 (
      {stage0_34[462]},
      {stage1_34[218]}
   );
   gpc1_1 gpc4099 (
      {stage0_34[463]},
      {stage1_34[219]}
   );
   gpc1_1 gpc4100 (
      {stage0_34[464]},
      {stage1_34[220]}
   );
   gpc1_1 gpc4101 (
      {stage0_34[465]},
      {stage1_34[221]}
   );
   gpc1_1 gpc4102 (
      {stage0_34[466]},
      {stage1_34[222]}
   );
   gpc1_1 gpc4103 (
      {stage0_34[467]},
      {stage1_34[223]}
   );
   gpc1_1 gpc4104 (
      {stage0_34[468]},
      {stage1_34[224]}
   );
   gpc1_1 gpc4105 (
      {stage0_34[469]},
      {stage1_34[225]}
   );
   gpc1_1 gpc4106 (
      {stage0_34[470]},
      {stage1_34[226]}
   );
   gpc1_1 gpc4107 (
      {stage0_34[471]},
      {stage1_34[227]}
   );
   gpc1_1 gpc4108 (
      {stage0_34[472]},
      {stage1_34[228]}
   );
   gpc1_1 gpc4109 (
      {stage0_34[473]},
      {stage1_34[229]}
   );
   gpc1_1 gpc4110 (
      {stage0_34[474]},
      {stage1_34[230]}
   );
   gpc1_1 gpc4111 (
      {stage0_34[475]},
      {stage1_34[231]}
   );
   gpc1_1 gpc4112 (
      {stage0_34[476]},
      {stage1_34[232]}
   );
   gpc1_1 gpc4113 (
      {stage0_34[477]},
      {stage1_34[233]}
   );
   gpc1_1 gpc4114 (
      {stage0_34[478]},
      {stage1_34[234]}
   );
   gpc1_1 gpc4115 (
      {stage0_34[479]},
      {stage1_34[235]}
   );
   gpc1_1 gpc4116 (
      {stage0_34[480]},
      {stage1_34[236]}
   );
   gpc1_1 gpc4117 (
      {stage0_34[481]},
      {stage1_34[237]}
   );
   gpc1_1 gpc4118 (
      {stage0_34[482]},
      {stage1_34[238]}
   );
   gpc1_1 gpc4119 (
      {stage0_34[483]},
      {stage1_34[239]}
   );
   gpc1_1 gpc4120 (
      {stage0_34[484]},
      {stage1_34[240]}
   );
   gpc1_1 gpc4121 (
      {stage0_34[485]},
      {stage1_34[241]}
   );
   gpc1_1 gpc4122 (
      {stage0_34[486]},
      {stage1_34[242]}
   );
   gpc1_1 gpc4123 (
      {stage0_34[487]},
      {stage1_34[243]}
   );
   gpc1_1 gpc4124 (
      {stage0_34[488]},
      {stage1_34[244]}
   );
   gpc1_1 gpc4125 (
      {stage0_34[489]},
      {stage1_34[245]}
   );
   gpc1_1 gpc4126 (
      {stage0_34[490]},
      {stage1_34[246]}
   );
   gpc1_1 gpc4127 (
      {stage0_34[491]},
      {stage1_34[247]}
   );
   gpc1_1 gpc4128 (
      {stage0_34[492]},
      {stage1_34[248]}
   );
   gpc1_1 gpc4129 (
      {stage0_34[493]},
      {stage1_34[249]}
   );
   gpc1_1 gpc4130 (
      {stage0_34[494]},
      {stage1_34[250]}
   );
   gpc1_1 gpc4131 (
      {stage0_34[495]},
      {stage1_34[251]}
   );
   gpc1_1 gpc4132 (
      {stage0_34[496]},
      {stage1_34[252]}
   );
   gpc1_1 gpc4133 (
      {stage0_34[497]},
      {stage1_34[253]}
   );
   gpc1_1 gpc4134 (
      {stage0_34[498]},
      {stage1_34[254]}
   );
   gpc1_1 gpc4135 (
      {stage0_34[499]},
      {stage1_34[255]}
   );
   gpc1_1 gpc4136 (
      {stage0_34[500]},
      {stage1_34[256]}
   );
   gpc1_1 gpc4137 (
      {stage0_34[501]},
      {stage1_34[257]}
   );
   gpc1_1 gpc4138 (
      {stage0_34[502]},
      {stage1_34[258]}
   );
   gpc1_1 gpc4139 (
      {stage0_34[503]},
      {stage1_34[259]}
   );
   gpc1_1 gpc4140 (
      {stage0_34[504]},
      {stage1_34[260]}
   );
   gpc1_1 gpc4141 (
      {stage0_34[505]},
      {stage1_34[261]}
   );
   gpc1_1 gpc4142 (
      {stage0_34[506]},
      {stage1_34[262]}
   );
   gpc1_1 gpc4143 (
      {stage0_34[507]},
      {stage1_34[263]}
   );
   gpc1_1 gpc4144 (
      {stage0_34[508]},
      {stage1_34[264]}
   );
   gpc1_1 gpc4145 (
      {stage0_34[509]},
      {stage1_34[265]}
   );
   gpc1_1 gpc4146 (
      {stage0_34[510]},
      {stage1_34[266]}
   );
   gpc1_1 gpc4147 (
      {stage0_34[511]},
      {stage1_34[267]}
   );
   gpc1_1 gpc4148 (
      {stage0_35[495]},
      {stage1_35[174]}
   );
   gpc1_1 gpc4149 (
      {stage0_35[496]},
      {stage1_35[175]}
   );
   gpc1_1 gpc4150 (
      {stage0_35[497]},
      {stage1_35[176]}
   );
   gpc1_1 gpc4151 (
      {stage0_35[498]},
      {stage1_35[177]}
   );
   gpc1_1 gpc4152 (
      {stage0_35[499]},
      {stage1_35[178]}
   );
   gpc1_1 gpc4153 (
      {stage0_35[500]},
      {stage1_35[179]}
   );
   gpc1_1 gpc4154 (
      {stage0_35[501]},
      {stage1_35[180]}
   );
   gpc1_1 gpc4155 (
      {stage0_35[502]},
      {stage1_35[181]}
   );
   gpc1_1 gpc4156 (
      {stage0_35[503]},
      {stage1_35[182]}
   );
   gpc1_1 gpc4157 (
      {stage0_35[504]},
      {stage1_35[183]}
   );
   gpc1_1 gpc4158 (
      {stage0_35[505]},
      {stage1_35[184]}
   );
   gpc1_1 gpc4159 (
      {stage0_35[506]},
      {stage1_35[185]}
   );
   gpc1_1 gpc4160 (
      {stage0_35[507]},
      {stage1_35[186]}
   );
   gpc1_1 gpc4161 (
      {stage0_35[508]},
      {stage1_35[187]}
   );
   gpc1_1 gpc4162 (
      {stage0_35[509]},
      {stage1_35[188]}
   );
   gpc1_1 gpc4163 (
      {stage0_35[510]},
      {stage1_35[189]}
   );
   gpc1_1 gpc4164 (
      {stage0_35[511]},
      {stage1_35[190]}
   );
   gpc1_1 gpc4165 (
      {stage0_36[367]},
      {stage1_36[186]}
   );
   gpc1_1 gpc4166 (
      {stage0_36[368]},
      {stage1_36[187]}
   );
   gpc1_1 gpc4167 (
      {stage0_36[369]},
      {stage1_36[188]}
   );
   gpc1_1 gpc4168 (
      {stage0_36[370]},
      {stage1_36[189]}
   );
   gpc1_1 gpc4169 (
      {stage0_36[371]},
      {stage1_36[190]}
   );
   gpc1_1 gpc4170 (
      {stage0_36[372]},
      {stage1_36[191]}
   );
   gpc1_1 gpc4171 (
      {stage0_36[373]},
      {stage1_36[192]}
   );
   gpc1_1 gpc4172 (
      {stage0_36[374]},
      {stage1_36[193]}
   );
   gpc1_1 gpc4173 (
      {stage0_36[375]},
      {stage1_36[194]}
   );
   gpc1_1 gpc4174 (
      {stage0_36[376]},
      {stage1_36[195]}
   );
   gpc1_1 gpc4175 (
      {stage0_36[377]},
      {stage1_36[196]}
   );
   gpc1_1 gpc4176 (
      {stage0_36[378]},
      {stage1_36[197]}
   );
   gpc1_1 gpc4177 (
      {stage0_36[379]},
      {stage1_36[198]}
   );
   gpc1_1 gpc4178 (
      {stage0_36[380]},
      {stage1_36[199]}
   );
   gpc1_1 gpc4179 (
      {stage0_36[381]},
      {stage1_36[200]}
   );
   gpc1_1 gpc4180 (
      {stage0_36[382]},
      {stage1_36[201]}
   );
   gpc1_1 gpc4181 (
      {stage0_36[383]},
      {stage1_36[202]}
   );
   gpc1_1 gpc4182 (
      {stage0_36[384]},
      {stage1_36[203]}
   );
   gpc1_1 gpc4183 (
      {stage0_36[385]},
      {stage1_36[204]}
   );
   gpc1_1 gpc4184 (
      {stage0_36[386]},
      {stage1_36[205]}
   );
   gpc1_1 gpc4185 (
      {stage0_36[387]},
      {stage1_36[206]}
   );
   gpc1_1 gpc4186 (
      {stage0_36[388]},
      {stage1_36[207]}
   );
   gpc1_1 gpc4187 (
      {stage0_36[389]},
      {stage1_36[208]}
   );
   gpc1_1 gpc4188 (
      {stage0_36[390]},
      {stage1_36[209]}
   );
   gpc1_1 gpc4189 (
      {stage0_36[391]},
      {stage1_36[210]}
   );
   gpc1_1 gpc4190 (
      {stage0_36[392]},
      {stage1_36[211]}
   );
   gpc1_1 gpc4191 (
      {stage0_36[393]},
      {stage1_36[212]}
   );
   gpc1_1 gpc4192 (
      {stage0_36[394]},
      {stage1_36[213]}
   );
   gpc1_1 gpc4193 (
      {stage0_36[395]},
      {stage1_36[214]}
   );
   gpc1_1 gpc4194 (
      {stage0_36[396]},
      {stage1_36[215]}
   );
   gpc1_1 gpc4195 (
      {stage0_36[397]},
      {stage1_36[216]}
   );
   gpc1_1 gpc4196 (
      {stage0_36[398]},
      {stage1_36[217]}
   );
   gpc1_1 gpc4197 (
      {stage0_36[399]},
      {stage1_36[218]}
   );
   gpc1_1 gpc4198 (
      {stage0_36[400]},
      {stage1_36[219]}
   );
   gpc1_1 gpc4199 (
      {stage0_36[401]},
      {stage1_36[220]}
   );
   gpc1_1 gpc4200 (
      {stage0_36[402]},
      {stage1_36[221]}
   );
   gpc1_1 gpc4201 (
      {stage0_36[403]},
      {stage1_36[222]}
   );
   gpc1_1 gpc4202 (
      {stage0_36[404]},
      {stage1_36[223]}
   );
   gpc1_1 gpc4203 (
      {stage0_36[405]},
      {stage1_36[224]}
   );
   gpc1_1 gpc4204 (
      {stage0_36[406]},
      {stage1_36[225]}
   );
   gpc1_1 gpc4205 (
      {stage0_36[407]},
      {stage1_36[226]}
   );
   gpc1_1 gpc4206 (
      {stage0_36[408]},
      {stage1_36[227]}
   );
   gpc1_1 gpc4207 (
      {stage0_36[409]},
      {stage1_36[228]}
   );
   gpc1_1 gpc4208 (
      {stage0_36[410]},
      {stage1_36[229]}
   );
   gpc1_1 gpc4209 (
      {stage0_36[411]},
      {stage1_36[230]}
   );
   gpc1_1 gpc4210 (
      {stage0_36[412]},
      {stage1_36[231]}
   );
   gpc1_1 gpc4211 (
      {stage0_36[413]},
      {stage1_36[232]}
   );
   gpc1_1 gpc4212 (
      {stage0_36[414]},
      {stage1_36[233]}
   );
   gpc1_1 gpc4213 (
      {stage0_36[415]},
      {stage1_36[234]}
   );
   gpc1_1 gpc4214 (
      {stage0_36[416]},
      {stage1_36[235]}
   );
   gpc1_1 gpc4215 (
      {stage0_36[417]},
      {stage1_36[236]}
   );
   gpc1_1 gpc4216 (
      {stage0_36[418]},
      {stage1_36[237]}
   );
   gpc1_1 gpc4217 (
      {stage0_36[419]},
      {stage1_36[238]}
   );
   gpc1_1 gpc4218 (
      {stage0_36[420]},
      {stage1_36[239]}
   );
   gpc1_1 gpc4219 (
      {stage0_36[421]},
      {stage1_36[240]}
   );
   gpc1_1 gpc4220 (
      {stage0_36[422]},
      {stage1_36[241]}
   );
   gpc1_1 gpc4221 (
      {stage0_36[423]},
      {stage1_36[242]}
   );
   gpc1_1 gpc4222 (
      {stage0_36[424]},
      {stage1_36[243]}
   );
   gpc1_1 gpc4223 (
      {stage0_36[425]},
      {stage1_36[244]}
   );
   gpc1_1 gpc4224 (
      {stage0_36[426]},
      {stage1_36[245]}
   );
   gpc1_1 gpc4225 (
      {stage0_36[427]},
      {stage1_36[246]}
   );
   gpc1_1 gpc4226 (
      {stage0_36[428]},
      {stage1_36[247]}
   );
   gpc1_1 gpc4227 (
      {stage0_36[429]},
      {stage1_36[248]}
   );
   gpc1_1 gpc4228 (
      {stage0_36[430]},
      {stage1_36[249]}
   );
   gpc1_1 gpc4229 (
      {stage0_36[431]},
      {stage1_36[250]}
   );
   gpc1_1 gpc4230 (
      {stage0_36[432]},
      {stage1_36[251]}
   );
   gpc1_1 gpc4231 (
      {stage0_36[433]},
      {stage1_36[252]}
   );
   gpc1_1 gpc4232 (
      {stage0_36[434]},
      {stage1_36[253]}
   );
   gpc1_1 gpc4233 (
      {stage0_36[435]},
      {stage1_36[254]}
   );
   gpc1_1 gpc4234 (
      {stage0_36[436]},
      {stage1_36[255]}
   );
   gpc1_1 gpc4235 (
      {stage0_36[437]},
      {stage1_36[256]}
   );
   gpc1_1 gpc4236 (
      {stage0_36[438]},
      {stage1_36[257]}
   );
   gpc1_1 gpc4237 (
      {stage0_36[439]},
      {stage1_36[258]}
   );
   gpc1_1 gpc4238 (
      {stage0_36[440]},
      {stage1_36[259]}
   );
   gpc1_1 gpc4239 (
      {stage0_36[441]},
      {stage1_36[260]}
   );
   gpc1_1 gpc4240 (
      {stage0_36[442]},
      {stage1_36[261]}
   );
   gpc1_1 gpc4241 (
      {stage0_36[443]},
      {stage1_36[262]}
   );
   gpc1_1 gpc4242 (
      {stage0_36[444]},
      {stage1_36[263]}
   );
   gpc1_1 gpc4243 (
      {stage0_36[445]},
      {stage1_36[264]}
   );
   gpc1_1 gpc4244 (
      {stage0_36[446]},
      {stage1_36[265]}
   );
   gpc1_1 gpc4245 (
      {stage0_36[447]},
      {stage1_36[266]}
   );
   gpc1_1 gpc4246 (
      {stage0_36[448]},
      {stage1_36[267]}
   );
   gpc1_1 gpc4247 (
      {stage0_36[449]},
      {stage1_36[268]}
   );
   gpc1_1 gpc4248 (
      {stage0_36[450]},
      {stage1_36[269]}
   );
   gpc1_1 gpc4249 (
      {stage0_36[451]},
      {stage1_36[270]}
   );
   gpc1_1 gpc4250 (
      {stage0_36[452]},
      {stage1_36[271]}
   );
   gpc1_1 gpc4251 (
      {stage0_36[453]},
      {stage1_36[272]}
   );
   gpc1_1 gpc4252 (
      {stage0_36[454]},
      {stage1_36[273]}
   );
   gpc1_1 gpc4253 (
      {stage0_36[455]},
      {stage1_36[274]}
   );
   gpc1_1 gpc4254 (
      {stage0_36[456]},
      {stage1_36[275]}
   );
   gpc1_1 gpc4255 (
      {stage0_36[457]},
      {stage1_36[276]}
   );
   gpc1_1 gpc4256 (
      {stage0_36[458]},
      {stage1_36[277]}
   );
   gpc1_1 gpc4257 (
      {stage0_36[459]},
      {stage1_36[278]}
   );
   gpc1_1 gpc4258 (
      {stage0_36[460]},
      {stage1_36[279]}
   );
   gpc1_1 gpc4259 (
      {stage0_36[461]},
      {stage1_36[280]}
   );
   gpc1_1 gpc4260 (
      {stage0_36[462]},
      {stage1_36[281]}
   );
   gpc1_1 gpc4261 (
      {stage0_36[463]},
      {stage1_36[282]}
   );
   gpc1_1 gpc4262 (
      {stage0_36[464]},
      {stage1_36[283]}
   );
   gpc1_1 gpc4263 (
      {stage0_36[465]},
      {stage1_36[284]}
   );
   gpc1_1 gpc4264 (
      {stage0_36[466]},
      {stage1_36[285]}
   );
   gpc1_1 gpc4265 (
      {stage0_36[467]},
      {stage1_36[286]}
   );
   gpc1_1 gpc4266 (
      {stage0_36[468]},
      {stage1_36[287]}
   );
   gpc1_1 gpc4267 (
      {stage0_36[469]},
      {stage1_36[288]}
   );
   gpc1_1 gpc4268 (
      {stage0_36[470]},
      {stage1_36[289]}
   );
   gpc1_1 gpc4269 (
      {stage0_36[471]},
      {stage1_36[290]}
   );
   gpc1_1 gpc4270 (
      {stage0_36[472]},
      {stage1_36[291]}
   );
   gpc1_1 gpc4271 (
      {stage0_36[473]},
      {stage1_36[292]}
   );
   gpc1_1 gpc4272 (
      {stage0_36[474]},
      {stage1_36[293]}
   );
   gpc1_1 gpc4273 (
      {stage0_36[475]},
      {stage1_36[294]}
   );
   gpc1_1 gpc4274 (
      {stage0_36[476]},
      {stage1_36[295]}
   );
   gpc1_1 gpc4275 (
      {stage0_36[477]},
      {stage1_36[296]}
   );
   gpc1_1 gpc4276 (
      {stage0_36[478]},
      {stage1_36[297]}
   );
   gpc1_1 gpc4277 (
      {stage0_36[479]},
      {stage1_36[298]}
   );
   gpc1_1 gpc4278 (
      {stage0_36[480]},
      {stage1_36[299]}
   );
   gpc1_1 gpc4279 (
      {stage0_36[481]},
      {stage1_36[300]}
   );
   gpc1_1 gpc4280 (
      {stage0_36[482]},
      {stage1_36[301]}
   );
   gpc1_1 gpc4281 (
      {stage0_36[483]},
      {stage1_36[302]}
   );
   gpc1_1 gpc4282 (
      {stage0_36[484]},
      {stage1_36[303]}
   );
   gpc1_1 gpc4283 (
      {stage0_36[485]},
      {stage1_36[304]}
   );
   gpc1_1 gpc4284 (
      {stage0_36[486]},
      {stage1_36[305]}
   );
   gpc1_1 gpc4285 (
      {stage0_36[487]},
      {stage1_36[306]}
   );
   gpc1_1 gpc4286 (
      {stage0_36[488]},
      {stage1_36[307]}
   );
   gpc1_1 gpc4287 (
      {stage0_36[489]},
      {stage1_36[308]}
   );
   gpc1_1 gpc4288 (
      {stage0_36[490]},
      {stage1_36[309]}
   );
   gpc1_1 gpc4289 (
      {stage0_36[491]},
      {stage1_36[310]}
   );
   gpc1_1 gpc4290 (
      {stage0_36[492]},
      {stage1_36[311]}
   );
   gpc1_1 gpc4291 (
      {stage0_36[493]},
      {stage1_36[312]}
   );
   gpc1_1 gpc4292 (
      {stage0_36[494]},
      {stage1_36[313]}
   );
   gpc1_1 gpc4293 (
      {stage0_36[495]},
      {stage1_36[314]}
   );
   gpc1_1 gpc4294 (
      {stage0_36[496]},
      {stage1_36[315]}
   );
   gpc1_1 gpc4295 (
      {stage0_36[497]},
      {stage1_36[316]}
   );
   gpc1_1 gpc4296 (
      {stage0_36[498]},
      {stage1_36[317]}
   );
   gpc1_1 gpc4297 (
      {stage0_36[499]},
      {stage1_36[318]}
   );
   gpc1_1 gpc4298 (
      {stage0_36[500]},
      {stage1_36[319]}
   );
   gpc1_1 gpc4299 (
      {stage0_36[501]},
      {stage1_36[320]}
   );
   gpc1_1 gpc4300 (
      {stage0_36[502]},
      {stage1_36[321]}
   );
   gpc1_1 gpc4301 (
      {stage0_36[503]},
      {stage1_36[322]}
   );
   gpc1_1 gpc4302 (
      {stage0_36[504]},
      {stage1_36[323]}
   );
   gpc1_1 gpc4303 (
      {stage0_36[505]},
      {stage1_36[324]}
   );
   gpc1_1 gpc4304 (
      {stage0_36[506]},
      {stage1_36[325]}
   );
   gpc1_1 gpc4305 (
      {stage0_36[507]},
      {stage1_36[326]}
   );
   gpc1_1 gpc4306 (
      {stage0_36[508]},
      {stage1_36[327]}
   );
   gpc1_1 gpc4307 (
      {stage0_36[509]},
      {stage1_36[328]}
   );
   gpc1_1 gpc4308 (
      {stage0_36[510]},
      {stage1_36[329]}
   );
   gpc1_1 gpc4309 (
      {stage0_36[511]},
      {stage1_36[330]}
   );
   gpc1_1 gpc4310 (
      {stage0_37[392]},
      {stage1_37[183]}
   );
   gpc1_1 gpc4311 (
      {stage0_37[393]},
      {stage1_37[184]}
   );
   gpc1_1 gpc4312 (
      {stage0_37[394]},
      {stage1_37[185]}
   );
   gpc1_1 gpc4313 (
      {stage0_37[395]},
      {stage1_37[186]}
   );
   gpc1_1 gpc4314 (
      {stage0_37[396]},
      {stage1_37[187]}
   );
   gpc1_1 gpc4315 (
      {stage0_37[397]},
      {stage1_37[188]}
   );
   gpc1_1 gpc4316 (
      {stage0_37[398]},
      {stage1_37[189]}
   );
   gpc1_1 gpc4317 (
      {stage0_37[399]},
      {stage1_37[190]}
   );
   gpc1_1 gpc4318 (
      {stage0_37[400]},
      {stage1_37[191]}
   );
   gpc1_1 gpc4319 (
      {stage0_37[401]},
      {stage1_37[192]}
   );
   gpc1_1 gpc4320 (
      {stage0_37[402]},
      {stage1_37[193]}
   );
   gpc1_1 gpc4321 (
      {stage0_37[403]},
      {stage1_37[194]}
   );
   gpc1_1 gpc4322 (
      {stage0_37[404]},
      {stage1_37[195]}
   );
   gpc1_1 gpc4323 (
      {stage0_37[405]},
      {stage1_37[196]}
   );
   gpc1_1 gpc4324 (
      {stage0_37[406]},
      {stage1_37[197]}
   );
   gpc1_1 gpc4325 (
      {stage0_37[407]},
      {stage1_37[198]}
   );
   gpc1_1 gpc4326 (
      {stage0_37[408]},
      {stage1_37[199]}
   );
   gpc1_1 gpc4327 (
      {stage0_37[409]},
      {stage1_37[200]}
   );
   gpc1_1 gpc4328 (
      {stage0_37[410]},
      {stage1_37[201]}
   );
   gpc1_1 gpc4329 (
      {stage0_37[411]},
      {stage1_37[202]}
   );
   gpc1_1 gpc4330 (
      {stage0_37[412]},
      {stage1_37[203]}
   );
   gpc1_1 gpc4331 (
      {stage0_37[413]},
      {stage1_37[204]}
   );
   gpc1_1 gpc4332 (
      {stage0_37[414]},
      {stage1_37[205]}
   );
   gpc1_1 gpc4333 (
      {stage0_37[415]},
      {stage1_37[206]}
   );
   gpc1_1 gpc4334 (
      {stage0_37[416]},
      {stage1_37[207]}
   );
   gpc1_1 gpc4335 (
      {stage0_37[417]},
      {stage1_37[208]}
   );
   gpc1_1 gpc4336 (
      {stage0_37[418]},
      {stage1_37[209]}
   );
   gpc1_1 gpc4337 (
      {stage0_37[419]},
      {stage1_37[210]}
   );
   gpc1_1 gpc4338 (
      {stage0_37[420]},
      {stage1_37[211]}
   );
   gpc1_1 gpc4339 (
      {stage0_37[421]},
      {stage1_37[212]}
   );
   gpc1_1 gpc4340 (
      {stage0_37[422]},
      {stage1_37[213]}
   );
   gpc1_1 gpc4341 (
      {stage0_37[423]},
      {stage1_37[214]}
   );
   gpc1_1 gpc4342 (
      {stage0_37[424]},
      {stage1_37[215]}
   );
   gpc1_1 gpc4343 (
      {stage0_37[425]},
      {stage1_37[216]}
   );
   gpc1_1 gpc4344 (
      {stage0_37[426]},
      {stage1_37[217]}
   );
   gpc1_1 gpc4345 (
      {stage0_37[427]},
      {stage1_37[218]}
   );
   gpc1_1 gpc4346 (
      {stage0_37[428]},
      {stage1_37[219]}
   );
   gpc1_1 gpc4347 (
      {stage0_37[429]},
      {stage1_37[220]}
   );
   gpc1_1 gpc4348 (
      {stage0_37[430]},
      {stage1_37[221]}
   );
   gpc1_1 gpc4349 (
      {stage0_37[431]},
      {stage1_37[222]}
   );
   gpc1_1 gpc4350 (
      {stage0_37[432]},
      {stage1_37[223]}
   );
   gpc1_1 gpc4351 (
      {stage0_37[433]},
      {stage1_37[224]}
   );
   gpc1_1 gpc4352 (
      {stage0_37[434]},
      {stage1_37[225]}
   );
   gpc1_1 gpc4353 (
      {stage0_37[435]},
      {stage1_37[226]}
   );
   gpc1_1 gpc4354 (
      {stage0_37[436]},
      {stage1_37[227]}
   );
   gpc1_1 gpc4355 (
      {stage0_37[437]},
      {stage1_37[228]}
   );
   gpc1_1 gpc4356 (
      {stage0_37[438]},
      {stage1_37[229]}
   );
   gpc1_1 gpc4357 (
      {stage0_37[439]},
      {stage1_37[230]}
   );
   gpc1_1 gpc4358 (
      {stage0_37[440]},
      {stage1_37[231]}
   );
   gpc1_1 gpc4359 (
      {stage0_37[441]},
      {stage1_37[232]}
   );
   gpc1_1 gpc4360 (
      {stage0_37[442]},
      {stage1_37[233]}
   );
   gpc1_1 gpc4361 (
      {stage0_37[443]},
      {stage1_37[234]}
   );
   gpc1_1 gpc4362 (
      {stage0_37[444]},
      {stage1_37[235]}
   );
   gpc1_1 gpc4363 (
      {stage0_37[445]},
      {stage1_37[236]}
   );
   gpc1_1 gpc4364 (
      {stage0_37[446]},
      {stage1_37[237]}
   );
   gpc1_1 gpc4365 (
      {stage0_37[447]},
      {stage1_37[238]}
   );
   gpc1_1 gpc4366 (
      {stage0_37[448]},
      {stage1_37[239]}
   );
   gpc1_1 gpc4367 (
      {stage0_37[449]},
      {stage1_37[240]}
   );
   gpc1_1 gpc4368 (
      {stage0_37[450]},
      {stage1_37[241]}
   );
   gpc1_1 gpc4369 (
      {stage0_37[451]},
      {stage1_37[242]}
   );
   gpc1_1 gpc4370 (
      {stage0_37[452]},
      {stage1_37[243]}
   );
   gpc1_1 gpc4371 (
      {stage0_37[453]},
      {stage1_37[244]}
   );
   gpc1_1 gpc4372 (
      {stage0_37[454]},
      {stage1_37[245]}
   );
   gpc1_1 gpc4373 (
      {stage0_37[455]},
      {stage1_37[246]}
   );
   gpc1_1 gpc4374 (
      {stage0_37[456]},
      {stage1_37[247]}
   );
   gpc1_1 gpc4375 (
      {stage0_37[457]},
      {stage1_37[248]}
   );
   gpc1_1 gpc4376 (
      {stage0_37[458]},
      {stage1_37[249]}
   );
   gpc1_1 gpc4377 (
      {stage0_37[459]},
      {stage1_37[250]}
   );
   gpc1_1 gpc4378 (
      {stage0_37[460]},
      {stage1_37[251]}
   );
   gpc1_1 gpc4379 (
      {stage0_37[461]},
      {stage1_37[252]}
   );
   gpc1_1 gpc4380 (
      {stage0_37[462]},
      {stage1_37[253]}
   );
   gpc1_1 gpc4381 (
      {stage0_37[463]},
      {stage1_37[254]}
   );
   gpc1_1 gpc4382 (
      {stage0_37[464]},
      {stage1_37[255]}
   );
   gpc1_1 gpc4383 (
      {stage0_37[465]},
      {stage1_37[256]}
   );
   gpc1_1 gpc4384 (
      {stage0_37[466]},
      {stage1_37[257]}
   );
   gpc1_1 gpc4385 (
      {stage0_37[467]},
      {stage1_37[258]}
   );
   gpc1_1 gpc4386 (
      {stage0_37[468]},
      {stage1_37[259]}
   );
   gpc1_1 gpc4387 (
      {stage0_37[469]},
      {stage1_37[260]}
   );
   gpc1_1 gpc4388 (
      {stage0_37[470]},
      {stage1_37[261]}
   );
   gpc1_1 gpc4389 (
      {stage0_37[471]},
      {stage1_37[262]}
   );
   gpc1_1 gpc4390 (
      {stage0_37[472]},
      {stage1_37[263]}
   );
   gpc1_1 gpc4391 (
      {stage0_37[473]},
      {stage1_37[264]}
   );
   gpc1_1 gpc4392 (
      {stage0_37[474]},
      {stage1_37[265]}
   );
   gpc1_1 gpc4393 (
      {stage0_37[475]},
      {stage1_37[266]}
   );
   gpc1_1 gpc4394 (
      {stage0_37[476]},
      {stage1_37[267]}
   );
   gpc1_1 gpc4395 (
      {stage0_37[477]},
      {stage1_37[268]}
   );
   gpc1_1 gpc4396 (
      {stage0_37[478]},
      {stage1_37[269]}
   );
   gpc1_1 gpc4397 (
      {stage0_37[479]},
      {stage1_37[270]}
   );
   gpc1_1 gpc4398 (
      {stage0_37[480]},
      {stage1_37[271]}
   );
   gpc1_1 gpc4399 (
      {stage0_37[481]},
      {stage1_37[272]}
   );
   gpc1_1 gpc4400 (
      {stage0_37[482]},
      {stage1_37[273]}
   );
   gpc1_1 gpc4401 (
      {stage0_37[483]},
      {stage1_37[274]}
   );
   gpc1_1 gpc4402 (
      {stage0_37[484]},
      {stage1_37[275]}
   );
   gpc1_1 gpc4403 (
      {stage0_37[485]},
      {stage1_37[276]}
   );
   gpc1_1 gpc4404 (
      {stage0_37[486]},
      {stage1_37[277]}
   );
   gpc1_1 gpc4405 (
      {stage0_37[487]},
      {stage1_37[278]}
   );
   gpc1_1 gpc4406 (
      {stage0_37[488]},
      {stage1_37[279]}
   );
   gpc1_1 gpc4407 (
      {stage0_37[489]},
      {stage1_37[280]}
   );
   gpc1_1 gpc4408 (
      {stage0_37[490]},
      {stage1_37[281]}
   );
   gpc1_1 gpc4409 (
      {stage0_37[491]},
      {stage1_37[282]}
   );
   gpc1_1 gpc4410 (
      {stage0_37[492]},
      {stage1_37[283]}
   );
   gpc1_1 gpc4411 (
      {stage0_37[493]},
      {stage1_37[284]}
   );
   gpc1_1 gpc4412 (
      {stage0_37[494]},
      {stage1_37[285]}
   );
   gpc1_1 gpc4413 (
      {stage0_37[495]},
      {stage1_37[286]}
   );
   gpc1_1 gpc4414 (
      {stage0_37[496]},
      {stage1_37[287]}
   );
   gpc1_1 gpc4415 (
      {stage0_37[497]},
      {stage1_37[288]}
   );
   gpc1_1 gpc4416 (
      {stage0_37[498]},
      {stage1_37[289]}
   );
   gpc1_1 gpc4417 (
      {stage0_37[499]},
      {stage1_37[290]}
   );
   gpc1_1 gpc4418 (
      {stage0_37[500]},
      {stage1_37[291]}
   );
   gpc1_1 gpc4419 (
      {stage0_37[501]},
      {stage1_37[292]}
   );
   gpc1_1 gpc4420 (
      {stage0_37[502]},
      {stage1_37[293]}
   );
   gpc1_1 gpc4421 (
      {stage0_37[503]},
      {stage1_37[294]}
   );
   gpc1_1 gpc4422 (
      {stage0_37[504]},
      {stage1_37[295]}
   );
   gpc1_1 gpc4423 (
      {stage0_37[505]},
      {stage1_37[296]}
   );
   gpc1_1 gpc4424 (
      {stage0_37[506]},
      {stage1_37[297]}
   );
   gpc1_1 gpc4425 (
      {stage0_37[507]},
      {stage1_37[298]}
   );
   gpc1_1 gpc4426 (
      {stage0_37[508]},
      {stage1_37[299]}
   );
   gpc1_1 gpc4427 (
      {stage0_37[509]},
      {stage1_37[300]}
   );
   gpc1_1 gpc4428 (
      {stage0_37[510]},
      {stage1_37[301]}
   );
   gpc1_1 gpc4429 (
      {stage0_37[511]},
      {stage1_37[302]}
   );
   gpc1_1 gpc4430 (
      {stage0_38[382]},
      {stage1_38[147]}
   );
   gpc1_1 gpc4431 (
      {stage0_38[383]},
      {stage1_38[148]}
   );
   gpc1_1 gpc4432 (
      {stage0_38[384]},
      {stage1_38[149]}
   );
   gpc1_1 gpc4433 (
      {stage0_38[385]},
      {stage1_38[150]}
   );
   gpc1_1 gpc4434 (
      {stage0_38[386]},
      {stage1_38[151]}
   );
   gpc1_1 gpc4435 (
      {stage0_38[387]},
      {stage1_38[152]}
   );
   gpc1_1 gpc4436 (
      {stage0_38[388]},
      {stage1_38[153]}
   );
   gpc1_1 gpc4437 (
      {stage0_38[389]},
      {stage1_38[154]}
   );
   gpc1_1 gpc4438 (
      {stage0_38[390]},
      {stage1_38[155]}
   );
   gpc1_1 gpc4439 (
      {stage0_38[391]},
      {stage1_38[156]}
   );
   gpc1_1 gpc4440 (
      {stage0_38[392]},
      {stage1_38[157]}
   );
   gpc1_1 gpc4441 (
      {stage0_38[393]},
      {stage1_38[158]}
   );
   gpc1_1 gpc4442 (
      {stage0_38[394]},
      {stage1_38[159]}
   );
   gpc1_1 gpc4443 (
      {stage0_38[395]},
      {stage1_38[160]}
   );
   gpc1_1 gpc4444 (
      {stage0_38[396]},
      {stage1_38[161]}
   );
   gpc1_1 gpc4445 (
      {stage0_38[397]},
      {stage1_38[162]}
   );
   gpc1_1 gpc4446 (
      {stage0_38[398]},
      {stage1_38[163]}
   );
   gpc1_1 gpc4447 (
      {stage0_38[399]},
      {stage1_38[164]}
   );
   gpc1_1 gpc4448 (
      {stage0_38[400]},
      {stage1_38[165]}
   );
   gpc1_1 gpc4449 (
      {stage0_38[401]},
      {stage1_38[166]}
   );
   gpc1_1 gpc4450 (
      {stage0_38[402]},
      {stage1_38[167]}
   );
   gpc1_1 gpc4451 (
      {stage0_38[403]},
      {stage1_38[168]}
   );
   gpc1_1 gpc4452 (
      {stage0_38[404]},
      {stage1_38[169]}
   );
   gpc1_1 gpc4453 (
      {stage0_38[405]},
      {stage1_38[170]}
   );
   gpc1_1 gpc4454 (
      {stage0_38[406]},
      {stage1_38[171]}
   );
   gpc1_1 gpc4455 (
      {stage0_38[407]},
      {stage1_38[172]}
   );
   gpc1_1 gpc4456 (
      {stage0_38[408]},
      {stage1_38[173]}
   );
   gpc1_1 gpc4457 (
      {stage0_38[409]},
      {stage1_38[174]}
   );
   gpc1_1 gpc4458 (
      {stage0_38[410]},
      {stage1_38[175]}
   );
   gpc1_1 gpc4459 (
      {stage0_38[411]},
      {stage1_38[176]}
   );
   gpc1_1 gpc4460 (
      {stage0_38[412]},
      {stage1_38[177]}
   );
   gpc1_1 gpc4461 (
      {stage0_38[413]},
      {stage1_38[178]}
   );
   gpc1_1 gpc4462 (
      {stage0_38[414]},
      {stage1_38[179]}
   );
   gpc1_1 gpc4463 (
      {stage0_38[415]},
      {stage1_38[180]}
   );
   gpc1_1 gpc4464 (
      {stage0_38[416]},
      {stage1_38[181]}
   );
   gpc1_1 gpc4465 (
      {stage0_38[417]},
      {stage1_38[182]}
   );
   gpc1_1 gpc4466 (
      {stage0_38[418]},
      {stage1_38[183]}
   );
   gpc1_1 gpc4467 (
      {stage0_38[419]},
      {stage1_38[184]}
   );
   gpc1_1 gpc4468 (
      {stage0_38[420]},
      {stage1_38[185]}
   );
   gpc1_1 gpc4469 (
      {stage0_38[421]},
      {stage1_38[186]}
   );
   gpc1_1 gpc4470 (
      {stage0_38[422]},
      {stage1_38[187]}
   );
   gpc1_1 gpc4471 (
      {stage0_38[423]},
      {stage1_38[188]}
   );
   gpc1_1 gpc4472 (
      {stage0_38[424]},
      {stage1_38[189]}
   );
   gpc1_1 gpc4473 (
      {stage0_38[425]},
      {stage1_38[190]}
   );
   gpc1_1 gpc4474 (
      {stage0_38[426]},
      {stage1_38[191]}
   );
   gpc1_1 gpc4475 (
      {stage0_38[427]},
      {stage1_38[192]}
   );
   gpc1_1 gpc4476 (
      {stage0_38[428]},
      {stage1_38[193]}
   );
   gpc1_1 gpc4477 (
      {stage0_38[429]},
      {stage1_38[194]}
   );
   gpc1_1 gpc4478 (
      {stage0_38[430]},
      {stage1_38[195]}
   );
   gpc1_1 gpc4479 (
      {stage0_38[431]},
      {stage1_38[196]}
   );
   gpc1_1 gpc4480 (
      {stage0_38[432]},
      {stage1_38[197]}
   );
   gpc1_1 gpc4481 (
      {stage0_38[433]},
      {stage1_38[198]}
   );
   gpc1_1 gpc4482 (
      {stage0_38[434]},
      {stage1_38[199]}
   );
   gpc1_1 gpc4483 (
      {stage0_38[435]},
      {stage1_38[200]}
   );
   gpc1_1 gpc4484 (
      {stage0_38[436]},
      {stage1_38[201]}
   );
   gpc1_1 gpc4485 (
      {stage0_38[437]},
      {stage1_38[202]}
   );
   gpc1_1 gpc4486 (
      {stage0_38[438]},
      {stage1_38[203]}
   );
   gpc1_1 gpc4487 (
      {stage0_38[439]},
      {stage1_38[204]}
   );
   gpc1_1 gpc4488 (
      {stage0_38[440]},
      {stage1_38[205]}
   );
   gpc1_1 gpc4489 (
      {stage0_38[441]},
      {stage1_38[206]}
   );
   gpc1_1 gpc4490 (
      {stage0_38[442]},
      {stage1_38[207]}
   );
   gpc1_1 gpc4491 (
      {stage0_38[443]},
      {stage1_38[208]}
   );
   gpc1_1 gpc4492 (
      {stage0_38[444]},
      {stage1_38[209]}
   );
   gpc1_1 gpc4493 (
      {stage0_38[445]},
      {stage1_38[210]}
   );
   gpc1_1 gpc4494 (
      {stage0_38[446]},
      {stage1_38[211]}
   );
   gpc1_1 gpc4495 (
      {stage0_38[447]},
      {stage1_38[212]}
   );
   gpc1_1 gpc4496 (
      {stage0_38[448]},
      {stage1_38[213]}
   );
   gpc1_1 gpc4497 (
      {stage0_38[449]},
      {stage1_38[214]}
   );
   gpc1_1 gpc4498 (
      {stage0_38[450]},
      {stage1_38[215]}
   );
   gpc1_1 gpc4499 (
      {stage0_38[451]},
      {stage1_38[216]}
   );
   gpc1_1 gpc4500 (
      {stage0_38[452]},
      {stage1_38[217]}
   );
   gpc1_1 gpc4501 (
      {stage0_38[453]},
      {stage1_38[218]}
   );
   gpc1_1 gpc4502 (
      {stage0_38[454]},
      {stage1_38[219]}
   );
   gpc1_1 gpc4503 (
      {stage0_38[455]},
      {stage1_38[220]}
   );
   gpc1_1 gpc4504 (
      {stage0_38[456]},
      {stage1_38[221]}
   );
   gpc1_1 gpc4505 (
      {stage0_38[457]},
      {stage1_38[222]}
   );
   gpc1_1 gpc4506 (
      {stage0_38[458]},
      {stage1_38[223]}
   );
   gpc1_1 gpc4507 (
      {stage0_38[459]},
      {stage1_38[224]}
   );
   gpc1_1 gpc4508 (
      {stage0_38[460]},
      {stage1_38[225]}
   );
   gpc1_1 gpc4509 (
      {stage0_38[461]},
      {stage1_38[226]}
   );
   gpc1_1 gpc4510 (
      {stage0_38[462]},
      {stage1_38[227]}
   );
   gpc1_1 gpc4511 (
      {stage0_38[463]},
      {stage1_38[228]}
   );
   gpc1_1 gpc4512 (
      {stage0_38[464]},
      {stage1_38[229]}
   );
   gpc1_1 gpc4513 (
      {stage0_38[465]},
      {stage1_38[230]}
   );
   gpc1_1 gpc4514 (
      {stage0_38[466]},
      {stage1_38[231]}
   );
   gpc1_1 gpc4515 (
      {stage0_38[467]},
      {stage1_38[232]}
   );
   gpc1_1 gpc4516 (
      {stage0_38[468]},
      {stage1_38[233]}
   );
   gpc1_1 gpc4517 (
      {stage0_38[469]},
      {stage1_38[234]}
   );
   gpc1_1 gpc4518 (
      {stage0_38[470]},
      {stage1_38[235]}
   );
   gpc1_1 gpc4519 (
      {stage0_38[471]},
      {stage1_38[236]}
   );
   gpc1_1 gpc4520 (
      {stage0_38[472]},
      {stage1_38[237]}
   );
   gpc1_1 gpc4521 (
      {stage0_38[473]},
      {stage1_38[238]}
   );
   gpc1_1 gpc4522 (
      {stage0_38[474]},
      {stage1_38[239]}
   );
   gpc1_1 gpc4523 (
      {stage0_38[475]},
      {stage1_38[240]}
   );
   gpc1_1 gpc4524 (
      {stage0_38[476]},
      {stage1_38[241]}
   );
   gpc1_1 gpc4525 (
      {stage0_38[477]},
      {stage1_38[242]}
   );
   gpc1_1 gpc4526 (
      {stage0_38[478]},
      {stage1_38[243]}
   );
   gpc1_1 gpc4527 (
      {stage0_38[479]},
      {stage1_38[244]}
   );
   gpc1_1 gpc4528 (
      {stage0_38[480]},
      {stage1_38[245]}
   );
   gpc1_1 gpc4529 (
      {stage0_38[481]},
      {stage1_38[246]}
   );
   gpc1_1 gpc4530 (
      {stage0_38[482]},
      {stage1_38[247]}
   );
   gpc1_1 gpc4531 (
      {stage0_38[483]},
      {stage1_38[248]}
   );
   gpc1_1 gpc4532 (
      {stage0_38[484]},
      {stage1_38[249]}
   );
   gpc1_1 gpc4533 (
      {stage0_38[485]},
      {stage1_38[250]}
   );
   gpc1_1 gpc4534 (
      {stage0_38[486]},
      {stage1_38[251]}
   );
   gpc1_1 gpc4535 (
      {stage0_38[487]},
      {stage1_38[252]}
   );
   gpc1_1 gpc4536 (
      {stage0_38[488]},
      {stage1_38[253]}
   );
   gpc1_1 gpc4537 (
      {stage0_38[489]},
      {stage1_38[254]}
   );
   gpc1_1 gpc4538 (
      {stage0_38[490]},
      {stage1_38[255]}
   );
   gpc1_1 gpc4539 (
      {stage0_38[491]},
      {stage1_38[256]}
   );
   gpc1_1 gpc4540 (
      {stage0_38[492]},
      {stage1_38[257]}
   );
   gpc1_1 gpc4541 (
      {stage0_38[493]},
      {stage1_38[258]}
   );
   gpc1_1 gpc4542 (
      {stage0_38[494]},
      {stage1_38[259]}
   );
   gpc1_1 gpc4543 (
      {stage0_38[495]},
      {stage1_38[260]}
   );
   gpc1_1 gpc4544 (
      {stage0_38[496]},
      {stage1_38[261]}
   );
   gpc1_1 gpc4545 (
      {stage0_38[497]},
      {stage1_38[262]}
   );
   gpc1_1 gpc4546 (
      {stage0_38[498]},
      {stage1_38[263]}
   );
   gpc1_1 gpc4547 (
      {stage0_38[499]},
      {stage1_38[264]}
   );
   gpc1_1 gpc4548 (
      {stage0_38[500]},
      {stage1_38[265]}
   );
   gpc1_1 gpc4549 (
      {stage0_38[501]},
      {stage1_38[266]}
   );
   gpc1_1 gpc4550 (
      {stage0_38[502]},
      {stage1_38[267]}
   );
   gpc1_1 gpc4551 (
      {stage0_38[503]},
      {stage1_38[268]}
   );
   gpc1_1 gpc4552 (
      {stage0_38[504]},
      {stage1_38[269]}
   );
   gpc1_1 gpc4553 (
      {stage0_38[505]},
      {stage1_38[270]}
   );
   gpc1_1 gpc4554 (
      {stage0_38[506]},
      {stage1_38[271]}
   );
   gpc1_1 gpc4555 (
      {stage0_38[507]},
      {stage1_38[272]}
   );
   gpc1_1 gpc4556 (
      {stage0_38[508]},
      {stage1_38[273]}
   );
   gpc1_1 gpc4557 (
      {stage0_38[509]},
      {stage1_38[274]}
   );
   gpc1_1 gpc4558 (
      {stage0_38[510]},
      {stage1_38[275]}
   );
   gpc1_1 gpc4559 (
      {stage0_38[511]},
      {stage1_38[276]}
   );
   gpc1_1 gpc4560 (
      {stage0_39[491]},
      {stage1_39[176]}
   );
   gpc1_1 gpc4561 (
      {stage0_39[492]},
      {stage1_39[177]}
   );
   gpc1_1 gpc4562 (
      {stage0_39[493]},
      {stage1_39[178]}
   );
   gpc1_1 gpc4563 (
      {stage0_39[494]},
      {stage1_39[179]}
   );
   gpc1_1 gpc4564 (
      {stage0_39[495]},
      {stage1_39[180]}
   );
   gpc1_1 gpc4565 (
      {stage0_39[496]},
      {stage1_39[181]}
   );
   gpc1_1 gpc4566 (
      {stage0_39[497]},
      {stage1_39[182]}
   );
   gpc1_1 gpc4567 (
      {stage0_39[498]},
      {stage1_39[183]}
   );
   gpc1_1 gpc4568 (
      {stage0_39[499]},
      {stage1_39[184]}
   );
   gpc1_1 gpc4569 (
      {stage0_39[500]},
      {stage1_39[185]}
   );
   gpc1_1 gpc4570 (
      {stage0_39[501]},
      {stage1_39[186]}
   );
   gpc1_1 gpc4571 (
      {stage0_39[502]},
      {stage1_39[187]}
   );
   gpc1_1 gpc4572 (
      {stage0_39[503]},
      {stage1_39[188]}
   );
   gpc1_1 gpc4573 (
      {stage0_39[504]},
      {stage1_39[189]}
   );
   gpc1_1 gpc4574 (
      {stage0_39[505]},
      {stage1_39[190]}
   );
   gpc1_1 gpc4575 (
      {stage0_39[506]},
      {stage1_39[191]}
   );
   gpc1_1 gpc4576 (
      {stage0_39[507]},
      {stage1_39[192]}
   );
   gpc1_1 gpc4577 (
      {stage0_39[508]},
      {stage1_39[193]}
   );
   gpc1_1 gpc4578 (
      {stage0_39[509]},
      {stage1_39[194]}
   );
   gpc1_1 gpc4579 (
      {stage0_39[510]},
      {stage1_39[195]}
   );
   gpc1_1 gpc4580 (
      {stage0_39[511]},
      {stage1_39[196]}
   );
   gpc1_1 gpc4581 (
      {stage0_40[489]},
      {stage1_40[207]}
   );
   gpc1_1 gpc4582 (
      {stage0_40[490]},
      {stage1_40[208]}
   );
   gpc1_1 gpc4583 (
      {stage0_40[491]},
      {stage1_40[209]}
   );
   gpc1_1 gpc4584 (
      {stage0_40[492]},
      {stage1_40[210]}
   );
   gpc1_1 gpc4585 (
      {stage0_40[493]},
      {stage1_40[211]}
   );
   gpc1_1 gpc4586 (
      {stage0_40[494]},
      {stage1_40[212]}
   );
   gpc1_1 gpc4587 (
      {stage0_40[495]},
      {stage1_40[213]}
   );
   gpc1_1 gpc4588 (
      {stage0_40[496]},
      {stage1_40[214]}
   );
   gpc1_1 gpc4589 (
      {stage0_40[497]},
      {stage1_40[215]}
   );
   gpc1_1 gpc4590 (
      {stage0_40[498]},
      {stage1_40[216]}
   );
   gpc1_1 gpc4591 (
      {stage0_40[499]},
      {stage1_40[217]}
   );
   gpc1_1 gpc4592 (
      {stage0_40[500]},
      {stage1_40[218]}
   );
   gpc1_1 gpc4593 (
      {stage0_40[501]},
      {stage1_40[219]}
   );
   gpc1_1 gpc4594 (
      {stage0_40[502]},
      {stage1_40[220]}
   );
   gpc1_1 gpc4595 (
      {stage0_40[503]},
      {stage1_40[221]}
   );
   gpc1_1 gpc4596 (
      {stage0_40[504]},
      {stage1_40[222]}
   );
   gpc1_1 gpc4597 (
      {stage0_40[505]},
      {stage1_40[223]}
   );
   gpc1_1 gpc4598 (
      {stage0_40[506]},
      {stage1_40[224]}
   );
   gpc1_1 gpc4599 (
      {stage0_40[507]},
      {stage1_40[225]}
   );
   gpc1_1 gpc4600 (
      {stage0_40[508]},
      {stage1_40[226]}
   );
   gpc1_1 gpc4601 (
      {stage0_40[509]},
      {stage1_40[227]}
   );
   gpc1_1 gpc4602 (
      {stage0_40[510]},
      {stage1_40[228]}
   );
   gpc1_1 gpc4603 (
      {stage0_40[511]},
      {stage1_40[229]}
   );
   gpc1_1 gpc4604 (
      {stage0_41[420]},
      {stage1_41[185]}
   );
   gpc1_1 gpc4605 (
      {stage0_41[421]},
      {stage1_41[186]}
   );
   gpc1_1 gpc4606 (
      {stage0_41[422]},
      {stage1_41[187]}
   );
   gpc1_1 gpc4607 (
      {stage0_41[423]},
      {stage1_41[188]}
   );
   gpc1_1 gpc4608 (
      {stage0_41[424]},
      {stage1_41[189]}
   );
   gpc1_1 gpc4609 (
      {stage0_41[425]},
      {stage1_41[190]}
   );
   gpc1_1 gpc4610 (
      {stage0_41[426]},
      {stage1_41[191]}
   );
   gpc1_1 gpc4611 (
      {stage0_41[427]},
      {stage1_41[192]}
   );
   gpc1_1 gpc4612 (
      {stage0_41[428]},
      {stage1_41[193]}
   );
   gpc1_1 gpc4613 (
      {stage0_41[429]},
      {stage1_41[194]}
   );
   gpc1_1 gpc4614 (
      {stage0_41[430]},
      {stage1_41[195]}
   );
   gpc1_1 gpc4615 (
      {stage0_41[431]},
      {stage1_41[196]}
   );
   gpc1_1 gpc4616 (
      {stage0_41[432]},
      {stage1_41[197]}
   );
   gpc1_1 gpc4617 (
      {stage0_41[433]},
      {stage1_41[198]}
   );
   gpc1_1 gpc4618 (
      {stage0_41[434]},
      {stage1_41[199]}
   );
   gpc1_1 gpc4619 (
      {stage0_41[435]},
      {stage1_41[200]}
   );
   gpc1_1 gpc4620 (
      {stage0_41[436]},
      {stage1_41[201]}
   );
   gpc1_1 gpc4621 (
      {stage0_41[437]},
      {stage1_41[202]}
   );
   gpc1_1 gpc4622 (
      {stage0_41[438]},
      {stage1_41[203]}
   );
   gpc1_1 gpc4623 (
      {stage0_41[439]},
      {stage1_41[204]}
   );
   gpc1_1 gpc4624 (
      {stage0_41[440]},
      {stage1_41[205]}
   );
   gpc1_1 gpc4625 (
      {stage0_41[441]},
      {stage1_41[206]}
   );
   gpc1_1 gpc4626 (
      {stage0_41[442]},
      {stage1_41[207]}
   );
   gpc1_1 gpc4627 (
      {stage0_41[443]},
      {stage1_41[208]}
   );
   gpc1_1 gpc4628 (
      {stage0_41[444]},
      {stage1_41[209]}
   );
   gpc1_1 gpc4629 (
      {stage0_41[445]},
      {stage1_41[210]}
   );
   gpc1_1 gpc4630 (
      {stage0_41[446]},
      {stage1_41[211]}
   );
   gpc1_1 gpc4631 (
      {stage0_41[447]},
      {stage1_41[212]}
   );
   gpc1_1 gpc4632 (
      {stage0_41[448]},
      {stage1_41[213]}
   );
   gpc1_1 gpc4633 (
      {stage0_41[449]},
      {stage1_41[214]}
   );
   gpc1_1 gpc4634 (
      {stage0_41[450]},
      {stage1_41[215]}
   );
   gpc1_1 gpc4635 (
      {stage0_41[451]},
      {stage1_41[216]}
   );
   gpc1_1 gpc4636 (
      {stage0_41[452]},
      {stage1_41[217]}
   );
   gpc1_1 gpc4637 (
      {stage0_41[453]},
      {stage1_41[218]}
   );
   gpc1_1 gpc4638 (
      {stage0_41[454]},
      {stage1_41[219]}
   );
   gpc1_1 gpc4639 (
      {stage0_41[455]},
      {stage1_41[220]}
   );
   gpc1_1 gpc4640 (
      {stage0_41[456]},
      {stage1_41[221]}
   );
   gpc1_1 gpc4641 (
      {stage0_41[457]},
      {stage1_41[222]}
   );
   gpc1_1 gpc4642 (
      {stage0_41[458]},
      {stage1_41[223]}
   );
   gpc1_1 gpc4643 (
      {stage0_41[459]},
      {stage1_41[224]}
   );
   gpc1_1 gpc4644 (
      {stage0_41[460]},
      {stage1_41[225]}
   );
   gpc1_1 gpc4645 (
      {stage0_41[461]},
      {stage1_41[226]}
   );
   gpc1_1 gpc4646 (
      {stage0_41[462]},
      {stage1_41[227]}
   );
   gpc1_1 gpc4647 (
      {stage0_41[463]},
      {stage1_41[228]}
   );
   gpc1_1 gpc4648 (
      {stage0_41[464]},
      {stage1_41[229]}
   );
   gpc1_1 gpc4649 (
      {stage0_41[465]},
      {stage1_41[230]}
   );
   gpc1_1 gpc4650 (
      {stage0_41[466]},
      {stage1_41[231]}
   );
   gpc1_1 gpc4651 (
      {stage0_41[467]},
      {stage1_41[232]}
   );
   gpc1_1 gpc4652 (
      {stage0_41[468]},
      {stage1_41[233]}
   );
   gpc1_1 gpc4653 (
      {stage0_41[469]},
      {stage1_41[234]}
   );
   gpc1_1 gpc4654 (
      {stage0_41[470]},
      {stage1_41[235]}
   );
   gpc1_1 gpc4655 (
      {stage0_41[471]},
      {stage1_41[236]}
   );
   gpc1_1 gpc4656 (
      {stage0_41[472]},
      {stage1_41[237]}
   );
   gpc1_1 gpc4657 (
      {stage0_41[473]},
      {stage1_41[238]}
   );
   gpc1_1 gpc4658 (
      {stage0_41[474]},
      {stage1_41[239]}
   );
   gpc1_1 gpc4659 (
      {stage0_41[475]},
      {stage1_41[240]}
   );
   gpc1_1 gpc4660 (
      {stage0_41[476]},
      {stage1_41[241]}
   );
   gpc1_1 gpc4661 (
      {stage0_41[477]},
      {stage1_41[242]}
   );
   gpc1_1 gpc4662 (
      {stage0_41[478]},
      {stage1_41[243]}
   );
   gpc1_1 gpc4663 (
      {stage0_41[479]},
      {stage1_41[244]}
   );
   gpc1_1 gpc4664 (
      {stage0_41[480]},
      {stage1_41[245]}
   );
   gpc1_1 gpc4665 (
      {stage0_41[481]},
      {stage1_41[246]}
   );
   gpc1_1 gpc4666 (
      {stage0_41[482]},
      {stage1_41[247]}
   );
   gpc1_1 gpc4667 (
      {stage0_41[483]},
      {stage1_41[248]}
   );
   gpc1_1 gpc4668 (
      {stage0_41[484]},
      {stage1_41[249]}
   );
   gpc1_1 gpc4669 (
      {stage0_41[485]},
      {stage1_41[250]}
   );
   gpc1_1 gpc4670 (
      {stage0_41[486]},
      {stage1_41[251]}
   );
   gpc1_1 gpc4671 (
      {stage0_41[487]},
      {stage1_41[252]}
   );
   gpc1_1 gpc4672 (
      {stage0_41[488]},
      {stage1_41[253]}
   );
   gpc1_1 gpc4673 (
      {stage0_41[489]},
      {stage1_41[254]}
   );
   gpc1_1 gpc4674 (
      {stage0_41[490]},
      {stage1_41[255]}
   );
   gpc1_1 gpc4675 (
      {stage0_41[491]},
      {stage1_41[256]}
   );
   gpc1_1 gpc4676 (
      {stage0_41[492]},
      {stage1_41[257]}
   );
   gpc1_1 gpc4677 (
      {stage0_41[493]},
      {stage1_41[258]}
   );
   gpc1_1 gpc4678 (
      {stage0_41[494]},
      {stage1_41[259]}
   );
   gpc1_1 gpc4679 (
      {stage0_41[495]},
      {stage1_41[260]}
   );
   gpc1_1 gpc4680 (
      {stage0_41[496]},
      {stage1_41[261]}
   );
   gpc1_1 gpc4681 (
      {stage0_41[497]},
      {stage1_41[262]}
   );
   gpc1_1 gpc4682 (
      {stage0_41[498]},
      {stage1_41[263]}
   );
   gpc1_1 gpc4683 (
      {stage0_41[499]},
      {stage1_41[264]}
   );
   gpc1_1 gpc4684 (
      {stage0_41[500]},
      {stage1_41[265]}
   );
   gpc1_1 gpc4685 (
      {stage0_41[501]},
      {stage1_41[266]}
   );
   gpc1_1 gpc4686 (
      {stage0_41[502]},
      {stage1_41[267]}
   );
   gpc1_1 gpc4687 (
      {stage0_41[503]},
      {stage1_41[268]}
   );
   gpc1_1 gpc4688 (
      {stage0_41[504]},
      {stage1_41[269]}
   );
   gpc1_1 gpc4689 (
      {stage0_41[505]},
      {stage1_41[270]}
   );
   gpc1_1 gpc4690 (
      {stage0_41[506]},
      {stage1_41[271]}
   );
   gpc1_1 gpc4691 (
      {stage0_41[507]},
      {stage1_41[272]}
   );
   gpc1_1 gpc4692 (
      {stage0_41[508]},
      {stage1_41[273]}
   );
   gpc1_1 gpc4693 (
      {stage0_41[509]},
      {stage1_41[274]}
   );
   gpc1_1 gpc4694 (
      {stage0_41[510]},
      {stage1_41[275]}
   );
   gpc1_1 gpc4695 (
      {stage0_41[511]},
      {stage1_41[276]}
   );
   gpc1_1 gpc4696 (
      {stage0_42[451]},
      {stage1_42[168]}
   );
   gpc1_1 gpc4697 (
      {stage0_42[452]},
      {stage1_42[169]}
   );
   gpc1_1 gpc4698 (
      {stage0_42[453]},
      {stage1_42[170]}
   );
   gpc1_1 gpc4699 (
      {stage0_42[454]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4700 (
      {stage0_42[455]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4701 (
      {stage0_42[456]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4702 (
      {stage0_42[457]},
      {stage1_42[174]}
   );
   gpc1_1 gpc4703 (
      {stage0_42[458]},
      {stage1_42[175]}
   );
   gpc1_1 gpc4704 (
      {stage0_42[459]},
      {stage1_42[176]}
   );
   gpc1_1 gpc4705 (
      {stage0_42[460]},
      {stage1_42[177]}
   );
   gpc1_1 gpc4706 (
      {stage0_42[461]},
      {stage1_42[178]}
   );
   gpc1_1 gpc4707 (
      {stage0_42[462]},
      {stage1_42[179]}
   );
   gpc1_1 gpc4708 (
      {stage0_42[463]},
      {stage1_42[180]}
   );
   gpc1_1 gpc4709 (
      {stage0_42[464]},
      {stage1_42[181]}
   );
   gpc1_1 gpc4710 (
      {stage0_42[465]},
      {stage1_42[182]}
   );
   gpc1_1 gpc4711 (
      {stage0_42[466]},
      {stage1_42[183]}
   );
   gpc1_1 gpc4712 (
      {stage0_42[467]},
      {stage1_42[184]}
   );
   gpc1_1 gpc4713 (
      {stage0_42[468]},
      {stage1_42[185]}
   );
   gpc1_1 gpc4714 (
      {stage0_42[469]},
      {stage1_42[186]}
   );
   gpc1_1 gpc4715 (
      {stage0_42[470]},
      {stage1_42[187]}
   );
   gpc1_1 gpc4716 (
      {stage0_42[471]},
      {stage1_42[188]}
   );
   gpc1_1 gpc4717 (
      {stage0_42[472]},
      {stage1_42[189]}
   );
   gpc1_1 gpc4718 (
      {stage0_42[473]},
      {stage1_42[190]}
   );
   gpc1_1 gpc4719 (
      {stage0_42[474]},
      {stage1_42[191]}
   );
   gpc1_1 gpc4720 (
      {stage0_42[475]},
      {stage1_42[192]}
   );
   gpc1_1 gpc4721 (
      {stage0_42[476]},
      {stage1_42[193]}
   );
   gpc1_1 gpc4722 (
      {stage0_42[477]},
      {stage1_42[194]}
   );
   gpc1_1 gpc4723 (
      {stage0_42[478]},
      {stage1_42[195]}
   );
   gpc1_1 gpc4724 (
      {stage0_42[479]},
      {stage1_42[196]}
   );
   gpc1_1 gpc4725 (
      {stage0_42[480]},
      {stage1_42[197]}
   );
   gpc1_1 gpc4726 (
      {stage0_42[481]},
      {stage1_42[198]}
   );
   gpc1_1 gpc4727 (
      {stage0_42[482]},
      {stage1_42[199]}
   );
   gpc1_1 gpc4728 (
      {stage0_42[483]},
      {stage1_42[200]}
   );
   gpc1_1 gpc4729 (
      {stage0_42[484]},
      {stage1_42[201]}
   );
   gpc1_1 gpc4730 (
      {stage0_42[485]},
      {stage1_42[202]}
   );
   gpc1_1 gpc4731 (
      {stage0_42[486]},
      {stage1_42[203]}
   );
   gpc1_1 gpc4732 (
      {stage0_42[487]},
      {stage1_42[204]}
   );
   gpc1_1 gpc4733 (
      {stage0_42[488]},
      {stage1_42[205]}
   );
   gpc1_1 gpc4734 (
      {stage0_42[489]},
      {stage1_42[206]}
   );
   gpc1_1 gpc4735 (
      {stage0_42[490]},
      {stage1_42[207]}
   );
   gpc1_1 gpc4736 (
      {stage0_42[491]},
      {stage1_42[208]}
   );
   gpc1_1 gpc4737 (
      {stage0_42[492]},
      {stage1_42[209]}
   );
   gpc1_1 gpc4738 (
      {stage0_42[493]},
      {stage1_42[210]}
   );
   gpc1_1 gpc4739 (
      {stage0_42[494]},
      {stage1_42[211]}
   );
   gpc1_1 gpc4740 (
      {stage0_42[495]},
      {stage1_42[212]}
   );
   gpc1_1 gpc4741 (
      {stage0_42[496]},
      {stage1_42[213]}
   );
   gpc1_1 gpc4742 (
      {stage0_42[497]},
      {stage1_42[214]}
   );
   gpc1_1 gpc4743 (
      {stage0_42[498]},
      {stage1_42[215]}
   );
   gpc1_1 gpc4744 (
      {stage0_42[499]},
      {stage1_42[216]}
   );
   gpc1_1 gpc4745 (
      {stage0_42[500]},
      {stage1_42[217]}
   );
   gpc1_1 gpc4746 (
      {stage0_42[501]},
      {stage1_42[218]}
   );
   gpc1_1 gpc4747 (
      {stage0_42[502]},
      {stage1_42[219]}
   );
   gpc1_1 gpc4748 (
      {stage0_42[503]},
      {stage1_42[220]}
   );
   gpc1_1 gpc4749 (
      {stage0_42[504]},
      {stage1_42[221]}
   );
   gpc1_1 gpc4750 (
      {stage0_42[505]},
      {stage1_42[222]}
   );
   gpc1_1 gpc4751 (
      {stage0_42[506]},
      {stage1_42[223]}
   );
   gpc1_1 gpc4752 (
      {stage0_42[507]},
      {stage1_42[224]}
   );
   gpc1_1 gpc4753 (
      {stage0_42[508]},
      {stage1_42[225]}
   );
   gpc1_1 gpc4754 (
      {stage0_42[509]},
      {stage1_42[226]}
   );
   gpc1_1 gpc4755 (
      {stage0_42[510]},
      {stage1_42[227]}
   );
   gpc1_1 gpc4756 (
      {stage0_42[511]},
      {stage1_42[228]}
   );
   gpc1_1 gpc4757 (
      {stage0_43[475]},
      {stage1_43[207]}
   );
   gpc1_1 gpc4758 (
      {stage0_43[476]},
      {stage1_43[208]}
   );
   gpc1_1 gpc4759 (
      {stage0_43[477]},
      {stage1_43[209]}
   );
   gpc1_1 gpc4760 (
      {stage0_43[478]},
      {stage1_43[210]}
   );
   gpc1_1 gpc4761 (
      {stage0_43[479]},
      {stage1_43[211]}
   );
   gpc1_1 gpc4762 (
      {stage0_43[480]},
      {stage1_43[212]}
   );
   gpc1_1 gpc4763 (
      {stage0_43[481]},
      {stage1_43[213]}
   );
   gpc1_1 gpc4764 (
      {stage0_43[482]},
      {stage1_43[214]}
   );
   gpc1_1 gpc4765 (
      {stage0_43[483]},
      {stage1_43[215]}
   );
   gpc1_1 gpc4766 (
      {stage0_43[484]},
      {stage1_43[216]}
   );
   gpc1_1 gpc4767 (
      {stage0_43[485]},
      {stage1_43[217]}
   );
   gpc1_1 gpc4768 (
      {stage0_43[486]},
      {stage1_43[218]}
   );
   gpc1_1 gpc4769 (
      {stage0_43[487]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4770 (
      {stage0_43[488]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4771 (
      {stage0_43[489]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4772 (
      {stage0_43[490]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4773 (
      {stage0_43[491]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4774 (
      {stage0_43[492]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4775 (
      {stage0_43[493]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4776 (
      {stage0_43[494]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4777 (
      {stage0_43[495]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4778 (
      {stage0_43[496]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4779 (
      {stage0_43[497]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4780 (
      {stage0_43[498]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4781 (
      {stage0_43[499]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4782 (
      {stage0_43[500]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4783 (
      {stage0_43[501]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4784 (
      {stage0_43[502]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4785 (
      {stage0_43[503]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4786 (
      {stage0_43[504]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4787 (
      {stage0_43[505]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4788 (
      {stage0_43[506]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4789 (
      {stage0_43[507]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4790 (
      {stage0_43[508]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4791 (
      {stage0_43[509]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4792 (
      {stage0_43[510]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4793 (
      {stage0_43[511]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4794 (
      {stage0_44[448]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4795 (
      {stage0_44[449]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4796 (
      {stage0_44[450]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4797 (
      {stage0_44[451]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4798 (
      {stage0_44[452]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4799 (
      {stage0_44[453]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4800 (
      {stage0_44[454]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4801 (
      {stage0_44[455]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4802 (
      {stage0_44[456]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4803 (
      {stage0_44[457]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4804 (
      {stage0_44[458]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4805 (
      {stage0_44[459]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4806 (
      {stage0_44[460]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4807 (
      {stage0_44[461]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4808 (
      {stage0_44[462]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4809 (
      {stage0_44[463]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4810 (
      {stage0_44[464]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4811 (
      {stage0_44[465]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4812 (
      {stage0_44[466]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4813 (
      {stage0_44[467]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4814 (
      {stage0_44[468]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4815 (
      {stage0_44[469]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4816 (
      {stage0_44[470]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4817 (
      {stage0_44[471]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4818 (
      {stage0_44[472]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4819 (
      {stage0_44[473]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4820 (
      {stage0_44[474]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4821 (
      {stage0_44[475]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4822 (
      {stage0_44[476]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4823 (
      {stage0_44[477]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4824 (
      {stage0_44[478]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4825 (
      {stage0_44[479]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4826 (
      {stage0_44[480]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4827 (
      {stage0_44[481]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4828 (
      {stage0_44[482]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4829 (
      {stage0_44[483]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4830 (
      {stage0_44[484]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4831 (
      {stage0_44[485]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4832 (
      {stage0_44[486]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4833 (
      {stage0_44[487]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4834 (
      {stage0_44[488]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4835 (
      {stage0_44[489]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4836 (
      {stage0_44[490]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4837 (
      {stage0_44[491]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4838 (
      {stage0_44[492]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4839 (
      {stage0_44[493]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4840 (
      {stage0_44[494]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4841 (
      {stage0_44[495]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4842 (
      {stage0_44[496]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4843 (
      {stage0_44[497]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4844 (
      {stage0_44[498]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4845 (
      {stage0_44[499]},
      {stage1_44[256]}
   );
   gpc1_1 gpc4846 (
      {stage0_44[500]},
      {stage1_44[257]}
   );
   gpc1_1 gpc4847 (
      {stage0_44[501]},
      {stage1_44[258]}
   );
   gpc1_1 gpc4848 (
      {stage0_44[502]},
      {stage1_44[259]}
   );
   gpc1_1 gpc4849 (
      {stage0_44[503]},
      {stage1_44[260]}
   );
   gpc1_1 gpc4850 (
      {stage0_44[504]},
      {stage1_44[261]}
   );
   gpc1_1 gpc4851 (
      {stage0_44[505]},
      {stage1_44[262]}
   );
   gpc1_1 gpc4852 (
      {stage0_44[506]},
      {stage1_44[263]}
   );
   gpc1_1 gpc4853 (
      {stage0_44[507]},
      {stage1_44[264]}
   );
   gpc1_1 gpc4854 (
      {stage0_44[508]},
      {stage1_44[265]}
   );
   gpc1_1 gpc4855 (
      {stage0_44[509]},
      {stage1_44[266]}
   );
   gpc1_1 gpc4856 (
      {stage0_44[510]},
      {stage1_44[267]}
   );
   gpc1_1 gpc4857 (
      {stage0_44[511]},
      {stage1_44[268]}
   );
   gpc1_1 gpc4858 (
      {stage0_45[498]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4859 (
      {stage0_45[499]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4860 (
      {stage0_45[500]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4861 (
      {stage0_45[501]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4862 (
      {stage0_45[502]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4863 (
      {stage0_45[503]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4864 (
      {stage0_45[504]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4865 (
      {stage0_45[505]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4866 (
      {stage0_45[506]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4867 (
      {stage0_45[507]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4868 (
      {stage0_45[508]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4869 (
      {stage0_45[509]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4870 (
      {stage0_45[510]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4871 (
      {stage0_45[511]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4872 (
      {stage0_46[388]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4873 (
      {stage0_46[389]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4874 (
      {stage0_46[390]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4875 (
      {stage0_46[391]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4876 (
      {stage0_46[392]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4877 (
      {stage0_46[393]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4878 (
      {stage0_46[394]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4879 (
      {stage0_46[395]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4880 (
      {stage0_46[396]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4881 (
      {stage0_46[397]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4882 (
      {stage0_46[398]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4883 (
      {stage0_46[399]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4884 (
      {stage0_46[400]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4885 (
      {stage0_46[401]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4886 (
      {stage0_46[402]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4887 (
      {stage0_46[403]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4888 (
      {stage0_46[404]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4889 (
      {stage0_46[405]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4890 (
      {stage0_46[406]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4891 (
      {stage0_46[407]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4892 (
      {stage0_46[408]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4893 (
      {stage0_46[409]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4894 (
      {stage0_46[410]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4895 (
      {stage0_46[411]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4896 (
      {stage0_46[412]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4897 (
      {stage0_46[413]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4898 (
      {stage0_46[414]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4899 (
      {stage0_46[415]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4900 (
      {stage0_46[416]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4901 (
      {stage0_46[417]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4902 (
      {stage0_46[418]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4903 (
      {stage0_46[419]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4904 (
      {stage0_46[420]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4905 (
      {stage0_46[421]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4906 (
      {stage0_46[422]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4907 (
      {stage0_46[423]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4908 (
      {stage0_46[424]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4909 (
      {stage0_46[425]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4910 (
      {stage0_46[426]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4911 (
      {stage0_46[427]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4912 (
      {stage0_46[428]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4913 (
      {stage0_46[429]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4914 (
      {stage0_46[430]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4915 (
      {stage0_46[431]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4916 (
      {stage0_46[432]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4917 (
      {stage0_46[433]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4918 (
      {stage0_46[434]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4919 (
      {stage0_46[435]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4920 (
      {stage0_46[436]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4921 (
      {stage0_46[437]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4922 (
      {stage0_46[438]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4923 (
      {stage0_46[439]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4924 (
      {stage0_46[440]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4925 (
      {stage0_46[441]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4926 (
      {stage0_46[442]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4927 (
      {stage0_46[443]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4928 (
      {stage0_46[444]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4929 (
      {stage0_46[445]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4930 (
      {stage0_46[446]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4931 (
      {stage0_46[447]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4932 (
      {stage0_46[448]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4933 (
      {stage0_46[449]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4934 (
      {stage0_46[450]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4935 (
      {stage0_46[451]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4936 (
      {stage0_46[452]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4937 (
      {stage0_46[453]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4938 (
      {stage0_46[454]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4939 (
      {stage0_46[455]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4940 (
      {stage0_46[456]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4941 (
      {stage0_46[457]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4942 (
      {stage0_46[458]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4943 (
      {stage0_46[459]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4944 (
      {stage0_46[460]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4945 (
      {stage0_46[461]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4946 (
      {stage0_46[462]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4947 (
      {stage0_46[463]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4948 (
      {stage0_46[464]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4949 (
      {stage0_46[465]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4950 (
      {stage0_46[466]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4951 (
      {stage0_46[467]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4952 (
      {stage0_46[468]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4953 (
      {stage0_46[469]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4954 (
      {stage0_46[470]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4955 (
      {stage0_46[471]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4956 (
      {stage0_46[472]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4957 (
      {stage0_46[473]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4958 (
      {stage0_46[474]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4959 (
      {stage0_46[475]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4960 (
      {stage0_46[476]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4961 (
      {stage0_46[477]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4962 (
      {stage0_46[478]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4963 (
      {stage0_46[479]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4964 (
      {stage0_46[480]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4965 (
      {stage0_46[481]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4966 (
      {stage0_46[482]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4967 (
      {stage0_46[483]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4968 (
      {stage0_46[484]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4969 (
      {stage0_46[485]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4970 (
      {stage0_46[486]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4971 (
      {stage0_46[487]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4972 (
      {stage0_46[488]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4973 (
      {stage0_46[489]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4974 (
      {stage0_46[490]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4975 (
      {stage0_46[491]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4976 (
      {stage0_46[492]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4977 (
      {stage0_46[493]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4978 (
      {stage0_46[494]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4979 (
      {stage0_46[495]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4980 (
      {stage0_46[496]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4981 (
      {stage0_46[497]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4982 (
      {stage0_46[498]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4983 (
      {stage0_46[499]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4984 (
      {stage0_46[500]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4985 (
      {stage0_46[501]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4986 (
      {stage0_46[502]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4987 (
      {stage0_46[503]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4988 (
      {stage0_46[504]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4989 (
      {stage0_46[505]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4990 (
      {stage0_46[506]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4991 (
      {stage0_46[507]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4992 (
      {stage0_46[508]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4993 (
      {stage0_46[509]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4994 (
      {stage0_46[510]},
      {stage1_46[298]}
   );
   gpc1_1 gpc4995 (
      {stage0_46[511]},
      {stage1_46[299]}
   );
   gpc1_1 gpc4996 (
      {stage0_47[437]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4997 (
      {stage0_47[438]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4998 (
      {stage0_47[439]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4999 (
      {stage0_47[440]},
      {stage1_47[206]}
   );
   gpc1_1 gpc5000 (
      {stage0_47[441]},
      {stage1_47[207]}
   );
   gpc1_1 gpc5001 (
      {stage0_47[442]},
      {stage1_47[208]}
   );
   gpc1_1 gpc5002 (
      {stage0_47[443]},
      {stage1_47[209]}
   );
   gpc1_1 gpc5003 (
      {stage0_47[444]},
      {stage1_47[210]}
   );
   gpc1_1 gpc5004 (
      {stage0_47[445]},
      {stage1_47[211]}
   );
   gpc1_1 gpc5005 (
      {stage0_47[446]},
      {stage1_47[212]}
   );
   gpc1_1 gpc5006 (
      {stage0_47[447]},
      {stage1_47[213]}
   );
   gpc1_1 gpc5007 (
      {stage0_47[448]},
      {stage1_47[214]}
   );
   gpc1_1 gpc5008 (
      {stage0_47[449]},
      {stage1_47[215]}
   );
   gpc1_1 gpc5009 (
      {stage0_47[450]},
      {stage1_47[216]}
   );
   gpc1_1 gpc5010 (
      {stage0_47[451]},
      {stage1_47[217]}
   );
   gpc1_1 gpc5011 (
      {stage0_47[452]},
      {stage1_47[218]}
   );
   gpc1_1 gpc5012 (
      {stage0_47[453]},
      {stage1_47[219]}
   );
   gpc1_1 gpc5013 (
      {stage0_47[454]},
      {stage1_47[220]}
   );
   gpc1_1 gpc5014 (
      {stage0_47[455]},
      {stage1_47[221]}
   );
   gpc1_1 gpc5015 (
      {stage0_47[456]},
      {stage1_47[222]}
   );
   gpc1_1 gpc5016 (
      {stage0_47[457]},
      {stage1_47[223]}
   );
   gpc1_1 gpc5017 (
      {stage0_47[458]},
      {stage1_47[224]}
   );
   gpc1_1 gpc5018 (
      {stage0_47[459]},
      {stage1_47[225]}
   );
   gpc1_1 gpc5019 (
      {stage0_47[460]},
      {stage1_47[226]}
   );
   gpc1_1 gpc5020 (
      {stage0_47[461]},
      {stage1_47[227]}
   );
   gpc1_1 gpc5021 (
      {stage0_47[462]},
      {stage1_47[228]}
   );
   gpc1_1 gpc5022 (
      {stage0_47[463]},
      {stage1_47[229]}
   );
   gpc1_1 gpc5023 (
      {stage0_47[464]},
      {stage1_47[230]}
   );
   gpc1_1 gpc5024 (
      {stage0_47[465]},
      {stage1_47[231]}
   );
   gpc1_1 gpc5025 (
      {stage0_47[466]},
      {stage1_47[232]}
   );
   gpc1_1 gpc5026 (
      {stage0_47[467]},
      {stage1_47[233]}
   );
   gpc1_1 gpc5027 (
      {stage0_47[468]},
      {stage1_47[234]}
   );
   gpc1_1 gpc5028 (
      {stage0_47[469]},
      {stage1_47[235]}
   );
   gpc1_1 gpc5029 (
      {stage0_47[470]},
      {stage1_47[236]}
   );
   gpc1_1 gpc5030 (
      {stage0_47[471]},
      {stage1_47[237]}
   );
   gpc1_1 gpc5031 (
      {stage0_47[472]},
      {stage1_47[238]}
   );
   gpc1_1 gpc5032 (
      {stage0_47[473]},
      {stage1_47[239]}
   );
   gpc1_1 gpc5033 (
      {stage0_47[474]},
      {stage1_47[240]}
   );
   gpc1_1 gpc5034 (
      {stage0_47[475]},
      {stage1_47[241]}
   );
   gpc1_1 gpc5035 (
      {stage0_47[476]},
      {stage1_47[242]}
   );
   gpc1_1 gpc5036 (
      {stage0_47[477]},
      {stage1_47[243]}
   );
   gpc1_1 gpc5037 (
      {stage0_47[478]},
      {stage1_47[244]}
   );
   gpc1_1 gpc5038 (
      {stage0_47[479]},
      {stage1_47[245]}
   );
   gpc1_1 gpc5039 (
      {stage0_47[480]},
      {stage1_47[246]}
   );
   gpc1_1 gpc5040 (
      {stage0_47[481]},
      {stage1_47[247]}
   );
   gpc1_1 gpc5041 (
      {stage0_47[482]},
      {stage1_47[248]}
   );
   gpc1_1 gpc5042 (
      {stage0_47[483]},
      {stage1_47[249]}
   );
   gpc1_1 gpc5043 (
      {stage0_47[484]},
      {stage1_47[250]}
   );
   gpc1_1 gpc5044 (
      {stage0_47[485]},
      {stage1_47[251]}
   );
   gpc1_1 gpc5045 (
      {stage0_47[486]},
      {stage1_47[252]}
   );
   gpc1_1 gpc5046 (
      {stage0_47[487]},
      {stage1_47[253]}
   );
   gpc1_1 gpc5047 (
      {stage0_47[488]},
      {stage1_47[254]}
   );
   gpc1_1 gpc5048 (
      {stage0_47[489]},
      {stage1_47[255]}
   );
   gpc1_1 gpc5049 (
      {stage0_47[490]},
      {stage1_47[256]}
   );
   gpc1_1 gpc5050 (
      {stage0_47[491]},
      {stage1_47[257]}
   );
   gpc1_1 gpc5051 (
      {stage0_47[492]},
      {stage1_47[258]}
   );
   gpc1_1 gpc5052 (
      {stage0_47[493]},
      {stage1_47[259]}
   );
   gpc1_1 gpc5053 (
      {stage0_47[494]},
      {stage1_47[260]}
   );
   gpc1_1 gpc5054 (
      {stage0_47[495]},
      {stage1_47[261]}
   );
   gpc1_1 gpc5055 (
      {stage0_47[496]},
      {stage1_47[262]}
   );
   gpc1_1 gpc5056 (
      {stage0_47[497]},
      {stage1_47[263]}
   );
   gpc1_1 gpc5057 (
      {stage0_47[498]},
      {stage1_47[264]}
   );
   gpc1_1 gpc5058 (
      {stage0_47[499]},
      {stage1_47[265]}
   );
   gpc1_1 gpc5059 (
      {stage0_47[500]},
      {stage1_47[266]}
   );
   gpc1_1 gpc5060 (
      {stage0_47[501]},
      {stage1_47[267]}
   );
   gpc1_1 gpc5061 (
      {stage0_47[502]},
      {stage1_47[268]}
   );
   gpc1_1 gpc5062 (
      {stage0_47[503]},
      {stage1_47[269]}
   );
   gpc1_1 gpc5063 (
      {stage0_47[504]},
      {stage1_47[270]}
   );
   gpc1_1 gpc5064 (
      {stage0_47[505]},
      {stage1_47[271]}
   );
   gpc1_1 gpc5065 (
      {stage0_47[506]},
      {stage1_47[272]}
   );
   gpc1_1 gpc5066 (
      {stage0_47[507]},
      {stage1_47[273]}
   );
   gpc1_1 gpc5067 (
      {stage0_47[508]},
      {stage1_47[274]}
   );
   gpc1_1 gpc5068 (
      {stage0_47[509]},
      {stage1_47[275]}
   );
   gpc1_1 gpc5069 (
      {stage0_47[510]},
      {stage1_47[276]}
   );
   gpc1_1 gpc5070 (
      {stage0_47[511]},
      {stage1_47[277]}
   );
   gpc1_1 gpc5071 (
      {stage0_48[495]},
      {stage1_48[194]}
   );
   gpc1_1 gpc5072 (
      {stage0_48[496]},
      {stage1_48[195]}
   );
   gpc1_1 gpc5073 (
      {stage0_48[497]},
      {stage1_48[196]}
   );
   gpc1_1 gpc5074 (
      {stage0_48[498]},
      {stage1_48[197]}
   );
   gpc1_1 gpc5075 (
      {stage0_48[499]},
      {stage1_48[198]}
   );
   gpc1_1 gpc5076 (
      {stage0_48[500]},
      {stage1_48[199]}
   );
   gpc1_1 gpc5077 (
      {stage0_48[501]},
      {stage1_48[200]}
   );
   gpc1_1 gpc5078 (
      {stage0_48[502]},
      {stage1_48[201]}
   );
   gpc1_1 gpc5079 (
      {stage0_48[503]},
      {stage1_48[202]}
   );
   gpc1_1 gpc5080 (
      {stage0_48[504]},
      {stage1_48[203]}
   );
   gpc1_1 gpc5081 (
      {stage0_48[505]},
      {stage1_48[204]}
   );
   gpc1_1 gpc5082 (
      {stage0_48[506]},
      {stage1_48[205]}
   );
   gpc1_1 gpc5083 (
      {stage0_48[507]},
      {stage1_48[206]}
   );
   gpc1_1 gpc5084 (
      {stage0_48[508]},
      {stage1_48[207]}
   );
   gpc1_1 gpc5085 (
      {stage0_48[509]},
      {stage1_48[208]}
   );
   gpc1_1 gpc5086 (
      {stage0_48[510]},
      {stage1_48[209]}
   );
   gpc1_1 gpc5087 (
      {stage0_48[511]},
      {stage1_48[210]}
   );
   gpc1_1 gpc5088 (
      {stage0_49[444]},
      {stage1_49[174]}
   );
   gpc1_1 gpc5089 (
      {stage0_49[445]},
      {stage1_49[175]}
   );
   gpc1_1 gpc5090 (
      {stage0_49[446]},
      {stage1_49[176]}
   );
   gpc1_1 gpc5091 (
      {stage0_49[447]},
      {stage1_49[177]}
   );
   gpc1_1 gpc5092 (
      {stage0_49[448]},
      {stage1_49[178]}
   );
   gpc1_1 gpc5093 (
      {stage0_49[449]},
      {stage1_49[179]}
   );
   gpc1_1 gpc5094 (
      {stage0_49[450]},
      {stage1_49[180]}
   );
   gpc1_1 gpc5095 (
      {stage0_49[451]},
      {stage1_49[181]}
   );
   gpc1_1 gpc5096 (
      {stage0_49[452]},
      {stage1_49[182]}
   );
   gpc1_1 gpc5097 (
      {stage0_49[453]},
      {stage1_49[183]}
   );
   gpc1_1 gpc5098 (
      {stage0_49[454]},
      {stage1_49[184]}
   );
   gpc1_1 gpc5099 (
      {stage0_49[455]},
      {stage1_49[185]}
   );
   gpc1_1 gpc5100 (
      {stage0_49[456]},
      {stage1_49[186]}
   );
   gpc1_1 gpc5101 (
      {stage0_49[457]},
      {stage1_49[187]}
   );
   gpc1_1 gpc5102 (
      {stage0_49[458]},
      {stage1_49[188]}
   );
   gpc1_1 gpc5103 (
      {stage0_49[459]},
      {stage1_49[189]}
   );
   gpc1_1 gpc5104 (
      {stage0_49[460]},
      {stage1_49[190]}
   );
   gpc1_1 gpc5105 (
      {stage0_49[461]},
      {stage1_49[191]}
   );
   gpc1_1 gpc5106 (
      {stage0_49[462]},
      {stage1_49[192]}
   );
   gpc1_1 gpc5107 (
      {stage0_49[463]},
      {stage1_49[193]}
   );
   gpc1_1 gpc5108 (
      {stage0_49[464]},
      {stage1_49[194]}
   );
   gpc1_1 gpc5109 (
      {stage0_49[465]},
      {stage1_49[195]}
   );
   gpc1_1 gpc5110 (
      {stage0_49[466]},
      {stage1_49[196]}
   );
   gpc1_1 gpc5111 (
      {stage0_49[467]},
      {stage1_49[197]}
   );
   gpc1_1 gpc5112 (
      {stage0_49[468]},
      {stage1_49[198]}
   );
   gpc1_1 gpc5113 (
      {stage0_49[469]},
      {stage1_49[199]}
   );
   gpc1_1 gpc5114 (
      {stage0_49[470]},
      {stage1_49[200]}
   );
   gpc1_1 gpc5115 (
      {stage0_49[471]},
      {stage1_49[201]}
   );
   gpc1_1 gpc5116 (
      {stage0_49[472]},
      {stage1_49[202]}
   );
   gpc1_1 gpc5117 (
      {stage0_49[473]},
      {stage1_49[203]}
   );
   gpc1_1 gpc5118 (
      {stage0_49[474]},
      {stage1_49[204]}
   );
   gpc1_1 gpc5119 (
      {stage0_49[475]},
      {stage1_49[205]}
   );
   gpc1_1 gpc5120 (
      {stage0_49[476]},
      {stage1_49[206]}
   );
   gpc1_1 gpc5121 (
      {stage0_49[477]},
      {stage1_49[207]}
   );
   gpc1_1 gpc5122 (
      {stage0_49[478]},
      {stage1_49[208]}
   );
   gpc1_1 gpc5123 (
      {stage0_49[479]},
      {stage1_49[209]}
   );
   gpc1_1 gpc5124 (
      {stage0_49[480]},
      {stage1_49[210]}
   );
   gpc1_1 gpc5125 (
      {stage0_49[481]},
      {stage1_49[211]}
   );
   gpc1_1 gpc5126 (
      {stage0_49[482]},
      {stage1_49[212]}
   );
   gpc1_1 gpc5127 (
      {stage0_49[483]},
      {stage1_49[213]}
   );
   gpc1_1 gpc5128 (
      {stage0_49[484]},
      {stage1_49[214]}
   );
   gpc1_1 gpc5129 (
      {stage0_49[485]},
      {stage1_49[215]}
   );
   gpc1_1 gpc5130 (
      {stage0_49[486]},
      {stage1_49[216]}
   );
   gpc1_1 gpc5131 (
      {stage0_49[487]},
      {stage1_49[217]}
   );
   gpc1_1 gpc5132 (
      {stage0_49[488]},
      {stage1_49[218]}
   );
   gpc1_1 gpc5133 (
      {stage0_49[489]},
      {stage1_49[219]}
   );
   gpc1_1 gpc5134 (
      {stage0_49[490]},
      {stage1_49[220]}
   );
   gpc1_1 gpc5135 (
      {stage0_49[491]},
      {stage1_49[221]}
   );
   gpc1_1 gpc5136 (
      {stage0_49[492]},
      {stage1_49[222]}
   );
   gpc1_1 gpc5137 (
      {stage0_49[493]},
      {stage1_49[223]}
   );
   gpc1_1 gpc5138 (
      {stage0_49[494]},
      {stage1_49[224]}
   );
   gpc1_1 gpc5139 (
      {stage0_49[495]},
      {stage1_49[225]}
   );
   gpc1_1 gpc5140 (
      {stage0_49[496]},
      {stage1_49[226]}
   );
   gpc1_1 gpc5141 (
      {stage0_49[497]},
      {stage1_49[227]}
   );
   gpc1_1 gpc5142 (
      {stage0_49[498]},
      {stage1_49[228]}
   );
   gpc1_1 gpc5143 (
      {stage0_49[499]},
      {stage1_49[229]}
   );
   gpc1_1 gpc5144 (
      {stage0_49[500]},
      {stage1_49[230]}
   );
   gpc1_1 gpc5145 (
      {stage0_49[501]},
      {stage1_49[231]}
   );
   gpc1_1 gpc5146 (
      {stage0_49[502]},
      {stage1_49[232]}
   );
   gpc1_1 gpc5147 (
      {stage0_49[503]},
      {stage1_49[233]}
   );
   gpc1_1 gpc5148 (
      {stage0_49[504]},
      {stage1_49[234]}
   );
   gpc1_1 gpc5149 (
      {stage0_49[505]},
      {stage1_49[235]}
   );
   gpc1_1 gpc5150 (
      {stage0_49[506]},
      {stage1_49[236]}
   );
   gpc1_1 gpc5151 (
      {stage0_49[507]},
      {stage1_49[237]}
   );
   gpc1_1 gpc5152 (
      {stage0_49[508]},
      {stage1_49[238]}
   );
   gpc1_1 gpc5153 (
      {stage0_49[509]},
      {stage1_49[239]}
   );
   gpc1_1 gpc5154 (
      {stage0_49[510]},
      {stage1_49[240]}
   );
   gpc1_1 gpc5155 (
      {stage0_49[511]},
      {stage1_49[241]}
   );
   gpc1_1 gpc5156 (
      {stage0_50[474]},
      {stage1_50[179]}
   );
   gpc1_1 gpc5157 (
      {stage0_50[475]},
      {stage1_50[180]}
   );
   gpc1_1 gpc5158 (
      {stage0_50[476]},
      {stage1_50[181]}
   );
   gpc1_1 gpc5159 (
      {stage0_50[477]},
      {stage1_50[182]}
   );
   gpc1_1 gpc5160 (
      {stage0_50[478]},
      {stage1_50[183]}
   );
   gpc1_1 gpc5161 (
      {stage0_50[479]},
      {stage1_50[184]}
   );
   gpc1_1 gpc5162 (
      {stage0_50[480]},
      {stage1_50[185]}
   );
   gpc1_1 gpc5163 (
      {stage0_50[481]},
      {stage1_50[186]}
   );
   gpc1_1 gpc5164 (
      {stage0_50[482]},
      {stage1_50[187]}
   );
   gpc1_1 gpc5165 (
      {stage0_50[483]},
      {stage1_50[188]}
   );
   gpc1_1 gpc5166 (
      {stage0_50[484]},
      {stage1_50[189]}
   );
   gpc1_1 gpc5167 (
      {stage0_50[485]},
      {stage1_50[190]}
   );
   gpc1_1 gpc5168 (
      {stage0_50[486]},
      {stage1_50[191]}
   );
   gpc1_1 gpc5169 (
      {stage0_50[487]},
      {stage1_50[192]}
   );
   gpc1_1 gpc5170 (
      {stage0_50[488]},
      {stage1_50[193]}
   );
   gpc1_1 gpc5171 (
      {stage0_50[489]},
      {stage1_50[194]}
   );
   gpc1_1 gpc5172 (
      {stage0_50[490]},
      {stage1_50[195]}
   );
   gpc1_1 gpc5173 (
      {stage0_50[491]},
      {stage1_50[196]}
   );
   gpc1_1 gpc5174 (
      {stage0_50[492]},
      {stage1_50[197]}
   );
   gpc1_1 gpc5175 (
      {stage0_50[493]},
      {stage1_50[198]}
   );
   gpc1_1 gpc5176 (
      {stage0_50[494]},
      {stage1_50[199]}
   );
   gpc1_1 gpc5177 (
      {stage0_50[495]},
      {stage1_50[200]}
   );
   gpc1_1 gpc5178 (
      {stage0_50[496]},
      {stage1_50[201]}
   );
   gpc1_1 gpc5179 (
      {stage0_50[497]},
      {stage1_50[202]}
   );
   gpc1_1 gpc5180 (
      {stage0_50[498]},
      {stage1_50[203]}
   );
   gpc1_1 gpc5181 (
      {stage0_50[499]},
      {stage1_50[204]}
   );
   gpc1_1 gpc5182 (
      {stage0_50[500]},
      {stage1_50[205]}
   );
   gpc1_1 gpc5183 (
      {stage0_50[501]},
      {stage1_50[206]}
   );
   gpc1_1 gpc5184 (
      {stage0_50[502]},
      {stage1_50[207]}
   );
   gpc1_1 gpc5185 (
      {stage0_50[503]},
      {stage1_50[208]}
   );
   gpc1_1 gpc5186 (
      {stage0_50[504]},
      {stage1_50[209]}
   );
   gpc1_1 gpc5187 (
      {stage0_50[505]},
      {stage1_50[210]}
   );
   gpc1_1 gpc5188 (
      {stage0_50[506]},
      {stage1_50[211]}
   );
   gpc1_1 gpc5189 (
      {stage0_50[507]},
      {stage1_50[212]}
   );
   gpc1_1 gpc5190 (
      {stage0_50[508]},
      {stage1_50[213]}
   );
   gpc1_1 gpc5191 (
      {stage0_50[509]},
      {stage1_50[214]}
   );
   gpc1_1 gpc5192 (
      {stage0_50[510]},
      {stage1_50[215]}
   );
   gpc1_1 gpc5193 (
      {stage0_50[511]},
      {stage1_50[216]}
   );
   gpc1_1 gpc5194 (
      {stage0_51[501]},
      {stage1_51[216]}
   );
   gpc1_1 gpc5195 (
      {stage0_51[502]},
      {stage1_51[217]}
   );
   gpc1_1 gpc5196 (
      {stage0_51[503]},
      {stage1_51[218]}
   );
   gpc1_1 gpc5197 (
      {stage0_51[504]},
      {stage1_51[219]}
   );
   gpc1_1 gpc5198 (
      {stage0_51[505]},
      {stage1_51[220]}
   );
   gpc1_1 gpc5199 (
      {stage0_51[506]},
      {stage1_51[221]}
   );
   gpc1_1 gpc5200 (
      {stage0_51[507]},
      {stage1_51[222]}
   );
   gpc1_1 gpc5201 (
      {stage0_51[508]},
      {stage1_51[223]}
   );
   gpc1_1 gpc5202 (
      {stage0_51[509]},
      {stage1_51[224]}
   );
   gpc1_1 gpc5203 (
      {stage0_51[510]},
      {stage1_51[225]}
   );
   gpc1_1 gpc5204 (
      {stage0_51[511]},
      {stage1_51[226]}
   );
   gpc1_1 gpc5205 (
      {stage0_52[410]},
      {stage1_52[202]}
   );
   gpc1_1 gpc5206 (
      {stage0_52[411]},
      {stage1_52[203]}
   );
   gpc1_1 gpc5207 (
      {stage0_52[412]},
      {stage1_52[204]}
   );
   gpc1_1 gpc5208 (
      {stage0_52[413]},
      {stage1_52[205]}
   );
   gpc1_1 gpc5209 (
      {stage0_52[414]},
      {stage1_52[206]}
   );
   gpc1_1 gpc5210 (
      {stage0_52[415]},
      {stage1_52[207]}
   );
   gpc1_1 gpc5211 (
      {stage0_52[416]},
      {stage1_52[208]}
   );
   gpc1_1 gpc5212 (
      {stage0_52[417]},
      {stage1_52[209]}
   );
   gpc1_1 gpc5213 (
      {stage0_52[418]},
      {stage1_52[210]}
   );
   gpc1_1 gpc5214 (
      {stage0_52[419]},
      {stage1_52[211]}
   );
   gpc1_1 gpc5215 (
      {stage0_52[420]},
      {stage1_52[212]}
   );
   gpc1_1 gpc5216 (
      {stage0_52[421]},
      {stage1_52[213]}
   );
   gpc1_1 gpc5217 (
      {stage0_52[422]},
      {stage1_52[214]}
   );
   gpc1_1 gpc5218 (
      {stage0_52[423]},
      {stage1_52[215]}
   );
   gpc1_1 gpc5219 (
      {stage0_52[424]},
      {stage1_52[216]}
   );
   gpc1_1 gpc5220 (
      {stage0_52[425]},
      {stage1_52[217]}
   );
   gpc1_1 gpc5221 (
      {stage0_52[426]},
      {stage1_52[218]}
   );
   gpc1_1 gpc5222 (
      {stage0_52[427]},
      {stage1_52[219]}
   );
   gpc1_1 gpc5223 (
      {stage0_52[428]},
      {stage1_52[220]}
   );
   gpc1_1 gpc5224 (
      {stage0_52[429]},
      {stage1_52[221]}
   );
   gpc1_1 gpc5225 (
      {stage0_52[430]},
      {stage1_52[222]}
   );
   gpc1_1 gpc5226 (
      {stage0_52[431]},
      {stage1_52[223]}
   );
   gpc1_1 gpc5227 (
      {stage0_52[432]},
      {stage1_52[224]}
   );
   gpc1_1 gpc5228 (
      {stage0_52[433]},
      {stage1_52[225]}
   );
   gpc1_1 gpc5229 (
      {stage0_52[434]},
      {stage1_52[226]}
   );
   gpc1_1 gpc5230 (
      {stage0_52[435]},
      {stage1_52[227]}
   );
   gpc1_1 gpc5231 (
      {stage0_52[436]},
      {stage1_52[228]}
   );
   gpc1_1 gpc5232 (
      {stage0_52[437]},
      {stage1_52[229]}
   );
   gpc1_1 gpc5233 (
      {stage0_52[438]},
      {stage1_52[230]}
   );
   gpc1_1 gpc5234 (
      {stage0_52[439]},
      {stage1_52[231]}
   );
   gpc1_1 gpc5235 (
      {stage0_52[440]},
      {stage1_52[232]}
   );
   gpc1_1 gpc5236 (
      {stage0_52[441]},
      {stage1_52[233]}
   );
   gpc1_1 gpc5237 (
      {stage0_52[442]},
      {stage1_52[234]}
   );
   gpc1_1 gpc5238 (
      {stage0_52[443]},
      {stage1_52[235]}
   );
   gpc1_1 gpc5239 (
      {stage0_52[444]},
      {stage1_52[236]}
   );
   gpc1_1 gpc5240 (
      {stage0_52[445]},
      {stage1_52[237]}
   );
   gpc1_1 gpc5241 (
      {stage0_52[446]},
      {stage1_52[238]}
   );
   gpc1_1 gpc5242 (
      {stage0_52[447]},
      {stage1_52[239]}
   );
   gpc1_1 gpc5243 (
      {stage0_52[448]},
      {stage1_52[240]}
   );
   gpc1_1 gpc5244 (
      {stage0_52[449]},
      {stage1_52[241]}
   );
   gpc1_1 gpc5245 (
      {stage0_52[450]},
      {stage1_52[242]}
   );
   gpc1_1 gpc5246 (
      {stage0_52[451]},
      {stage1_52[243]}
   );
   gpc1_1 gpc5247 (
      {stage0_52[452]},
      {stage1_52[244]}
   );
   gpc1_1 gpc5248 (
      {stage0_52[453]},
      {stage1_52[245]}
   );
   gpc1_1 gpc5249 (
      {stage0_52[454]},
      {stage1_52[246]}
   );
   gpc1_1 gpc5250 (
      {stage0_52[455]},
      {stage1_52[247]}
   );
   gpc1_1 gpc5251 (
      {stage0_52[456]},
      {stage1_52[248]}
   );
   gpc1_1 gpc5252 (
      {stage0_52[457]},
      {stage1_52[249]}
   );
   gpc1_1 gpc5253 (
      {stage0_52[458]},
      {stage1_52[250]}
   );
   gpc1_1 gpc5254 (
      {stage0_52[459]},
      {stage1_52[251]}
   );
   gpc1_1 gpc5255 (
      {stage0_52[460]},
      {stage1_52[252]}
   );
   gpc1_1 gpc5256 (
      {stage0_52[461]},
      {stage1_52[253]}
   );
   gpc1_1 gpc5257 (
      {stage0_52[462]},
      {stage1_52[254]}
   );
   gpc1_1 gpc5258 (
      {stage0_52[463]},
      {stage1_52[255]}
   );
   gpc1_1 gpc5259 (
      {stage0_52[464]},
      {stage1_52[256]}
   );
   gpc1_1 gpc5260 (
      {stage0_52[465]},
      {stage1_52[257]}
   );
   gpc1_1 gpc5261 (
      {stage0_52[466]},
      {stage1_52[258]}
   );
   gpc1_1 gpc5262 (
      {stage0_52[467]},
      {stage1_52[259]}
   );
   gpc1_1 gpc5263 (
      {stage0_52[468]},
      {stage1_52[260]}
   );
   gpc1_1 gpc5264 (
      {stage0_52[469]},
      {stage1_52[261]}
   );
   gpc1_1 gpc5265 (
      {stage0_52[470]},
      {stage1_52[262]}
   );
   gpc1_1 gpc5266 (
      {stage0_52[471]},
      {stage1_52[263]}
   );
   gpc1_1 gpc5267 (
      {stage0_52[472]},
      {stage1_52[264]}
   );
   gpc1_1 gpc5268 (
      {stage0_52[473]},
      {stage1_52[265]}
   );
   gpc1_1 gpc5269 (
      {stage0_52[474]},
      {stage1_52[266]}
   );
   gpc1_1 gpc5270 (
      {stage0_52[475]},
      {stage1_52[267]}
   );
   gpc1_1 gpc5271 (
      {stage0_52[476]},
      {stage1_52[268]}
   );
   gpc1_1 gpc5272 (
      {stage0_52[477]},
      {stage1_52[269]}
   );
   gpc1_1 gpc5273 (
      {stage0_52[478]},
      {stage1_52[270]}
   );
   gpc1_1 gpc5274 (
      {stage0_52[479]},
      {stage1_52[271]}
   );
   gpc1_1 gpc5275 (
      {stage0_52[480]},
      {stage1_52[272]}
   );
   gpc1_1 gpc5276 (
      {stage0_52[481]},
      {stage1_52[273]}
   );
   gpc1_1 gpc5277 (
      {stage0_52[482]},
      {stage1_52[274]}
   );
   gpc1_1 gpc5278 (
      {stage0_52[483]},
      {stage1_52[275]}
   );
   gpc1_1 gpc5279 (
      {stage0_52[484]},
      {stage1_52[276]}
   );
   gpc1_1 gpc5280 (
      {stage0_52[485]},
      {stage1_52[277]}
   );
   gpc1_1 gpc5281 (
      {stage0_52[486]},
      {stage1_52[278]}
   );
   gpc1_1 gpc5282 (
      {stage0_52[487]},
      {stage1_52[279]}
   );
   gpc1_1 gpc5283 (
      {stage0_52[488]},
      {stage1_52[280]}
   );
   gpc1_1 gpc5284 (
      {stage0_52[489]},
      {stage1_52[281]}
   );
   gpc1_1 gpc5285 (
      {stage0_52[490]},
      {stage1_52[282]}
   );
   gpc1_1 gpc5286 (
      {stage0_52[491]},
      {stage1_52[283]}
   );
   gpc1_1 gpc5287 (
      {stage0_52[492]},
      {stage1_52[284]}
   );
   gpc1_1 gpc5288 (
      {stage0_52[493]},
      {stage1_52[285]}
   );
   gpc1_1 gpc5289 (
      {stage0_52[494]},
      {stage1_52[286]}
   );
   gpc1_1 gpc5290 (
      {stage0_52[495]},
      {stage1_52[287]}
   );
   gpc1_1 gpc5291 (
      {stage0_52[496]},
      {stage1_52[288]}
   );
   gpc1_1 gpc5292 (
      {stage0_52[497]},
      {stage1_52[289]}
   );
   gpc1_1 gpc5293 (
      {stage0_52[498]},
      {stage1_52[290]}
   );
   gpc1_1 gpc5294 (
      {stage0_52[499]},
      {stage1_52[291]}
   );
   gpc1_1 gpc5295 (
      {stage0_52[500]},
      {stage1_52[292]}
   );
   gpc1_1 gpc5296 (
      {stage0_52[501]},
      {stage1_52[293]}
   );
   gpc1_1 gpc5297 (
      {stage0_52[502]},
      {stage1_52[294]}
   );
   gpc1_1 gpc5298 (
      {stage0_52[503]},
      {stage1_52[295]}
   );
   gpc1_1 gpc5299 (
      {stage0_52[504]},
      {stage1_52[296]}
   );
   gpc1_1 gpc5300 (
      {stage0_52[505]},
      {stage1_52[297]}
   );
   gpc1_1 gpc5301 (
      {stage0_52[506]},
      {stage1_52[298]}
   );
   gpc1_1 gpc5302 (
      {stage0_52[507]},
      {stage1_52[299]}
   );
   gpc1_1 gpc5303 (
      {stage0_52[508]},
      {stage1_52[300]}
   );
   gpc1_1 gpc5304 (
      {stage0_52[509]},
      {stage1_52[301]}
   );
   gpc1_1 gpc5305 (
      {stage0_52[510]},
      {stage1_52[302]}
   );
   gpc1_1 gpc5306 (
      {stage0_52[511]},
      {stage1_52[303]}
   );
   gpc1_1 gpc5307 (
      {stage0_53[497]},
      {stage1_53[172]}
   );
   gpc1_1 gpc5308 (
      {stage0_53[498]},
      {stage1_53[173]}
   );
   gpc1_1 gpc5309 (
      {stage0_53[499]},
      {stage1_53[174]}
   );
   gpc1_1 gpc5310 (
      {stage0_53[500]},
      {stage1_53[175]}
   );
   gpc1_1 gpc5311 (
      {stage0_53[501]},
      {stage1_53[176]}
   );
   gpc1_1 gpc5312 (
      {stage0_53[502]},
      {stage1_53[177]}
   );
   gpc1_1 gpc5313 (
      {stage0_53[503]},
      {stage1_53[178]}
   );
   gpc1_1 gpc5314 (
      {stage0_53[504]},
      {stage1_53[179]}
   );
   gpc1_1 gpc5315 (
      {stage0_53[505]},
      {stage1_53[180]}
   );
   gpc1_1 gpc5316 (
      {stage0_53[506]},
      {stage1_53[181]}
   );
   gpc1_1 gpc5317 (
      {stage0_53[507]},
      {stage1_53[182]}
   );
   gpc1_1 gpc5318 (
      {stage0_53[508]},
      {stage1_53[183]}
   );
   gpc1_1 gpc5319 (
      {stage0_53[509]},
      {stage1_53[184]}
   );
   gpc1_1 gpc5320 (
      {stage0_53[510]},
      {stage1_53[185]}
   );
   gpc1_1 gpc5321 (
      {stage0_53[511]},
      {stage1_53[186]}
   );
   gpc1_1 gpc5322 (
      {stage0_54[441]},
      {stage1_54[192]}
   );
   gpc1_1 gpc5323 (
      {stage0_54[442]},
      {stage1_54[193]}
   );
   gpc1_1 gpc5324 (
      {stage0_54[443]},
      {stage1_54[194]}
   );
   gpc1_1 gpc5325 (
      {stage0_54[444]},
      {stage1_54[195]}
   );
   gpc1_1 gpc5326 (
      {stage0_54[445]},
      {stage1_54[196]}
   );
   gpc1_1 gpc5327 (
      {stage0_54[446]},
      {stage1_54[197]}
   );
   gpc1_1 gpc5328 (
      {stage0_54[447]},
      {stage1_54[198]}
   );
   gpc1_1 gpc5329 (
      {stage0_54[448]},
      {stage1_54[199]}
   );
   gpc1_1 gpc5330 (
      {stage0_54[449]},
      {stage1_54[200]}
   );
   gpc1_1 gpc5331 (
      {stage0_54[450]},
      {stage1_54[201]}
   );
   gpc1_1 gpc5332 (
      {stage0_54[451]},
      {stage1_54[202]}
   );
   gpc1_1 gpc5333 (
      {stage0_54[452]},
      {stage1_54[203]}
   );
   gpc1_1 gpc5334 (
      {stage0_54[453]},
      {stage1_54[204]}
   );
   gpc1_1 gpc5335 (
      {stage0_54[454]},
      {stage1_54[205]}
   );
   gpc1_1 gpc5336 (
      {stage0_54[455]},
      {stage1_54[206]}
   );
   gpc1_1 gpc5337 (
      {stage0_54[456]},
      {stage1_54[207]}
   );
   gpc1_1 gpc5338 (
      {stage0_54[457]},
      {stage1_54[208]}
   );
   gpc1_1 gpc5339 (
      {stage0_54[458]},
      {stage1_54[209]}
   );
   gpc1_1 gpc5340 (
      {stage0_54[459]},
      {stage1_54[210]}
   );
   gpc1_1 gpc5341 (
      {stage0_54[460]},
      {stage1_54[211]}
   );
   gpc1_1 gpc5342 (
      {stage0_54[461]},
      {stage1_54[212]}
   );
   gpc1_1 gpc5343 (
      {stage0_54[462]},
      {stage1_54[213]}
   );
   gpc1_1 gpc5344 (
      {stage0_54[463]},
      {stage1_54[214]}
   );
   gpc1_1 gpc5345 (
      {stage0_54[464]},
      {stage1_54[215]}
   );
   gpc1_1 gpc5346 (
      {stage0_54[465]},
      {stage1_54[216]}
   );
   gpc1_1 gpc5347 (
      {stage0_54[466]},
      {stage1_54[217]}
   );
   gpc1_1 gpc5348 (
      {stage0_54[467]},
      {stage1_54[218]}
   );
   gpc1_1 gpc5349 (
      {stage0_54[468]},
      {stage1_54[219]}
   );
   gpc1_1 gpc5350 (
      {stage0_54[469]},
      {stage1_54[220]}
   );
   gpc1_1 gpc5351 (
      {stage0_54[470]},
      {stage1_54[221]}
   );
   gpc1_1 gpc5352 (
      {stage0_54[471]},
      {stage1_54[222]}
   );
   gpc1_1 gpc5353 (
      {stage0_54[472]},
      {stage1_54[223]}
   );
   gpc1_1 gpc5354 (
      {stage0_54[473]},
      {stage1_54[224]}
   );
   gpc1_1 gpc5355 (
      {stage0_54[474]},
      {stage1_54[225]}
   );
   gpc1_1 gpc5356 (
      {stage0_54[475]},
      {stage1_54[226]}
   );
   gpc1_1 gpc5357 (
      {stage0_54[476]},
      {stage1_54[227]}
   );
   gpc1_1 gpc5358 (
      {stage0_54[477]},
      {stage1_54[228]}
   );
   gpc1_1 gpc5359 (
      {stage0_54[478]},
      {stage1_54[229]}
   );
   gpc1_1 gpc5360 (
      {stage0_54[479]},
      {stage1_54[230]}
   );
   gpc1_1 gpc5361 (
      {stage0_54[480]},
      {stage1_54[231]}
   );
   gpc1_1 gpc5362 (
      {stage0_54[481]},
      {stage1_54[232]}
   );
   gpc1_1 gpc5363 (
      {stage0_54[482]},
      {stage1_54[233]}
   );
   gpc1_1 gpc5364 (
      {stage0_54[483]},
      {stage1_54[234]}
   );
   gpc1_1 gpc5365 (
      {stage0_54[484]},
      {stage1_54[235]}
   );
   gpc1_1 gpc5366 (
      {stage0_54[485]},
      {stage1_54[236]}
   );
   gpc1_1 gpc5367 (
      {stage0_54[486]},
      {stage1_54[237]}
   );
   gpc1_1 gpc5368 (
      {stage0_54[487]},
      {stage1_54[238]}
   );
   gpc1_1 gpc5369 (
      {stage0_54[488]},
      {stage1_54[239]}
   );
   gpc1_1 gpc5370 (
      {stage0_54[489]},
      {stage1_54[240]}
   );
   gpc1_1 gpc5371 (
      {stage0_54[490]},
      {stage1_54[241]}
   );
   gpc1_1 gpc5372 (
      {stage0_54[491]},
      {stage1_54[242]}
   );
   gpc1_1 gpc5373 (
      {stage0_54[492]},
      {stage1_54[243]}
   );
   gpc1_1 gpc5374 (
      {stage0_54[493]},
      {stage1_54[244]}
   );
   gpc1_1 gpc5375 (
      {stage0_54[494]},
      {stage1_54[245]}
   );
   gpc1_1 gpc5376 (
      {stage0_54[495]},
      {stage1_54[246]}
   );
   gpc1_1 gpc5377 (
      {stage0_54[496]},
      {stage1_54[247]}
   );
   gpc1_1 gpc5378 (
      {stage0_54[497]},
      {stage1_54[248]}
   );
   gpc1_1 gpc5379 (
      {stage0_54[498]},
      {stage1_54[249]}
   );
   gpc1_1 gpc5380 (
      {stage0_54[499]},
      {stage1_54[250]}
   );
   gpc1_1 gpc5381 (
      {stage0_54[500]},
      {stage1_54[251]}
   );
   gpc1_1 gpc5382 (
      {stage0_54[501]},
      {stage1_54[252]}
   );
   gpc1_1 gpc5383 (
      {stage0_54[502]},
      {stage1_54[253]}
   );
   gpc1_1 gpc5384 (
      {stage0_54[503]},
      {stage1_54[254]}
   );
   gpc1_1 gpc5385 (
      {stage0_54[504]},
      {stage1_54[255]}
   );
   gpc1_1 gpc5386 (
      {stage0_54[505]},
      {stage1_54[256]}
   );
   gpc1_1 gpc5387 (
      {stage0_54[506]},
      {stage1_54[257]}
   );
   gpc1_1 gpc5388 (
      {stage0_54[507]},
      {stage1_54[258]}
   );
   gpc1_1 gpc5389 (
      {stage0_54[508]},
      {stage1_54[259]}
   );
   gpc1_1 gpc5390 (
      {stage0_54[509]},
      {stage1_54[260]}
   );
   gpc1_1 gpc5391 (
      {stage0_54[510]},
      {stage1_54[261]}
   );
   gpc1_1 gpc5392 (
      {stage0_54[511]},
      {stage1_54[262]}
   );
   gpc1_1 gpc5393 (
      {stage0_55[508]},
      {stage1_55[222]}
   );
   gpc1_1 gpc5394 (
      {stage0_55[509]},
      {stage1_55[223]}
   );
   gpc1_1 gpc5395 (
      {stage0_55[510]},
      {stage1_55[224]}
   );
   gpc1_1 gpc5396 (
      {stage0_55[511]},
      {stage1_55[225]}
   );
   gpc1_1 gpc5397 (
      {stage0_56[444]},
      {stage1_56[189]}
   );
   gpc1_1 gpc5398 (
      {stage0_56[445]},
      {stage1_56[190]}
   );
   gpc1_1 gpc5399 (
      {stage0_56[446]},
      {stage1_56[191]}
   );
   gpc1_1 gpc5400 (
      {stage0_56[447]},
      {stage1_56[192]}
   );
   gpc1_1 gpc5401 (
      {stage0_56[448]},
      {stage1_56[193]}
   );
   gpc1_1 gpc5402 (
      {stage0_56[449]},
      {stage1_56[194]}
   );
   gpc1_1 gpc5403 (
      {stage0_56[450]},
      {stage1_56[195]}
   );
   gpc1_1 gpc5404 (
      {stage0_56[451]},
      {stage1_56[196]}
   );
   gpc1_1 gpc5405 (
      {stage0_56[452]},
      {stage1_56[197]}
   );
   gpc1_1 gpc5406 (
      {stage0_56[453]},
      {stage1_56[198]}
   );
   gpc1_1 gpc5407 (
      {stage0_56[454]},
      {stage1_56[199]}
   );
   gpc1_1 gpc5408 (
      {stage0_56[455]},
      {stage1_56[200]}
   );
   gpc1_1 gpc5409 (
      {stage0_56[456]},
      {stage1_56[201]}
   );
   gpc1_1 gpc5410 (
      {stage0_56[457]},
      {stage1_56[202]}
   );
   gpc1_1 gpc5411 (
      {stage0_56[458]},
      {stage1_56[203]}
   );
   gpc1_1 gpc5412 (
      {stage0_56[459]},
      {stage1_56[204]}
   );
   gpc1_1 gpc5413 (
      {stage0_56[460]},
      {stage1_56[205]}
   );
   gpc1_1 gpc5414 (
      {stage0_56[461]},
      {stage1_56[206]}
   );
   gpc1_1 gpc5415 (
      {stage0_56[462]},
      {stage1_56[207]}
   );
   gpc1_1 gpc5416 (
      {stage0_56[463]},
      {stage1_56[208]}
   );
   gpc1_1 gpc5417 (
      {stage0_56[464]},
      {stage1_56[209]}
   );
   gpc1_1 gpc5418 (
      {stage0_56[465]},
      {stage1_56[210]}
   );
   gpc1_1 gpc5419 (
      {stage0_56[466]},
      {stage1_56[211]}
   );
   gpc1_1 gpc5420 (
      {stage0_56[467]},
      {stage1_56[212]}
   );
   gpc1_1 gpc5421 (
      {stage0_56[468]},
      {stage1_56[213]}
   );
   gpc1_1 gpc5422 (
      {stage0_56[469]},
      {stage1_56[214]}
   );
   gpc1_1 gpc5423 (
      {stage0_56[470]},
      {stage1_56[215]}
   );
   gpc1_1 gpc5424 (
      {stage0_56[471]},
      {stage1_56[216]}
   );
   gpc1_1 gpc5425 (
      {stage0_56[472]},
      {stage1_56[217]}
   );
   gpc1_1 gpc5426 (
      {stage0_56[473]},
      {stage1_56[218]}
   );
   gpc1_1 gpc5427 (
      {stage0_56[474]},
      {stage1_56[219]}
   );
   gpc1_1 gpc5428 (
      {stage0_56[475]},
      {stage1_56[220]}
   );
   gpc1_1 gpc5429 (
      {stage0_56[476]},
      {stage1_56[221]}
   );
   gpc1_1 gpc5430 (
      {stage0_56[477]},
      {stage1_56[222]}
   );
   gpc1_1 gpc5431 (
      {stage0_56[478]},
      {stage1_56[223]}
   );
   gpc1_1 gpc5432 (
      {stage0_56[479]},
      {stage1_56[224]}
   );
   gpc1_1 gpc5433 (
      {stage0_56[480]},
      {stage1_56[225]}
   );
   gpc1_1 gpc5434 (
      {stage0_56[481]},
      {stage1_56[226]}
   );
   gpc1_1 gpc5435 (
      {stage0_56[482]},
      {stage1_56[227]}
   );
   gpc1_1 gpc5436 (
      {stage0_56[483]},
      {stage1_56[228]}
   );
   gpc1_1 gpc5437 (
      {stage0_56[484]},
      {stage1_56[229]}
   );
   gpc1_1 gpc5438 (
      {stage0_56[485]},
      {stage1_56[230]}
   );
   gpc1_1 gpc5439 (
      {stage0_56[486]},
      {stage1_56[231]}
   );
   gpc1_1 gpc5440 (
      {stage0_56[487]},
      {stage1_56[232]}
   );
   gpc1_1 gpc5441 (
      {stage0_56[488]},
      {stage1_56[233]}
   );
   gpc1_1 gpc5442 (
      {stage0_56[489]},
      {stage1_56[234]}
   );
   gpc1_1 gpc5443 (
      {stage0_56[490]},
      {stage1_56[235]}
   );
   gpc1_1 gpc5444 (
      {stage0_56[491]},
      {stage1_56[236]}
   );
   gpc1_1 gpc5445 (
      {stage0_56[492]},
      {stage1_56[237]}
   );
   gpc1_1 gpc5446 (
      {stage0_56[493]},
      {stage1_56[238]}
   );
   gpc1_1 gpc5447 (
      {stage0_56[494]},
      {stage1_56[239]}
   );
   gpc1_1 gpc5448 (
      {stage0_56[495]},
      {stage1_56[240]}
   );
   gpc1_1 gpc5449 (
      {stage0_56[496]},
      {stage1_56[241]}
   );
   gpc1_1 gpc5450 (
      {stage0_56[497]},
      {stage1_56[242]}
   );
   gpc1_1 gpc5451 (
      {stage0_56[498]},
      {stage1_56[243]}
   );
   gpc1_1 gpc5452 (
      {stage0_56[499]},
      {stage1_56[244]}
   );
   gpc1_1 gpc5453 (
      {stage0_56[500]},
      {stage1_56[245]}
   );
   gpc1_1 gpc5454 (
      {stage0_56[501]},
      {stage1_56[246]}
   );
   gpc1_1 gpc5455 (
      {stage0_56[502]},
      {stage1_56[247]}
   );
   gpc1_1 gpc5456 (
      {stage0_56[503]},
      {stage1_56[248]}
   );
   gpc1_1 gpc5457 (
      {stage0_56[504]},
      {stage1_56[249]}
   );
   gpc1_1 gpc5458 (
      {stage0_56[505]},
      {stage1_56[250]}
   );
   gpc1_1 gpc5459 (
      {stage0_56[506]},
      {stage1_56[251]}
   );
   gpc1_1 gpc5460 (
      {stage0_56[507]},
      {stage1_56[252]}
   );
   gpc1_1 gpc5461 (
      {stage0_56[508]},
      {stage1_56[253]}
   );
   gpc1_1 gpc5462 (
      {stage0_56[509]},
      {stage1_56[254]}
   );
   gpc1_1 gpc5463 (
      {stage0_56[510]},
      {stage1_56[255]}
   );
   gpc1_1 gpc5464 (
      {stage0_56[511]},
      {stage1_56[256]}
   );
   gpc1_1 gpc5465 (
      {stage0_57[510]},
      {stage1_57[178]}
   );
   gpc1_1 gpc5466 (
      {stage0_57[511]},
      {stage1_57[179]}
   );
   gpc1_1 gpc5467 (
      {stage0_58[493]},
      {stage1_58[224]}
   );
   gpc1_1 gpc5468 (
      {stage0_58[494]},
      {stage1_58[225]}
   );
   gpc1_1 gpc5469 (
      {stage0_58[495]},
      {stage1_58[226]}
   );
   gpc1_1 gpc5470 (
      {stage0_58[496]},
      {stage1_58[227]}
   );
   gpc1_1 gpc5471 (
      {stage0_58[497]},
      {stage1_58[228]}
   );
   gpc1_1 gpc5472 (
      {stage0_58[498]},
      {stage1_58[229]}
   );
   gpc1_1 gpc5473 (
      {stage0_58[499]},
      {stage1_58[230]}
   );
   gpc1_1 gpc5474 (
      {stage0_58[500]},
      {stage1_58[231]}
   );
   gpc1_1 gpc5475 (
      {stage0_58[501]},
      {stage1_58[232]}
   );
   gpc1_1 gpc5476 (
      {stage0_58[502]},
      {stage1_58[233]}
   );
   gpc1_1 gpc5477 (
      {stage0_58[503]},
      {stage1_58[234]}
   );
   gpc1_1 gpc5478 (
      {stage0_58[504]},
      {stage1_58[235]}
   );
   gpc1_1 gpc5479 (
      {stage0_58[505]},
      {stage1_58[236]}
   );
   gpc1_1 gpc5480 (
      {stage0_58[506]},
      {stage1_58[237]}
   );
   gpc1_1 gpc5481 (
      {stage0_58[507]},
      {stage1_58[238]}
   );
   gpc1_1 gpc5482 (
      {stage0_58[508]},
      {stage1_58[239]}
   );
   gpc1_1 gpc5483 (
      {stage0_58[509]},
      {stage1_58[240]}
   );
   gpc1_1 gpc5484 (
      {stage0_58[510]},
      {stage1_58[241]}
   );
   gpc1_1 gpc5485 (
      {stage0_58[511]},
      {stage1_58[242]}
   );
   gpc1_1 gpc5486 (
      {stage0_59[412]},
      {stage1_59[194]}
   );
   gpc1_1 gpc5487 (
      {stage0_59[413]},
      {stage1_59[195]}
   );
   gpc1_1 gpc5488 (
      {stage0_59[414]},
      {stage1_59[196]}
   );
   gpc1_1 gpc5489 (
      {stage0_59[415]},
      {stage1_59[197]}
   );
   gpc1_1 gpc5490 (
      {stage0_59[416]},
      {stage1_59[198]}
   );
   gpc1_1 gpc5491 (
      {stage0_59[417]},
      {stage1_59[199]}
   );
   gpc1_1 gpc5492 (
      {stage0_59[418]},
      {stage1_59[200]}
   );
   gpc1_1 gpc5493 (
      {stage0_59[419]},
      {stage1_59[201]}
   );
   gpc1_1 gpc5494 (
      {stage0_59[420]},
      {stage1_59[202]}
   );
   gpc1_1 gpc5495 (
      {stage0_59[421]},
      {stage1_59[203]}
   );
   gpc1_1 gpc5496 (
      {stage0_59[422]},
      {stage1_59[204]}
   );
   gpc1_1 gpc5497 (
      {stage0_59[423]},
      {stage1_59[205]}
   );
   gpc1_1 gpc5498 (
      {stage0_59[424]},
      {stage1_59[206]}
   );
   gpc1_1 gpc5499 (
      {stage0_59[425]},
      {stage1_59[207]}
   );
   gpc1_1 gpc5500 (
      {stage0_59[426]},
      {stage1_59[208]}
   );
   gpc1_1 gpc5501 (
      {stage0_59[427]},
      {stage1_59[209]}
   );
   gpc1_1 gpc5502 (
      {stage0_59[428]},
      {stage1_59[210]}
   );
   gpc1_1 gpc5503 (
      {stage0_59[429]},
      {stage1_59[211]}
   );
   gpc1_1 gpc5504 (
      {stage0_59[430]},
      {stage1_59[212]}
   );
   gpc1_1 gpc5505 (
      {stage0_59[431]},
      {stage1_59[213]}
   );
   gpc1_1 gpc5506 (
      {stage0_59[432]},
      {stage1_59[214]}
   );
   gpc1_1 gpc5507 (
      {stage0_59[433]},
      {stage1_59[215]}
   );
   gpc1_1 gpc5508 (
      {stage0_59[434]},
      {stage1_59[216]}
   );
   gpc1_1 gpc5509 (
      {stage0_59[435]},
      {stage1_59[217]}
   );
   gpc1_1 gpc5510 (
      {stage0_59[436]},
      {stage1_59[218]}
   );
   gpc1_1 gpc5511 (
      {stage0_59[437]},
      {stage1_59[219]}
   );
   gpc1_1 gpc5512 (
      {stage0_59[438]},
      {stage1_59[220]}
   );
   gpc1_1 gpc5513 (
      {stage0_59[439]},
      {stage1_59[221]}
   );
   gpc1_1 gpc5514 (
      {stage0_59[440]},
      {stage1_59[222]}
   );
   gpc1_1 gpc5515 (
      {stage0_59[441]},
      {stage1_59[223]}
   );
   gpc1_1 gpc5516 (
      {stage0_59[442]},
      {stage1_59[224]}
   );
   gpc1_1 gpc5517 (
      {stage0_59[443]},
      {stage1_59[225]}
   );
   gpc1_1 gpc5518 (
      {stage0_59[444]},
      {stage1_59[226]}
   );
   gpc1_1 gpc5519 (
      {stage0_59[445]},
      {stage1_59[227]}
   );
   gpc1_1 gpc5520 (
      {stage0_59[446]},
      {stage1_59[228]}
   );
   gpc1_1 gpc5521 (
      {stage0_59[447]},
      {stage1_59[229]}
   );
   gpc1_1 gpc5522 (
      {stage0_59[448]},
      {stage1_59[230]}
   );
   gpc1_1 gpc5523 (
      {stage0_59[449]},
      {stage1_59[231]}
   );
   gpc1_1 gpc5524 (
      {stage0_59[450]},
      {stage1_59[232]}
   );
   gpc1_1 gpc5525 (
      {stage0_59[451]},
      {stage1_59[233]}
   );
   gpc1_1 gpc5526 (
      {stage0_59[452]},
      {stage1_59[234]}
   );
   gpc1_1 gpc5527 (
      {stage0_59[453]},
      {stage1_59[235]}
   );
   gpc1_1 gpc5528 (
      {stage0_59[454]},
      {stage1_59[236]}
   );
   gpc1_1 gpc5529 (
      {stage0_59[455]},
      {stage1_59[237]}
   );
   gpc1_1 gpc5530 (
      {stage0_59[456]},
      {stage1_59[238]}
   );
   gpc1_1 gpc5531 (
      {stage0_59[457]},
      {stage1_59[239]}
   );
   gpc1_1 gpc5532 (
      {stage0_59[458]},
      {stage1_59[240]}
   );
   gpc1_1 gpc5533 (
      {stage0_59[459]},
      {stage1_59[241]}
   );
   gpc1_1 gpc5534 (
      {stage0_59[460]},
      {stage1_59[242]}
   );
   gpc1_1 gpc5535 (
      {stage0_59[461]},
      {stage1_59[243]}
   );
   gpc1_1 gpc5536 (
      {stage0_59[462]},
      {stage1_59[244]}
   );
   gpc1_1 gpc5537 (
      {stage0_59[463]},
      {stage1_59[245]}
   );
   gpc1_1 gpc5538 (
      {stage0_59[464]},
      {stage1_59[246]}
   );
   gpc1_1 gpc5539 (
      {stage0_59[465]},
      {stage1_59[247]}
   );
   gpc1_1 gpc5540 (
      {stage0_59[466]},
      {stage1_59[248]}
   );
   gpc1_1 gpc5541 (
      {stage0_59[467]},
      {stage1_59[249]}
   );
   gpc1_1 gpc5542 (
      {stage0_59[468]},
      {stage1_59[250]}
   );
   gpc1_1 gpc5543 (
      {stage0_59[469]},
      {stage1_59[251]}
   );
   gpc1_1 gpc5544 (
      {stage0_59[470]},
      {stage1_59[252]}
   );
   gpc1_1 gpc5545 (
      {stage0_59[471]},
      {stage1_59[253]}
   );
   gpc1_1 gpc5546 (
      {stage0_59[472]},
      {stage1_59[254]}
   );
   gpc1_1 gpc5547 (
      {stage0_59[473]},
      {stage1_59[255]}
   );
   gpc1_1 gpc5548 (
      {stage0_59[474]},
      {stage1_59[256]}
   );
   gpc1_1 gpc5549 (
      {stage0_59[475]},
      {stage1_59[257]}
   );
   gpc1_1 gpc5550 (
      {stage0_59[476]},
      {stage1_59[258]}
   );
   gpc1_1 gpc5551 (
      {stage0_59[477]},
      {stage1_59[259]}
   );
   gpc1_1 gpc5552 (
      {stage0_59[478]},
      {stage1_59[260]}
   );
   gpc1_1 gpc5553 (
      {stage0_59[479]},
      {stage1_59[261]}
   );
   gpc1_1 gpc5554 (
      {stage0_59[480]},
      {stage1_59[262]}
   );
   gpc1_1 gpc5555 (
      {stage0_59[481]},
      {stage1_59[263]}
   );
   gpc1_1 gpc5556 (
      {stage0_59[482]},
      {stage1_59[264]}
   );
   gpc1_1 gpc5557 (
      {stage0_59[483]},
      {stage1_59[265]}
   );
   gpc1_1 gpc5558 (
      {stage0_59[484]},
      {stage1_59[266]}
   );
   gpc1_1 gpc5559 (
      {stage0_59[485]},
      {stage1_59[267]}
   );
   gpc1_1 gpc5560 (
      {stage0_59[486]},
      {stage1_59[268]}
   );
   gpc1_1 gpc5561 (
      {stage0_59[487]},
      {stage1_59[269]}
   );
   gpc1_1 gpc5562 (
      {stage0_59[488]},
      {stage1_59[270]}
   );
   gpc1_1 gpc5563 (
      {stage0_59[489]},
      {stage1_59[271]}
   );
   gpc1_1 gpc5564 (
      {stage0_59[490]},
      {stage1_59[272]}
   );
   gpc1_1 gpc5565 (
      {stage0_59[491]},
      {stage1_59[273]}
   );
   gpc1_1 gpc5566 (
      {stage0_59[492]},
      {stage1_59[274]}
   );
   gpc1_1 gpc5567 (
      {stage0_59[493]},
      {stage1_59[275]}
   );
   gpc1_1 gpc5568 (
      {stage0_59[494]},
      {stage1_59[276]}
   );
   gpc1_1 gpc5569 (
      {stage0_59[495]},
      {stage1_59[277]}
   );
   gpc1_1 gpc5570 (
      {stage0_59[496]},
      {stage1_59[278]}
   );
   gpc1_1 gpc5571 (
      {stage0_59[497]},
      {stage1_59[279]}
   );
   gpc1_1 gpc5572 (
      {stage0_59[498]},
      {stage1_59[280]}
   );
   gpc1_1 gpc5573 (
      {stage0_59[499]},
      {stage1_59[281]}
   );
   gpc1_1 gpc5574 (
      {stage0_59[500]},
      {stage1_59[282]}
   );
   gpc1_1 gpc5575 (
      {stage0_59[501]},
      {stage1_59[283]}
   );
   gpc1_1 gpc5576 (
      {stage0_59[502]},
      {stage1_59[284]}
   );
   gpc1_1 gpc5577 (
      {stage0_59[503]},
      {stage1_59[285]}
   );
   gpc1_1 gpc5578 (
      {stage0_59[504]},
      {stage1_59[286]}
   );
   gpc1_1 gpc5579 (
      {stage0_59[505]},
      {stage1_59[287]}
   );
   gpc1_1 gpc5580 (
      {stage0_59[506]},
      {stage1_59[288]}
   );
   gpc1_1 gpc5581 (
      {stage0_59[507]},
      {stage1_59[289]}
   );
   gpc1_1 gpc5582 (
      {stage0_59[508]},
      {stage1_59[290]}
   );
   gpc1_1 gpc5583 (
      {stage0_59[509]},
      {stage1_59[291]}
   );
   gpc1_1 gpc5584 (
      {stage0_59[510]},
      {stage1_59[292]}
   );
   gpc1_1 gpc5585 (
      {stage0_59[511]},
      {stage1_59[293]}
   );
   gpc1_1 gpc5586 (
      {stage0_60[502]},
      {stage1_60[190]}
   );
   gpc1_1 gpc5587 (
      {stage0_60[503]},
      {stage1_60[191]}
   );
   gpc1_1 gpc5588 (
      {stage0_60[504]},
      {stage1_60[192]}
   );
   gpc1_1 gpc5589 (
      {stage0_60[505]},
      {stage1_60[193]}
   );
   gpc1_1 gpc5590 (
      {stage0_60[506]},
      {stage1_60[194]}
   );
   gpc1_1 gpc5591 (
      {stage0_60[507]},
      {stage1_60[195]}
   );
   gpc1_1 gpc5592 (
      {stage0_60[508]},
      {stage1_60[196]}
   );
   gpc1_1 gpc5593 (
      {stage0_60[509]},
      {stage1_60[197]}
   );
   gpc1_1 gpc5594 (
      {stage0_60[510]},
      {stage1_60[198]}
   );
   gpc1_1 gpc5595 (
      {stage0_60[511]},
      {stage1_60[199]}
   );
   gpc1_1 gpc5596 (
      {stage0_62[330]},
      {stage1_62[191]}
   );
   gpc1_1 gpc5597 (
      {stage0_62[331]},
      {stage1_62[192]}
   );
   gpc1_1 gpc5598 (
      {stage0_62[332]},
      {stage1_62[193]}
   );
   gpc1_1 gpc5599 (
      {stage0_62[333]},
      {stage1_62[194]}
   );
   gpc1_1 gpc5600 (
      {stage0_62[334]},
      {stage1_62[195]}
   );
   gpc1_1 gpc5601 (
      {stage0_62[335]},
      {stage1_62[196]}
   );
   gpc1_1 gpc5602 (
      {stage0_62[336]},
      {stage1_62[197]}
   );
   gpc1_1 gpc5603 (
      {stage0_62[337]},
      {stage1_62[198]}
   );
   gpc1_1 gpc5604 (
      {stage0_62[338]},
      {stage1_62[199]}
   );
   gpc1_1 gpc5605 (
      {stage0_62[339]},
      {stage1_62[200]}
   );
   gpc1_1 gpc5606 (
      {stage0_62[340]},
      {stage1_62[201]}
   );
   gpc1_1 gpc5607 (
      {stage0_62[341]},
      {stage1_62[202]}
   );
   gpc1_1 gpc5608 (
      {stage0_62[342]},
      {stage1_62[203]}
   );
   gpc1_1 gpc5609 (
      {stage0_62[343]},
      {stage1_62[204]}
   );
   gpc1_1 gpc5610 (
      {stage0_62[344]},
      {stage1_62[205]}
   );
   gpc1_1 gpc5611 (
      {stage0_62[345]},
      {stage1_62[206]}
   );
   gpc1_1 gpc5612 (
      {stage0_62[346]},
      {stage1_62[207]}
   );
   gpc1_1 gpc5613 (
      {stage0_62[347]},
      {stage1_62[208]}
   );
   gpc1_1 gpc5614 (
      {stage0_62[348]},
      {stage1_62[209]}
   );
   gpc1_1 gpc5615 (
      {stage0_62[349]},
      {stage1_62[210]}
   );
   gpc1_1 gpc5616 (
      {stage0_62[350]},
      {stage1_62[211]}
   );
   gpc1_1 gpc5617 (
      {stage0_62[351]},
      {stage1_62[212]}
   );
   gpc1_1 gpc5618 (
      {stage0_62[352]},
      {stage1_62[213]}
   );
   gpc1_1 gpc5619 (
      {stage0_62[353]},
      {stage1_62[214]}
   );
   gpc1_1 gpc5620 (
      {stage0_62[354]},
      {stage1_62[215]}
   );
   gpc1_1 gpc5621 (
      {stage0_62[355]},
      {stage1_62[216]}
   );
   gpc1_1 gpc5622 (
      {stage0_62[356]},
      {stage1_62[217]}
   );
   gpc1_1 gpc5623 (
      {stage0_62[357]},
      {stage1_62[218]}
   );
   gpc1_1 gpc5624 (
      {stage0_62[358]},
      {stage1_62[219]}
   );
   gpc1_1 gpc5625 (
      {stage0_62[359]},
      {stage1_62[220]}
   );
   gpc1_1 gpc5626 (
      {stage0_62[360]},
      {stage1_62[221]}
   );
   gpc1_1 gpc5627 (
      {stage0_62[361]},
      {stage1_62[222]}
   );
   gpc1_1 gpc5628 (
      {stage0_62[362]},
      {stage1_62[223]}
   );
   gpc1_1 gpc5629 (
      {stage0_62[363]},
      {stage1_62[224]}
   );
   gpc1_1 gpc5630 (
      {stage0_62[364]},
      {stage1_62[225]}
   );
   gpc1_1 gpc5631 (
      {stage0_62[365]},
      {stage1_62[226]}
   );
   gpc1_1 gpc5632 (
      {stage0_62[366]},
      {stage1_62[227]}
   );
   gpc1_1 gpc5633 (
      {stage0_62[367]},
      {stage1_62[228]}
   );
   gpc1_1 gpc5634 (
      {stage0_62[368]},
      {stage1_62[229]}
   );
   gpc1_1 gpc5635 (
      {stage0_62[369]},
      {stage1_62[230]}
   );
   gpc1_1 gpc5636 (
      {stage0_62[370]},
      {stage1_62[231]}
   );
   gpc1_1 gpc5637 (
      {stage0_62[371]},
      {stage1_62[232]}
   );
   gpc1_1 gpc5638 (
      {stage0_62[372]},
      {stage1_62[233]}
   );
   gpc1_1 gpc5639 (
      {stage0_62[373]},
      {stage1_62[234]}
   );
   gpc1_1 gpc5640 (
      {stage0_62[374]},
      {stage1_62[235]}
   );
   gpc1_1 gpc5641 (
      {stage0_62[375]},
      {stage1_62[236]}
   );
   gpc1_1 gpc5642 (
      {stage0_62[376]},
      {stage1_62[237]}
   );
   gpc1_1 gpc5643 (
      {stage0_62[377]},
      {stage1_62[238]}
   );
   gpc1_1 gpc5644 (
      {stage0_62[378]},
      {stage1_62[239]}
   );
   gpc1_1 gpc5645 (
      {stage0_62[379]},
      {stage1_62[240]}
   );
   gpc1_1 gpc5646 (
      {stage0_62[380]},
      {stage1_62[241]}
   );
   gpc1_1 gpc5647 (
      {stage0_62[381]},
      {stage1_62[242]}
   );
   gpc1_1 gpc5648 (
      {stage0_62[382]},
      {stage1_62[243]}
   );
   gpc1_1 gpc5649 (
      {stage0_62[383]},
      {stage1_62[244]}
   );
   gpc1_1 gpc5650 (
      {stage0_62[384]},
      {stage1_62[245]}
   );
   gpc1_1 gpc5651 (
      {stage0_62[385]},
      {stage1_62[246]}
   );
   gpc1_1 gpc5652 (
      {stage0_62[386]},
      {stage1_62[247]}
   );
   gpc1_1 gpc5653 (
      {stage0_62[387]},
      {stage1_62[248]}
   );
   gpc1_1 gpc5654 (
      {stage0_62[388]},
      {stage1_62[249]}
   );
   gpc1_1 gpc5655 (
      {stage0_62[389]},
      {stage1_62[250]}
   );
   gpc1_1 gpc5656 (
      {stage0_62[390]},
      {stage1_62[251]}
   );
   gpc1_1 gpc5657 (
      {stage0_62[391]},
      {stage1_62[252]}
   );
   gpc1_1 gpc5658 (
      {stage0_62[392]},
      {stage1_62[253]}
   );
   gpc1_1 gpc5659 (
      {stage0_62[393]},
      {stage1_62[254]}
   );
   gpc1_1 gpc5660 (
      {stage0_62[394]},
      {stage1_62[255]}
   );
   gpc1_1 gpc5661 (
      {stage0_62[395]},
      {stage1_62[256]}
   );
   gpc1_1 gpc5662 (
      {stage0_62[396]},
      {stage1_62[257]}
   );
   gpc1_1 gpc5663 (
      {stage0_62[397]},
      {stage1_62[258]}
   );
   gpc1_1 gpc5664 (
      {stage0_62[398]},
      {stage1_62[259]}
   );
   gpc1_1 gpc5665 (
      {stage0_62[399]},
      {stage1_62[260]}
   );
   gpc1_1 gpc5666 (
      {stage0_62[400]},
      {stage1_62[261]}
   );
   gpc1_1 gpc5667 (
      {stage0_62[401]},
      {stage1_62[262]}
   );
   gpc1_1 gpc5668 (
      {stage0_62[402]},
      {stage1_62[263]}
   );
   gpc1_1 gpc5669 (
      {stage0_62[403]},
      {stage1_62[264]}
   );
   gpc1_1 gpc5670 (
      {stage0_62[404]},
      {stage1_62[265]}
   );
   gpc1_1 gpc5671 (
      {stage0_62[405]},
      {stage1_62[266]}
   );
   gpc1_1 gpc5672 (
      {stage0_62[406]},
      {stage1_62[267]}
   );
   gpc1_1 gpc5673 (
      {stage0_62[407]},
      {stage1_62[268]}
   );
   gpc1_1 gpc5674 (
      {stage0_62[408]},
      {stage1_62[269]}
   );
   gpc1_1 gpc5675 (
      {stage0_62[409]},
      {stage1_62[270]}
   );
   gpc1_1 gpc5676 (
      {stage0_62[410]},
      {stage1_62[271]}
   );
   gpc1_1 gpc5677 (
      {stage0_62[411]},
      {stage1_62[272]}
   );
   gpc1_1 gpc5678 (
      {stage0_62[412]},
      {stage1_62[273]}
   );
   gpc1_1 gpc5679 (
      {stage0_62[413]},
      {stage1_62[274]}
   );
   gpc1_1 gpc5680 (
      {stage0_62[414]},
      {stage1_62[275]}
   );
   gpc1_1 gpc5681 (
      {stage0_62[415]},
      {stage1_62[276]}
   );
   gpc1_1 gpc5682 (
      {stage0_62[416]},
      {stage1_62[277]}
   );
   gpc1_1 gpc5683 (
      {stage0_62[417]},
      {stage1_62[278]}
   );
   gpc1_1 gpc5684 (
      {stage0_62[418]},
      {stage1_62[279]}
   );
   gpc1_1 gpc5685 (
      {stage0_62[419]},
      {stage1_62[280]}
   );
   gpc1_1 gpc5686 (
      {stage0_62[420]},
      {stage1_62[281]}
   );
   gpc1_1 gpc5687 (
      {stage0_62[421]},
      {stage1_62[282]}
   );
   gpc1_1 gpc5688 (
      {stage0_62[422]},
      {stage1_62[283]}
   );
   gpc1_1 gpc5689 (
      {stage0_62[423]},
      {stage1_62[284]}
   );
   gpc1_1 gpc5690 (
      {stage0_62[424]},
      {stage1_62[285]}
   );
   gpc1_1 gpc5691 (
      {stage0_62[425]},
      {stage1_62[286]}
   );
   gpc1_1 gpc5692 (
      {stage0_62[426]},
      {stage1_62[287]}
   );
   gpc1_1 gpc5693 (
      {stage0_62[427]},
      {stage1_62[288]}
   );
   gpc1_1 gpc5694 (
      {stage0_62[428]},
      {stage1_62[289]}
   );
   gpc1_1 gpc5695 (
      {stage0_62[429]},
      {stage1_62[290]}
   );
   gpc1_1 gpc5696 (
      {stage0_62[430]},
      {stage1_62[291]}
   );
   gpc1_1 gpc5697 (
      {stage0_62[431]},
      {stage1_62[292]}
   );
   gpc1_1 gpc5698 (
      {stage0_62[432]},
      {stage1_62[293]}
   );
   gpc1_1 gpc5699 (
      {stage0_62[433]},
      {stage1_62[294]}
   );
   gpc1_1 gpc5700 (
      {stage0_62[434]},
      {stage1_62[295]}
   );
   gpc1_1 gpc5701 (
      {stage0_62[435]},
      {stage1_62[296]}
   );
   gpc1_1 gpc5702 (
      {stage0_62[436]},
      {stage1_62[297]}
   );
   gpc1_1 gpc5703 (
      {stage0_62[437]},
      {stage1_62[298]}
   );
   gpc1_1 gpc5704 (
      {stage0_62[438]},
      {stage1_62[299]}
   );
   gpc1_1 gpc5705 (
      {stage0_62[439]},
      {stage1_62[300]}
   );
   gpc1_1 gpc5706 (
      {stage0_62[440]},
      {stage1_62[301]}
   );
   gpc1_1 gpc5707 (
      {stage0_62[441]},
      {stage1_62[302]}
   );
   gpc1_1 gpc5708 (
      {stage0_62[442]},
      {stage1_62[303]}
   );
   gpc1_1 gpc5709 (
      {stage0_62[443]},
      {stage1_62[304]}
   );
   gpc1_1 gpc5710 (
      {stage0_62[444]},
      {stage1_62[305]}
   );
   gpc1_1 gpc5711 (
      {stage0_62[445]},
      {stage1_62[306]}
   );
   gpc1_1 gpc5712 (
      {stage0_62[446]},
      {stage1_62[307]}
   );
   gpc1_1 gpc5713 (
      {stage0_62[447]},
      {stage1_62[308]}
   );
   gpc1_1 gpc5714 (
      {stage0_62[448]},
      {stage1_62[309]}
   );
   gpc1_1 gpc5715 (
      {stage0_62[449]},
      {stage1_62[310]}
   );
   gpc1_1 gpc5716 (
      {stage0_62[450]},
      {stage1_62[311]}
   );
   gpc1_1 gpc5717 (
      {stage0_62[451]},
      {stage1_62[312]}
   );
   gpc1_1 gpc5718 (
      {stage0_62[452]},
      {stage1_62[313]}
   );
   gpc1_1 gpc5719 (
      {stage0_62[453]},
      {stage1_62[314]}
   );
   gpc1_1 gpc5720 (
      {stage0_62[454]},
      {stage1_62[315]}
   );
   gpc1_1 gpc5721 (
      {stage0_62[455]},
      {stage1_62[316]}
   );
   gpc1_1 gpc5722 (
      {stage0_62[456]},
      {stage1_62[317]}
   );
   gpc1_1 gpc5723 (
      {stage0_62[457]},
      {stage1_62[318]}
   );
   gpc1_1 gpc5724 (
      {stage0_62[458]},
      {stage1_62[319]}
   );
   gpc1_1 gpc5725 (
      {stage0_62[459]},
      {stage1_62[320]}
   );
   gpc1_1 gpc5726 (
      {stage0_62[460]},
      {stage1_62[321]}
   );
   gpc1_1 gpc5727 (
      {stage0_62[461]},
      {stage1_62[322]}
   );
   gpc1_1 gpc5728 (
      {stage0_62[462]},
      {stage1_62[323]}
   );
   gpc1_1 gpc5729 (
      {stage0_62[463]},
      {stage1_62[324]}
   );
   gpc1_1 gpc5730 (
      {stage0_62[464]},
      {stage1_62[325]}
   );
   gpc1_1 gpc5731 (
      {stage0_62[465]},
      {stage1_62[326]}
   );
   gpc1_1 gpc5732 (
      {stage0_62[466]},
      {stage1_62[327]}
   );
   gpc1_1 gpc5733 (
      {stage0_62[467]},
      {stage1_62[328]}
   );
   gpc1_1 gpc5734 (
      {stage0_62[468]},
      {stage1_62[329]}
   );
   gpc1_1 gpc5735 (
      {stage0_62[469]},
      {stage1_62[330]}
   );
   gpc1_1 gpc5736 (
      {stage0_62[470]},
      {stage1_62[331]}
   );
   gpc1_1 gpc5737 (
      {stage0_62[471]},
      {stage1_62[332]}
   );
   gpc1_1 gpc5738 (
      {stage0_62[472]},
      {stage1_62[333]}
   );
   gpc1_1 gpc5739 (
      {stage0_62[473]},
      {stage1_62[334]}
   );
   gpc1_1 gpc5740 (
      {stage0_62[474]},
      {stage1_62[335]}
   );
   gpc1_1 gpc5741 (
      {stage0_62[475]},
      {stage1_62[336]}
   );
   gpc1_1 gpc5742 (
      {stage0_62[476]},
      {stage1_62[337]}
   );
   gpc1_1 gpc5743 (
      {stage0_62[477]},
      {stage1_62[338]}
   );
   gpc1_1 gpc5744 (
      {stage0_62[478]},
      {stage1_62[339]}
   );
   gpc1_1 gpc5745 (
      {stage0_62[479]},
      {stage1_62[340]}
   );
   gpc1_1 gpc5746 (
      {stage0_62[480]},
      {stage1_62[341]}
   );
   gpc1_1 gpc5747 (
      {stage0_62[481]},
      {stage1_62[342]}
   );
   gpc1_1 gpc5748 (
      {stage0_62[482]},
      {stage1_62[343]}
   );
   gpc1_1 gpc5749 (
      {stage0_62[483]},
      {stage1_62[344]}
   );
   gpc1_1 gpc5750 (
      {stage0_62[484]},
      {stage1_62[345]}
   );
   gpc1_1 gpc5751 (
      {stage0_62[485]},
      {stage1_62[346]}
   );
   gpc1_1 gpc5752 (
      {stage0_62[486]},
      {stage1_62[347]}
   );
   gpc1_1 gpc5753 (
      {stage0_62[487]},
      {stage1_62[348]}
   );
   gpc1_1 gpc5754 (
      {stage0_62[488]},
      {stage1_62[349]}
   );
   gpc1_1 gpc5755 (
      {stage0_62[489]},
      {stage1_62[350]}
   );
   gpc1_1 gpc5756 (
      {stage0_62[490]},
      {stage1_62[351]}
   );
   gpc1_1 gpc5757 (
      {stage0_62[491]},
      {stage1_62[352]}
   );
   gpc1_1 gpc5758 (
      {stage0_62[492]},
      {stage1_62[353]}
   );
   gpc1_1 gpc5759 (
      {stage0_62[493]},
      {stage1_62[354]}
   );
   gpc1_1 gpc5760 (
      {stage0_62[494]},
      {stage1_62[355]}
   );
   gpc1_1 gpc5761 (
      {stage0_62[495]},
      {stage1_62[356]}
   );
   gpc1_1 gpc5762 (
      {stage0_62[496]},
      {stage1_62[357]}
   );
   gpc1_1 gpc5763 (
      {stage0_62[497]},
      {stage1_62[358]}
   );
   gpc1_1 gpc5764 (
      {stage0_62[498]},
      {stage1_62[359]}
   );
   gpc1_1 gpc5765 (
      {stage0_62[499]},
      {stage1_62[360]}
   );
   gpc1_1 gpc5766 (
      {stage0_62[500]},
      {stage1_62[361]}
   );
   gpc1_1 gpc5767 (
      {stage0_62[501]},
      {stage1_62[362]}
   );
   gpc1_1 gpc5768 (
      {stage0_62[502]},
      {stage1_62[363]}
   );
   gpc1_1 gpc5769 (
      {stage0_62[503]},
      {stage1_62[364]}
   );
   gpc1_1 gpc5770 (
      {stage0_62[504]},
      {stage1_62[365]}
   );
   gpc1_1 gpc5771 (
      {stage0_62[505]},
      {stage1_62[366]}
   );
   gpc1_1 gpc5772 (
      {stage0_62[506]},
      {stage1_62[367]}
   );
   gpc1_1 gpc5773 (
      {stage0_62[507]},
      {stage1_62[368]}
   );
   gpc1_1 gpc5774 (
      {stage0_62[508]},
      {stage1_62[369]}
   );
   gpc1_1 gpc5775 (
      {stage0_62[509]},
      {stage1_62[370]}
   );
   gpc1_1 gpc5776 (
      {stage0_62[510]},
      {stage1_62[371]}
   );
   gpc1_1 gpc5777 (
      {stage0_62[511]},
      {stage1_62[372]}
   );
   gpc1_1 gpc5778 (
      {stage0_63[342]},
      {stage1_63[125]}
   );
   gpc1_1 gpc5779 (
      {stage0_63[343]},
      {stage1_63[126]}
   );
   gpc1_1 gpc5780 (
      {stage0_63[344]},
      {stage1_63[127]}
   );
   gpc1_1 gpc5781 (
      {stage0_63[345]},
      {stage1_63[128]}
   );
   gpc1_1 gpc5782 (
      {stage0_63[346]},
      {stage1_63[129]}
   );
   gpc1_1 gpc5783 (
      {stage0_63[347]},
      {stage1_63[130]}
   );
   gpc1_1 gpc5784 (
      {stage0_63[348]},
      {stage1_63[131]}
   );
   gpc1_1 gpc5785 (
      {stage0_63[349]},
      {stage1_63[132]}
   );
   gpc1_1 gpc5786 (
      {stage0_63[350]},
      {stage1_63[133]}
   );
   gpc1_1 gpc5787 (
      {stage0_63[351]},
      {stage1_63[134]}
   );
   gpc1_1 gpc5788 (
      {stage0_63[352]},
      {stage1_63[135]}
   );
   gpc1_1 gpc5789 (
      {stage0_63[353]},
      {stage1_63[136]}
   );
   gpc1_1 gpc5790 (
      {stage0_63[354]},
      {stage1_63[137]}
   );
   gpc1_1 gpc5791 (
      {stage0_63[355]},
      {stage1_63[138]}
   );
   gpc1_1 gpc5792 (
      {stage0_63[356]},
      {stage1_63[139]}
   );
   gpc1_1 gpc5793 (
      {stage0_63[357]},
      {stage1_63[140]}
   );
   gpc1_1 gpc5794 (
      {stage0_63[358]},
      {stage1_63[141]}
   );
   gpc1_1 gpc5795 (
      {stage0_63[359]},
      {stage1_63[142]}
   );
   gpc1_1 gpc5796 (
      {stage0_63[360]},
      {stage1_63[143]}
   );
   gpc1_1 gpc5797 (
      {stage0_63[361]},
      {stage1_63[144]}
   );
   gpc1_1 gpc5798 (
      {stage0_63[362]},
      {stage1_63[145]}
   );
   gpc1_1 gpc5799 (
      {stage0_63[363]},
      {stage1_63[146]}
   );
   gpc1_1 gpc5800 (
      {stage0_63[364]},
      {stage1_63[147]}
   );
   gpc1_1 gpc5801 (
      {stage0_63[365]},
      {stage1_63[148]}
   );
   gpc1_1 gpc5802 (
      {stage0_63[366]},
      {stage1_63[149]}
   );
   gpc1_1 gpc5803 (
      {stage0_63[367]},
      {stage1_63[150]}
   );
   gpc1_1 gpc5804 (
      {stage0_63[368]},
      {stage1_63[151]}
   );
   gpc1_1 gpc5805 (
      {stage0_63[369]},
      {stage1_63[152]}
   );
   gpc1_1 gpc5806 (
      {stage0_63[370]},
      {stage1_63[153]}
   );
   gpc1_1 gpc5807 (
      {stage0_63[371]},
      {stage1_63[154]}
   );
   gpc1_1 gpc5808 (
      {stage0_63[372]},
      {stage1_63[155]}
   );
   gpc1_1 gpc5809 (
      {stage0_63[373]},
      {stage1_63[156]}
   );
   gpc1_1 gpc5810 (
      {stage0_63[374]},
      {stage1_63[157]}
   );
   gpc1_1 gpc5811 (
      {stage0_63[375]},
      {stage1_63[158]}
   );
   gpc1_1 gpc5812 (
      {stage0_63[376]},
      {stage1_63[159]}
   );
   gpc1_1 gpc5813 (
      {stage0_63[377]},
      {stage1_63[160]}
   );
   gpc1_1 gpc5814 (
      {stage0_63[378]},
      {stage1_63[161]}
   );
   gpc1_1 gpc5815 (
      {stage0_63[379]},
      {stage1_63[162]}
   );
   gpc1_1 gpc5816 (
      {stage0_63[380]},
      {stage1_63[163]}
   );
   gpc1_1 gpc5817 (
      {stage0_63[381]},
      {stage1_63[164]}
   );
   gpc1_1 gpc5818 (
      {stage0_63[382]},
      {stage1_63[165]}
   );
   gpc1_1 gpc5819 (
      {stage0_63[383]},
      {stage1_63[166]}
   );
   gpc1_1 gpc5820 (
      {stage0_63[384]},
      {stage1_63[167]}
   );
   gpc1_1 gpc5821 (
      {stage0_63[385]},
      {stage1_63[168]}
   );
   gpc1_1 gpc5822 (
      {stage0_63[386]},
      {stage1_63[169]}
   );
   gpc1_1 gpc5823 (
      {stage0_63[387]},
      {stage1_63[170]}
   );
   gpc1_1 gpc5824 (
      {stage0_63[388]},
      {stage1_63[171]}
   );
   gpc1_1 gpc5825 (
      {stage0_63[389]},
      {stage1_63[172]}
   );
   gpc1_1 gpc5826 (
      {stage0_63[390]},
      {stage1_63[173]}
   );
   gpc1_1 gpc5827 (
      {stage0_63[391]},
      {stage1_63[174]}
   );
   gpc1_1 gpc5828 (
      {stage0_63[392]},
      {stage1_63[175]}
   );
   gpc1_1 gpc5829 (
      {stage0_63[393]},
      {stage1_63[176]}
   );
   gpc1_1 gpc5830 (
      {stage0_63[394]},
      {stage1_63[177]}
   );
   gpc1_1 gpc5831 (
      {stage0_63[395]},
      {stage1_63[178]}
   );
   gpc1_1 gpc5832 (
      {stage0_63[396]},
      {stage1_63[179]}
   );
   gpc1_1 gpc5833 (
      {stage0_63[397]},
      {stage1_63[180]}
   );
   gpc1_1 gpc5834 (
      {stage0_63[398]},
      {stage1_63[181]}
   );
   gpc1_1 gpc5835 (
      {stage0_63[399]},
      {stage1_63[182]}
   );
   gpc1_1 gpc5836 (
      {stage0_63[400]},
      {stage1_63[183]}
   );
   gpc1_1 gpc5837 (
      {stage0_63[401]},
      {stage1_63[184]}
   );
   gpc1_1 gpc5838 (
      {stage0_63[402]},
      {stage1_63[185]}
   );
   gpc1_1 gpc5839 (
      {stage0_63[403]},
      {stage1_63[186]}
   );
   gpc1_1 gpc5840 (
      {stage0_63[404]},
      {stage1_63[187]}
   );
   gpc1_1 gpc5841 (
      {stage0_63[405]},
      {stage1_63[188]}
   );
   gpc1_1 gpc5842 (
      {stage0_63[406]},
      {stage1_63[189]}
   );
   gpc1_1 gpc5843 (
      {stage0_63[407]},
      {stage1_63[190]}
   );
   gpc1_1 gpc5844 (
      {stage0_63[408]},
      {stage1_63[191]}
   );
   gpc1_1 gpc5845 (
      {stage0_63[409]},
      {stage1_63[192]}
   );
   gpc1_1 gpc5846 (
      {stage0_63[410]},
      {stage1_63[193]}
   );
   gpc1_1 gpc5847 (
      {stage0_63[411]},
      {stage1_63[194]}
   );
   gpc1_1 gpc5848 (
      {stage0_63[412]},
      {stage1_63[195]}
   );
   gpc1_1 gpc5849 (
      {stage0_63[413]},
      {stage1_63[196]}
   );
   gpc1_1 gpc5850 (
      {stage0_63[414]},
      {stage1_63[197]}
   );
   gpc1_1 gpc5851 (
      {stage0_63[415]},
      {stage1_63[198]}
   );
   gpc1_1 gpc5852 (
      {stage0_63[416]},
      {stage1_63[199]}
   );
   gpc1_1 gpc5853 (
      {stage0_63[417]},
      {stage1_63[200]}
   );
   gpc1_1 gpc5854 (
      {stage0_63[418]},
      {stage1_63[201]}
   );
   gpc1_1 gpc5855 (
      {stage0_63[419]},
      {stage1_63[202]}
   );
   gpc1_1 gpc5856 (
      {stage0_63[420]},
      {stage1_63[203]}
   );
   gpc1_1 gpc5857 (
      {stage0_63[421]},
      {stage1_63[204]}
   );
   gpc1_1 gpc5858 (
      {stage0_63[422]},
      {stage1_63[205]}
   );
   gpc1_1 gpc5859 (
      {stage0_63[423]},
      {stage1_63[206]}
   );
   gpc1_1 gpc5860 (
      {stage0_63[424]},
      {stage1_63[207]}
   );
   gpc1_1 gpc5861 (
      {stage0_63[425]},
      {stage1_63[208]}
   );
   gpc1_1 gpc5862 (
      {stage0_63[426]},
      {stage1_63[209]}
   );
   gpc1_1 gpc5863 (
      {stage0_63[427]},
      {stage1_63[210]}
   );
   gpc1_1 gpc5864 (
      {stage0_63[428]},
      {stage1_63[211]}
   );
   gpc1_1 gpc5865 (
      {stage0_63[429]},
      {stage1_63[212]}
   );
   gpc1_1 gpc5866 (
      {stage0_63[430]},
      {stage1_63[213]}
   );
   gpc1_1 gpc5867 (
      {stage0_63[431]},
      {stage1_63[214]}
   );
   gpc1_1 gpc5868 (
      {stage0_63[432]},
      {stage1_63[215]}
   );
   gpc1_1 gpc5869 (
      {stage0_63[433]},
      {stage1_63[216]}
   );
   gpc1_1 gpc5870 (
      {stage0_63[434]},
      {stage1_63[217]}
   );
   gpc1_1 gpc5871 (
      {stage0_63[435]},
      {stage1_63[218]}
   );
   gpc1_1 gpc5872 (
      {stage0_63[436]},
      {stage1_63[219]}
   );
   gpc1_1 gpc5873 (
      {stage0_63[437]},
      {stage1_63[220]}
   );
   gpc1_1 gpc5874 (
      {stage0_63[438]},
      {stage1_63[221]}
   );
   gpc1_1 gpc5875 (
      {stage0_63[439]},
      {stage1_63[222]}
   );
   gpc1_1 gpc5876 (
      {stage0_63[440]},
      {stage1_63[223]}
   );
   gpc1_1 gpc5877 (
      {stage0_63[441]},
      {stage1_63[224]}
   );
   gpc1_1 gpc5878 (
      {stage0_63[442]},
      {stage1_63[225]}
   );
   gpc1_1 gpc5879 (
      {stage0_63[443]},
      {stage1_63[226]}
   );
   gpc1_1 gpc5880 (
      {stage0_63[444]},
      {stage1_63[227]}
   );
   gpc1_1 gpc5881 (
      {stage0_63[445]},
      {stage1_63[228]}
   );
   gpc1_1 gpc5882 (
      {stage0_63[446]},
      {stage1_63[229]}
   );
   gpc1_1 gpc5883 (
      {stage0_63[447]},
      {stage1_63[230]}
   );
   gpc1_1 gpc5884 (
      {stage0_63[448]},
      {stage1_63[231]}
   );
   gpc1_1 gpc5885 (
      {stage0_63[449]},
      {stage1_63[232]}
   );
   gpc1_1 gpc5886 (
      {stage0_63[450]},
      {stage1_63[233]}
   );
   gpc1_1 gpc5887 (
      {stage0_63[451]},
      {stage1_63[234]}
   );
   gpc1_1 gpc5888 (
      {stage0_63[452]},
      {stage1_63[235]}
   );
   gpc1_1 gpc5889 (
      {stage0_63[453]},
      {stage1_63[236]}
   );
   gpc1_1 gpc5890 (
      {stage0_63[454]},
      {stage1_63[237]}
   );
   gpc1_1 gpc5891 (
      {stage0_63[455]},
      {stage1_63[238]}
   );
   gpc1_1 gpc5892 (
      {stage0_63[456]},
      {stage1_63[239]}
   );
   gpc1_1 gpc5893 (
      {stage0_63[457]},
      {stage1_63[240]}
   );
   gpc1_1 gpc5894 (
      {stage0_63[458]},
      {stage1_63[241]}
   );
   gpc1_1 gpc5895 (
      {stage0_63[459]},
      {stage1_63[242]}
   );
   gpc1_1 gpc5896 (
      {stage0_63[460]},
      {stage1_63[243]}
   );
   gpc1_1 gpc5897 (
      {stage0_63[461]},
      {stage1_63[244]}
   );
   gpc1_1 gpc5898 (
      {stage0_63[462]},
      {stage1_63[245]}
   );
   gpc1_1 gpc5899 (
      {stage0_63[463]},
      {stage1_63[246]}
   );
   gpc1_1 gpc5900 (
      {stage0_63[464]},
      {stage1_63[247]}
   );
   gpc1_1 gpc5901 (
      {stage0_63[465]},
      {stage1_63[248]}
   );
   gpc1_1 gpc5902 (
      {stage0_63[466]},
      {stage1_63[249]}
   );
   gpc1_1 gpc5903 (
      {stage0_63[467]},
      {stage1_63[250]}
   );
   gpc1_1 gpc5904 (
      {stage0_63[468]},
      {stage1_63[251]}
   );
   gpc1_1 gpc5905 (
      {stage0_63[469]},
      {stage1_63[252]}
   );
   gpc1_1 gpc5906 (
      {stage0_63[470]},
      {stage1_63[253]}
   );
   gpc1_1 gpc5907 (
      {stage0_63[471]},
      {stage1_63[254]}
   );
   gpc1_1 gpc5908 (
      {stage0_63[472]},
      {stage1_63[255]}
   );
   gpc1_1 gpc5909 (
      {stage0_63[473]},
      {stage1_63[256]}
   );
   gpc1_1 gpc5910 (
      {stage0_63[474]},
      {stage1_63[257]}
   );
   gpc1_1 gpc5911 (
      {stage0_63[475]},
      {stage1_63[258]}
   );
   gpc1_1 gpc5912 (
      {stage0_63[476]},
      {stage1_63[259]}
   );
   gpc1_1 gpc5913 (
      {stage0_63[477]},
      {stage1_63[260]}
   );
   gpc1_1 gpc5914 (
      {stage0_63[478]},
      {stage1_63[261]}
   );
   gpc1_1 gpc5915 (
      {stage0_63[479]},
      {stage1_63[262]}
   );
   gpc1_1 gpc5916 (
      {stage0_63[480]},
      {stage1_63[263]}
   );
   gpc1_1 gpc5917 (
      {stage0_63[481]},
      {stage1_63[264]}
   );
   gpc1_1 gpc5918 (
      {stage0_63[482]},
      {stage1_63[265]}
   );
   gpc1_1 gpc5919 (
      {stage0_63[483]},
      {stage1_63[266]}
   );
   gpc1_1 gpc5920 (
      {stage0_63[484]},
      {stage1_63[267]}
   );
   gpc1_1 gpc5921 (
      {stage0_63[485]},
      {stage1_63[268]}
   );
   gpc1_1 gpc5922 (
      {stage0_63[486]},
      {stage1_63[269]}
   );
   gpc1_1 gpc5923 (
      {stage0_63[487]},
      {stage1_63[270]}
   );
   gpc1_1 gpc5924 (
      {stage0_63[488]},
      {stage1_63[271]}
   );
   gpc1_1 gpc5925 (
      {stage0_63[489]},
      {stage1_63[272]}
   );
   gpc1_1 gpc5926 (
      {stage0_63[490]},
      {stage1_63[273]}
   );
   gpc1_1 gpc5927 (
      {stage0_63[491]},
      {stage1_63[274]}
   );
   gpc1_1 gpc5928 (
      {stage0_63[492]},
      {stage1_63[275]}
   );
   gpc1_1 gpc5929 (
      {stage0_63[493]},
      {stage1_63[276]}
   );
   gpc1_1 gpc5930 (
      {stage0_63[494]},
      {stage1_63[277]}
   );
   gpc1_1 gpc5931 (
      {stage0_63[495]},
      {stage1_63[278]}
   );
   gpc1_1 gpc5932 (
      {stage0_63[496]},
      {stage1_63[279]}
   );
   gpc1_1 gpc5933 (
      {stage0_63[497]},
      {stage1_63[280]}
   );
   gpc1_1 gpc5934 (
      {stage0_63[498]},
      {stage1_63[281]}
   );
   gpc1_1 gpc5935 (
      {stage0_63[499]},
      {stage1_63[282]}
   );
   gpc1_1 gpc5936 (
      {stage0_63[500]},
      {stage1_63[283]}
   );
   gpc1_1 gpc5937 (
      {stage0_63[501]},
      {stage1_63[284]}
   );
   gpc1_1 gpc5938 (
      {stage0_63[502]},
      {stage1_63[285]}
   );
   gpc1_1 gpc5939 (
      {stage0_63[503]},
      {stage1_63[286]}
   );
   gpc1_1 gpc5940 (
      {stage0_63[504]},
      {stage1_63[287]}
   );
   gpc1_1 gpc5941 (
      {stage0_63[505]},
      {stage1_63[288]}
   );
   gpc1_1 gpc5942 (
      {stage0_63[506]},
      {stage1_63[289]}
   );
   gpc1_1 gpc5943 (
      {stage0_63[507]},
      {stage1_63[290]}
   );
   gpc1_1 gpc5944 (
      {stage0_63[508]},
      {stage1_63[291]}
   );
   gpc1_1 gpc5945 (
      {stage0_63[509]},
      {stage1_63[292]}
   );
   gpc1_1 gpc5946 (
      {stage0_63[510]},
      {stage1_63[293]}
   );
   gpc1_1 gpc5947 (
      {stage0_63[511]},
      {stage1_63[294]}
   );
   gpc1163_5 gpc5948 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc5949 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc5950 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc5951 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc5952 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc5953 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc5954 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc5955 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc5956 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc5957 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc5958 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc5959 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc5960 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc5961 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc5962 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc5963 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc5964 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc5965 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc5966 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc5967 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc5968 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc5969 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc5970 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc5971 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc5972 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc615_5 gpc5973 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106]},
      {stage1_1[96]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc615_5 gpc5974 (
      {stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111]},
      {stage1_1[97]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc5975 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[0],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc5976 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[1],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc5977 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[2],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc5978 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[3],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc5979 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[4],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc5980 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[5],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc5981 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[6],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc5982 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage2_5[7],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc5983 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69]},
      {stage2_5[8],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc5984 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage2_5[9],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc5985 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage2_5[10],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc5986 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], 1'b0},
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87]},
      {stage2_5[11],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc5987 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[12],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc5988 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[13],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc5989 (
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[14],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc5990 (
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[15],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc5991 (
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[16],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc606_5 gpc5992 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[17],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc606_5 gpc5993 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[18],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc606_5 gpc5994 (
      {stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[19],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc5995 (
      {stage1_2[130], stage1_2[131], stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[20],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc5996 (
      {stage1_2[136], stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[21],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc606_5 gpc5997 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[22],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc606_5 gpc5998 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152], stage1_2[153]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[23],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc606_5 gpc5999 (
      {stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157], stage1_2[158], stage1_2[159]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[24],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc606_5 gpc6000 (
      {stage1_2[160], stage1_2[161], stage1_2[162], stage1_2[163], stage1_2[164], stage1_2[165]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[25],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc606_5 gpc6001 (
      {stage1_2[166], stage1_2[167], stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[26],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc606_5 gpc6002 (
      {stage1_2[172], stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[27],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc606_5 gpc6003 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182], stage1_2[183]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[28],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc606_5 gpc6004 (
      {stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187], stage1_2[188], stage1_2[189]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[29],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc606_5 gpc6005 (
      {stage1_2[190], stage1_2[191], stage1_2[192], stage1_2[193], stage1_2[194], stage1_2[195]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[30],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc606_5 gpc6006 (
      {stage1_2[196], stage1_2[197], stage1_2[198], stage1_2[199], stage1_2[200], stage1_2[201]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[31],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc606_5 gpc6007 (
      {stage1_2[202], stage1_2[203], stage1_2[204], stage1_2[205], stage1_2[206], stage1_2[207]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[32],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc1415_5 gpc6008 (
      {stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92]},
      {stage1_4[126]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[21],stage2_5[33],stage2_4[60],stage2_3[60]}
   );
   gpc1415_5 gpc6009 (
      {stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage1_4[127]},
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7]},
      {stage1_6[1]},
      {stage2_7[1],stage2_6[22],stage2_5[34],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc6010 (
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102]},
      {stage1_4[128]},
      {stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13]},
      {stage2_7[2],stage2_6[23],stage2_5[35],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc6011 (
      {stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage1_4[129]},
      {stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19]},
      {stage2_7[3],stage2_6[24],stage2_5[36],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc6012 (
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112]},
      {stage1_4[130]},
      {stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25]},
      {stage2_7[4],stage2_6[25],stage2_5[37],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc6013 (
      {stage1_3[113], stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117]},
      {stage1_4[131]},
      {stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31]},
      {stage2_7[5],stage2_6[26],stage2_5[38],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc6014 (
      {stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122]},
      {stage1_4[132]},
      {stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37]},
      {stage2_7[6],stage2_6[27],stage2_5[39],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc6015 (
      {stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage1_4[133]},
      {stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43]},
      {stage2_7[7],stage2_6[28],stage2_5[40],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc6016 (
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132]},
      {stage1_4[134]},
      {stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49]},
      {stage2_7[8],stage2_6[29],stage2_5[41],stage2_4[68],stage2_3[68]}
   );
   gpc623_5 gpc6017 (
      {stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[135], stage1_4[136]},
      {stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55]},
      {stage2_7[9],stage2_6[30],stage2_5[42],stage2_4[69],stage2_3[69]}
   );
   gpc623_5 gpc6018 (
      {stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[137], stage1_4[138]},
      {stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61]},
      {stage2_7[10],stage2_6[31],stage2_5[43],stage2_4[70],stage2_3[70]}
   );
   gpc606_5 gpc6019 (
      {stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[11],stage2_6[32],stage2_5[44],stage2_4[71]}
   );
   gpc606_5 gpc6020 (
      {stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[12],stage2_6[33],stage2_5[45],stage2_4[72]}
   );
   gpc606_5 gpc6021 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[13],stage2_6[34],stage2_5[46],stage2_4[73]}
   );
   gpc606_5 gpc6022 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162]},
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage2_8[3],stage2_7[14],stage2_6[35],stage2_5[47],stage2_4[74]}
   );
   gpc606_5 gpc6023 (
      {stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168]},
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage2_8[4],stage2_7[15],stage2_6[36],stage2_5[48],stage2_4[75]}
   );
   gpc606_5 gpc6024 (
      {stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174]},
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36], stage1_6[37]},
      {stage2_8[5],stage2_7[16],stage2_6[37],stage2_5[49],stage2_4[76]}
   );
   gpc606_5 gpc6025 (
      {stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42], stage1_6[43]},
      {stage2_8[6],stage2_7[17],stage2_6[38],stage2_5[50],stage2_4[77]}
   );
   gpc606_5 gpc6026 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49]},
      {stage2_8[7],stage2_7[18],stage2_6[39],stage2_5[51],stage2_4[78]}
   );
   gpc606_5 gpc6027 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192]},
      {stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage2_8[8],stage2_7[19],stage2_6[40],stage2_5[52],stage2_4[79]}
   );
   gpc606_5 gpc6028 (
      {stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198]},
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage2_8[9],stage2_7[20],stage2_6[41],stage2_5[53],stage2_4[80]}
   );
   gpc606_5 gpc6029 (
      {stage1_4[199], stage1_4[200], stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204]},
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66], stage1_6[67]},
      {stage2_8[10],stage2_7[21],stage2_6[42],stage2_5[54],stage2_4[81]}
   );
   gpc606_5 gpc6030 (
      {stage1_4[205], stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72], stage1_6[73]},
      {stage2_8[11],stage2_7[22],stage2_6[43],stage2_5[55],stage2_4[82]}
   );
   gpc606_5 gpc6031 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79]},
      {stage2_8[12],stage2_7[23],stage2_6[44],stage2_5[56],stage2_4[83]}
   );
   gpc606_5 gpc6032 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221], stage1_4[222]},
      {stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage2_8[13],stage2_7[24],stage2_6[45],stage2_5[57],stage2_4[84]}
   );
   gpc606_5 gpc6033 (
      {stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227], stage1_4[228]},
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage2_8[14],stage2_7[25],stage2_6[46],stage2_5[58],stage2_4[85]}
   );
   gpc606_5 gpc6034 (
      {stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233], stage1_4[234]},
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96], stage1_6[97]},
      {stage2_8[15],stage2_7[26],stage2_6[47],stage2_5[59],stage2_4[86]}
   );
   gpc606_5 gpc6035 (
      {stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239], stage1_4[240]},
      {stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102], stage1_6[103]},
      {stage2_8[16],stage2_7[27],stage2_6[48],stage2_5[60],stage2_4[87]}
   );
   gpc606_5 gpc6036 (
      {stage1_4[241], stage1_4[242], stage1_4[243], stage1_4[244], stage1_4[245], stage1_4[246]},
      {stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108], stage1_6[109]},
      {stage2_8[17],stage2_7[28],stage2_6[49],stage2_5[61],stage2_4[88]}
   );
   gpc606_5 gpc6037 (
      {stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[18],stage2_7[29],stage2_6[50],stage2_5[62]}
   );
   gpc606_5 gpc6038 (
      {stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[19],stage2_7[30],stage2_6[51],stage2_5[63]}
   );
   gpc606_5 gpc6039 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[20],stage2_7[31],stage2_6[52],stage2_5[64]}
   );
   gpc606_5 gpc6040 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[21],stage2_7[32],stage2_6[53],stage2_5[65]}
   );
   gpc606_5 gpc6041 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[22],stage2_7[33],stage2_6[54],stage2_5[66]}
   );
   gpc606_5 gpc6042 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[23],stage2_7[34],stage2_6[55],stage2_5[67]}
   );
   gpc606_5 gpc6043 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[24],stage2_7[35],stage2_6[56],stage2_5[68]}
   );
   gpc606_5 gpc6044 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[25],stage2_7[36],stage2_6[57],stage2_5[69]}
   );
   gpc606_5 gpc6045 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[26],stage2_7[37],stage2_6[58],stage2_5[70]}
   );
   gpc606_5 gpc6046 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[27],stage2_7[38],stage2_6[59],stage2_5[71]}
   );
   gpc606_5 gpc6047 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[28],stage2_7[39],stage2_6[60],stage2_5[72]}
   );
   gpc606_5 gpc6048 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[29],stage2_7[40],stage2_6[61],stage2_5[73]}
   );
   gpc606_5 gpc6049 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[30],stage2_7[41],stage2_6[62],stage2_5[74]}
   );
   gpc606_5 gpc6050 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[31],stage2_7[42],stage2_6[63],stage2_5[75]}
   );
   gpc606_5 gpc6051 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[32],stage2_7[43],stage2_6[64],stage2_5[76]}
   );
   gpc606_5 gpc6052 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[33],stage2_7[44],stage2_6[65],stage2_5[77]}
   );
   gpc606_5 gpc6053 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[34],stage2_7[45],stage2_6[66],stage2_5[78]}
   );
   gpc606_5 gpc6054 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[35],stage2_7[46],stage2_6[67],stage2_5[79]}
   );
   gpc606_5 gpc6055 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[36],stage2_7[47],stage2_6[68],stage2_5[80]}
   );
   gpc606_5 gpc6056 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[114], stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage2_9[19],stage2_8[37],stage2_7[48],stage2_6[69],stage2_5[81]}
   );
   gpc606_5 gpc6057 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage2_9[20],stage2_8[38],stage2_7[49],stage2_6[70],stage2_5[82]}
   );
   gpc615_5 gpc6058 (
      {stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_7[126]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[21],stage2_8[39],stage2_7[50],stage2_6[71]}
   );
   gpc615_5 gpc6059 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_7[127]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[22],stage2_8[40],stage2_7[51],stage2_6[72]}
   );
   gpc615_5 gpc6060 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124]},
      {stage1_7[128]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[23],stage2_8[41],stage2_7[52],stage2_6[73]}
   );
   gpc615_5 gpc6061 (
      {stage1_6[125], stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129]},
      {stage1_7[129]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[24],stage2_8[42],stage2_7[53],stage2_6[74]}
   );
   gpc615_5 gpc6062 (
      {stage1_6[130], stage1_6[131], stage1_6[132], stage1_6[133], stage1_6[134]},
      {stage1_7[130]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[25],stage2_8[43],stage2_7[54],stage2_6[75]}
   );
   gpc615_5 gpc6063 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[26],stage2_8[44],stage2_7[55]}
   );
   gpc615_5 gpc6064 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[27],stage2_8[45],stage2_7[56]}
   );
   gpc615_5 gpc6065 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[28],stage2_8[46],stage2_7[57]}
   );
   gpc615_5 gpc6066 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[29],stage2_8[47],stage2_7[58]}
   );
   gpc615_5 gpc6067 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[30],stage2_8[48],stage2_7[59]}
   );
   gpc615_5 gpc6068 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[31],stage2_8[49],stage2_7[60]}
   );
   gpc615_5 gpc6069 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[36]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[32],stage2_8[50],stage2_7[61]}
   );
   gpc615_5 gpc6070 (
      {stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170]},
      {stage1_8[37]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[33],stage2_8[51],stage2_7[62]}
   );
   gpc615_5 gpc6071 (
      {stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175]},
      {stage1_8[38]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[34],stage2_8[52],stage2_7[63]}
   );
   gpc615_5 gpc6072 (
      {stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_8[39]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[35],stage2_8[53],stage2_7[64]}
   );
   gpc615_5 gpc6073 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185]},
      {stage1_8[40]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[36],stage2_8[54],stage2_7[65]}
   );
   gpc615_5 gpc6074 (
      {stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190]},
      {stage1_8[41]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[37],stage2_8[55],stage2_7[66]}
   );
   gpc615_5 gpc6075 (
      {stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195]},
      {stage1_8[42]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[38],stage2_8[56],stage2_7[67]}
   );
   gpc615_5 gpc6076 (
      {stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200]},
      {stage1_8[43]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[39],stage2_8[57],stage2_7[68]}
   );
   gpc615_5 gpc6077 (
      {stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205]},
      {stage1_8[44]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[40],stage2_8[58],stage2_7[69]}
   );
   gpc615_5 gpc6078 (
      {stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_8[45]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[41],stage2_8[59],stage2_7[70]}
   );
   gpc615_5 gpc6079 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215]},
      {stage1_8[46]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[42],stage2_8[60],stage2_7[71]}
   );
   gpc615_5 gpc6080 (
      {stage1_7[216], stage1_7[217], stage1_7[218], stage1_7[219], stage1_7[220]},
      {stage1_8[47]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[43],stage2_8[61],stage2_7[72]}
   );
   gpc615_5 gpc6081 (
      {stage1_7[221], stage1_7[222], stage1_7[223], stage1_7[224], stage1_7[225]},
      {stage1_8[48]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[44],stage2_8[62],stage2_7[73]}
   );
   gpc615_5 gpc6082 (
      {stage1_7[226], stage1_7[227], stage1_7[228], stage1_7[229], stage1_7[230]},
      {stage1_8[49]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[45],stage2_8[63],stage2_7[74]}
   );
   gpc615_5 gpc6083 (
      {stage1_7[231], stage1_7[232], stage1_7[233], stage1_7[234], stage1_7[235]},
      {stage1_8[50]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[46],stage2_8[64],stage2_7[75]}
   );
   gpc615_5 gpc6084 (
      {stage1_7[236], stage1_7[237], stage1_7[238], stage1_7[239], stage1_7[240]},
      {stage1_8[51]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[26],stage2_9[47],stage2_8[65],stage2_7[76]}
   );
   gpc615_5 gpc6085 (
      {stage1_7[241], stage1_7[242], stage1_7[243], stage1_7[244], stage1_7[245]},
      {stage1_8[52]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[27],stage2_9[48],stage2_8[66],stage2_7[77]}
   );
   gpc615_5 gpc6086 (
      {stage1_7[246], stage1_7[247], stage1_7[248], stage1_7[249], stage1_7[250]},
      {stage1_8[53]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[28],stage2_9[49],stage2_8[67],stage2_7[78]}
   );
   gpc615_5 gpc6087 (
      {stage1_7[251], stage1_7[252], stage1_7[253], stage1_7[254], stage1_7[255]},
      {stage1_8[54]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[29],stage2_9[50],stage2_8[68],stage2_7[79]}
   );
   gpc615_5 gpc6088 (
      {stage1_7[256], stage1_7[257], stage1_7[258], stage1_7[259], stage1_7[260]},
      {stage1_8[55]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[30],stage2_9[51],stage2_8[69],stage2_7[80]}
   );
   gpc615_5 gpc6089 (
      {stage1_7[261], stage1_7[262], stage1_7[263], stage1_7[264], stage1_7[265]},
      {stage1_8[56]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[31],stage2_9[52],stage2_8[70],stage2_7[81]}
   );
   gpc615_5 gpc6090 (
      {stage1_7[266], stage1_7[267], stage1_7[268], stage1_7[269], stage1_7[270]},
      {stage1_8[57]},
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage2_11[27],stage2_10[32],stage2_9[53],stage2_8[71],stage2_7[82]}
   );
   gpc615_5 gpc6091 (
      {stage1_7[271], stage1_7[272], stage1_7[273], stage1_7[274], stage1_7[275]},
      {stage1_8[58]},
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage2_11[28],stage2_10[33],stage2_9[54],stage2_8[72],stage2_7[83]}
   );
   gpc615_5 gpc6092 (
      {stage1_7[276], stage1_7[277], stage1_7[278], stage1_7[279], stage1_7[280]},
      {stage1_8[59]},
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage2_11[29],stage2_10[34],stage2_9[55],stage2_8[73],stage2_7[84]}
   );
   gpc615_5 gpc6093 (
      {stage1_7[281], stage1_7[282], stage1_7[283], stage1_7[284], stage1_7[285]},
      {stage1_8[60]},
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage2_11[30],stage2_10[35],stage2_9[56],stage2_8[74],stage2_7[85]}
   );
   gpc615_5 gpc6094 (
      {stage1_7[286], stage1_7[287], stage1_7[288], stage1_7[289], stage1_7[290]},
      {stage1_8[61]},
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage2_11[31],stage2_10[36],stage2_9[57],stage2_8[75],stage2_7[86]}
   );
   gpc615_5 gpc6095 (
      {stage1_7[291], stage1_7[292], stage1_7[293], stage1_7[294], stage1_7[295]},
      {stage1_8[62]},
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage2_11[32],stage2_10[37],stage2_9[58],stage2_8[76],stage2_7[87]}
   );
   gpc615_5 gpc6096 (
      {stage1_7[296], stage1_7[297], stage1_7[298], stage1_7[299], stage1_7[300]},
      {stage1_8[63]},
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage2_11[33],stage2_10[38],stage2_9[59],stage2_8[77],stage2_7[88]}
   );
   gpc615_5 gpc6097 (
      {stage1_7[301], stage1_7[302], stage1_7[303], stage1_7[304], stage1_7[305]},
      {stage1_8[64]},
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage2_11[34],stage2_10[39],stage2_9[60],stage2_8[78],stage2_7[89]}
   );
   gpc615_5 gpc6098 (
      {stage1_7[306], stage1_7[307], stage1_7[308], stage1_7[309], stage1_7[310]},
      {stage1_8[65]},
      {stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213], stage1_9[214], stage1_9[215]},
      {stage2_11[35],stage2_10[40],stage2_9[61],stage2_8[79],stage2_7[90]}
   );
   gpc615_5 gpc6099 (
      {stage1_7[311], stage1_7[312], stage1_7[313], stage1_7[314], stage1_7[315]},
      {stage1_8[66]},
      {stage1_9[216], stage1_9[217], stage1_9[218], stage1_9[219], stage1_9[220], stage1_9[221]},
      {stage2_11[36],stage2_10[41],stage2_9[62],stage2_8[80],stage2_7[91]}
   );
   gpc615_5 gpc6100 (
      {stage1_7[316], stage1_7[317], stage1_7[318], stage1_7[319], stage1_7[320]},
      {stage1_8[67]},
      {stage1_9[222], stage1_9[223], stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227]},
      {stage2_11[37],stage2_10[42],stage2_9[63],stage2_8[81],stage2_7[92]}
   );
   gpc615_5 gpc6101 (
      {stage1_7[321], stage1_7[322], stage1_7[323], stage1_7[324], stage1_7[325]},
      {stage1_8[68]},
      {stage1_9[228], stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage2_11[38],stage2_10[43],stage2_9[64],stage2_8[82],stage2_7[93]}
   );
   gpc615_5 gpc6102 (
      {stage1_7[326], stage1_7[327], stage1_7[328], stage1_7[329], stage1_7[330]},
      {stage1_8[69]},
      {stage1_9[234], stage1_9[235], stage1_9[236], stage1_9[237], stage1_9[238], stage1_9[239]},
      {stage2_11[39],stage2_10[44],stage2_9[65],stage2_8[83],stage2_7[94]}
   );
   gpc615_5 gpc6103 (
      {stage1_7[331], stage1_7[332], stage1_7[333], stage1_7[334], stage1_7[335]},
      {stage1_8[70]},
      {stage1_9[240], stage1_9[241], stage1_9[242], stage1_9[243], stage1_9[244], stage1_9[245]},
      {stage2_11[40],stage2_10[45],stage2_9[66],stage2_8[84],stage2_7[95]}
   );
   gpc615_5 gpc6104 (
      {stage1_7[336], stage1_7[337], stage1_7[338], stage1_7[339], 1'b0},
      {stage1_8[71]},
      {stage1_9[246], stage1_9[247], stage1_9[248], stage1_9[249], stage1_9[250], stage1_9[251]},
      {stage2_11[41],stage2_10[46],stage2_9[67],stage2_8[85],stage2_7[96]}
   );
   gpc606_5 gpc6105 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[42],stage2_10[47],stage2_9[68],stage2_8[86]}
   );
   gpc606_5 gpc6106 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[43],stage2_10[48],stage2_9[69],stage2_8[87]}
   );
   gpc606_5 gpc6107 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[44],stage2_10[49],stage2_9[70],stage2_8[88]}
   );
   gpc606_5 gpc6108 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[45],stage2_10[50],stage2_9[71],stage2_8[89]}
   );
   gpc606_5 gpc6109 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[46],stage2_10[51],stage2_9[72],stage2_8[90]}
   );
   gpc606_5 gpc6110 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[47],stage2_10[52],stage2_9[73],stage2_8[91]}
   );
   gpc606_5 gpc6111 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[48],stage2_10[53],stage2_9[74],stage2_8[92]}
   );
   gpc606_5 gpc6112 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[49],stage2_10[54],stage2_9[75],stage2_8[93]}
   );
   gpc606_5 gpc6113 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[50],stage2_10[55],stage2_9[76],stage2_8[94]}
   );
   gpc606_5 gpc6114 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[51],stage2_10[56],stage2_9[77],stage2_8[95]}
   );
   gpc606_5 gpc6115 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[52],stage2_10[57],stage2_9[78],stage2_8[96]}
   );
   gpc606_5 gpc6116 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[53],stage2_10[58],stage2_9[79],stage2_8[97]}
   );
   gpc606_5 gpc6117 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[54],stage2_10[59],stage2_9[80],stage2_8[98]}
   );
   gpc606_5 gpc6118 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[55],stage2_10[60],stage2_9[81],stage2_8[99]}
   );
   gpc606_5 gpc6119 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[56],stage2_10[61],stage2_9[82],stage2_8[100]}
   );
   gpc606_5 gpc6120 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[57],stage2_10[62],stage2_9[83],stage2_8[101]}
   );
   gpc606_5 gpc6121 (
      {stage1_9[252], stage1_9[253], stage1_9[254], stage1_9[255], stage1_9[256], stage1_9[257]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[16],stage2_11[58],stage2_10[63],stage2_9[84]}
   );
   gpc606_5 gpc6122 (
      {stage1_9[258], stage1_9[259], stage1_9[260], stage1_9[261], stage1_9[262], stage1_9[263]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[17],stage2_11[59],stage2_10[64],stage2_9[85]}
   );
   gpc606_5 gpc6123 (
      {stage1_9[264], stage1_9[265], stage1_9[266], stage1_9[267], stage1_9[268], stage1_9[269]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[18],stage2_11[60],stage2_10[65],stage2_9[86]}
   );
   gpc606_5 gpc6124 (
      {stage1_9[270], stage1_9[271], stage1_9[272], stage1_9[273], stage1_9[274], stage1_9[275]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[19],stage2_11[61],stage2_10[66],stage2_9[87]}
   );
   gpc606_5 gpc6125 (
      {stage1_9[276], stage1_9[277], stage1_9[278], stage1_9[279], stage1_9[280], stage1_9[281]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[20],stage2_11[62],stage2_10[67],stage2_9[88]}
   );
   gpc606_5 gpc6126 (
      {stage1_9[282], stage1_9[283], stage1_9[284], stage1_9[285], stage1_9[286], stage1_9[287]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[21],stage2_11[63],stage2_10[68],stage2_9[89]}
   );
   gpc606_5 gpc6127 (
      {stage1_9[288], stage1_9[289], stage1_9[290], stage1_9[291], stage1_9[292], stage1_9[293]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[22],stage2_11[64],stage2_10[69],stage2_9[90]}
   );
   gpc606_5 gpc6128 (
      {stage1_9[294], stage1_9[295], stage1_9[296], stage1_9[297], stage1_9[298], stage1_9[299]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[23],stage2_11[65],stage2_10[70],stage2_9[91]}
   );
   gpc606_5 gpc6129 (
      {stage1_9[300], stage1_9[301], stage1_9[302], stage1_9[303], stage1_9[304], stage1_9[305]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[24],stage2_11[66],stage2_10[71],stage2_9[92]}
   );
   gpc606_5 gpc6130 (
      {stage1_9[306], stage1_9[307], stage1_9[308], stage1_9[309], stage1_9[310], stage1_9[311]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[25],stage2_11[67],stage2_10[72],stage2_9[93]}
   );
   gpc606_5 gpc6131 (
      {stage1_9[312], stage1_9[313], stage1_9[314], stage1_9[315], stage1_9[316], stage1_9[317]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[26],stage2_11[68],stage2_10[73],stage2_9[94]}
   );
   gpc606_5 gpc6132 (
      {stage1_9[318], stage1_9[319], stage1_9[320], stage1_9[321], stage1_9[322], stage1_9[323]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[27],stage2_11[69],stage2_10[74],stage2_9[95]}
   );
   gpc606_5 gpc6133 (
      {stage1_9[324], stage1_9[325], stage1_9[326], stage1_9[327], stage1_9[328], stage1_9[329]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[28],stage2_11[70],stage2_10[75],stage2_9[96]}
   );
   gpc606_5 gpc6134 (
      {stage1_9[330], stage1_9[331], stage1_9[332], stage1_9[333], stage1_9[334], stage1_9[335]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[29],stage2_11[71],stage2_10[76],stage2_9[97]}
   );
   gpc606_5 gpc6135 (
      {stage1_9[336], stage1_9[337], stage1_9[338], stage1_9[339], stage1_9[340], stage1_9[341]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[30],stage2_11[72],stage2_10[77],stage2_9[98]}
   );
   gpc606_5 gpc6136 (
      {stage1_9[342], stage1_9[343], stage1_9[344], stage1_9[345], stage1_9[346], stage1_9[347]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[31],stage2_11[73],stage2_10[78],stage2_9[99]}
   );
   gpc606_5 gpc6137 (
      {stage1_9[348], stage1_9[349], stage1_9[350], stage1_9[351], stage1_9[352], stage1_9[353]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[32],stage2_11[74],stage2_10[79],stage2_9[100]}
   );
   gpc606_5 gpc6138 (
      {stage1_9[354], stage1_9[355], stage1_9[356], stage1_9[357], stage1_9[358], stage1_9[359]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[33],stage2_11[75],stage2_10[80],stage2_9[101]}
   );
   gpc615_5 gpc6139 (
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_11[108]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[34],stage2_11[76],stage2_10[81]}
   );
   gpc1163_5 gpc6140 (
      {stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_13[0]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[19],stage2_12[35],stage2_11[77]}
   );
   gpc1163_5 gpc6141 (
      {stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage1_13[1]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[20],stage2_12[36],stage2_11[78]}
   );
   gpc1163_5 gpc6142 (
      {stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage1_13[2]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[21],stage2_12[37],stage2_11[79]}
   );
   gpc1163_5 gpc6143 (
      {stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage1_13[3]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[22],stage2_12[38],stage2_11[80]}
   );
   gpc1163_5 gpc6144 (
      {stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage1_13[4]},
      {stage1_14[4]},
      {stage2_15[4],stage2_14[5],stage2_13[23],stage2_12[39],stage2_11[81]}
   );
   gpc1163_5 gpc6145 (
      {stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[5]},
      {stage1_14[5]},
      {stage2_15[5],stage2_14[6],stage2_13[24],stage2_12[40],stage2_11[82]}
   );
   gpc1163_5 gpc6146 (
      {stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_13[6]},
      {stage1_14[6]},
      {stage2_15[6],stage2_14[7],stage2_13[25],stage2_12[41],stage2_11[83]}
   );
   gpc1163_5 gpc6147 (
      {stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_13[7]},
      {stage1_14[7]},
      {stage2_15[7],stage2_14[8],stage2_13[26],stage2_12[42],stage2_11[84]}
   );
   gpc1163_5 gpc6148 (
      {stage1_11[133], stage1_11[134], stage1_11[135]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[8]},
      {stage1_14[8]},
      {stage2_15[8],stage2_14[9],stage2_13[27],stage2_12[43],stage2_11[85]}
   );
   gpc1163_5 gpc6149 (
      {stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_13[9]},
      {stage1_14[9]},
      {stage2_15[9],stage2_14[10],stage2_13[28],stage2_12[44],stage2_11[86]}
   );
   gpc1163_5 gpc6150 (
      {stage1_11[139], stage1_11[140], stage1_11[141]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage1_13[10]},
      {stage1_14[10]},
      {stage2_15[10],stage2_14[11],stage2_13[29],stage2_12[45],stage2_11[87]}
   );
   gpc1163_5 gpc6151 (
      {stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage1_13[11]},
      {stage1_14[11]},
      {stage2_15[11],stage2_14[12],stage2_13[30],stage2_12[46],stage2_11[88]}
   );
   gpc1163_5 gpc6152 (
      {stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage1_13[12]},
      {stage1_14[12]},
      {stage2_15[12],stage2_14[13],stage2_13[31],stage2_12[47],stage2_11[89]}
   );
   gpc1163_5 gpc6153 (
      {stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[13]},
      {stage1_14[13]},
      {stage2_15[13],stage2_14[14],stage2_13[32],stage2_12[48],stage2_11[90]}
   );
   gpc1163_5 gpc6154 (
      {stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage1_13[14]},
      {stage1_14[14]},
      {stage2_15[14],stage2_14[15],stage2_13[33],stage2_12[49],stage2_11[91]}
   );
   gpc1163_5 gpc6155 (
      {stage1_11[154], stage1_11[155], stage1_11[156]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_13[15]},
      {stage1_14[15]},
      {stage2_15[15],stage2_14[16],stage2_13[34],stage2_12[50],stage2_11[92]}
   );
   gpc1163_5 gpc6156 (
      {stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage1_13[16]},
      {stage1_14[16]},
      {stage2_15[16],stage2_14[17],stage2_13[35],stage2_12[51],stage2_11[93]}
   );
   gpc1163_5 gpc6157 (
      {stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_13[17]},
      {stage1_14[17]},
      {stage2_15[17],stage2_14[18],stage2_13[36],stage2_12[52],stage2_11[94]}
   );
   gpc1163_5 gpc6158 (
      {stage1_11[163], stage1_11[164], stage1_11[165]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[18]},
      {stage1_14[18]},
      {stage2_15[18],stage2_14[19],stage2_13[37],stage2_12[53],stage2_11[95]}
   );
   gpc1163_5 gpc6159 (
      {stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_13[19]},
      {stage1_14[19]},
      {stage2_15[19],stage2_14[20],stage2_13[38],stage2_12[54],stage2_11[96]}
   );
   gpc1163_5 gpc6160 (
      {stage1_11[169], stage1_11[170], stage1_11[171]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_13[20]},
      {stage1_14[20]},
      {stage2_15[20],stage2_14[21],stage2_13[39],stage2_12[55],stage2_11[97]}
   );
   gpc615_5 gpc6161 (
      {stage1_11[172], stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176]},
      {stage1_12[132]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[21],stage2_14[22],stage2_13[40],stage2_12[56],stage2_11[98]}
   );
   gpc615_5 gpc6162 (
      {stage1_11[177], stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181]},
      {stage1_12[133]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[22],stage2_14[23],stage2_13[41],stage2_12[57],stage2_11[99]}
   );
   gpc615_5 gpc6163 (
      {stage1_11[182], stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186]},
      {stage1_12[134]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[23],stage2_14[24],stage2_13[42],stage2_12[58],stage2_11[100]}
   );
   gpc615_5 gpc6164 (
      {stage1_11[187], stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191]},
      {stage1_12[135]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[24],stage2_14[25],stage2_13[43],stage2_12[59],stage2_11[101]}
   );
   gpc615_5 gpc6165 (
      {stage1_11[192], stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196]},
      {stage1_12[136]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[25],stage2_14[26],stage2_13[44],stage2_12[60],stage2_11[102]}
   );
   gpc615_5 gpc6166 (
      {stage1_11[197], stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201]},
      {stage1_12[137]},
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage2_15[26],stage2_14[27],stage2_13[45],stage2_12[61],stage2_11[103]}
   );
   gpc615_5 gpc6167 (
      {stage1_11[202], stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206]},
      {stage1_12[138]},
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage2_15[27],stage2_14[28],stage2_13[46],stage2_12[62],stage2_11[104]}
   );
   gpc615_5 gpc6168 (
      {stage1_11[207], stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211]},
      {stage1_12[139]},
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage2_15[28],stage2_14[29],stage2_13[47],stage2_12[63],stage2_11[105]}
   );
   gpc615_5 gpc6169 (
      {stage1_11[212], stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216]},
      {stage1_12[140]},
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage2_15[29],stage2_14[30],stage2_13[48],stage2_12[64],stage2_11[106]}
   );
   gpc615_5 gpc6170 (
      {stage1_11[217], stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221]},
      {stage1_12[141]},
      {stage1_13[75], stage1_13[76], stage1_13[77], stage1_13[78], stage1_13[79], stage1_13[80]},
      {stage2_15[30],stage2_14[31],stage2_13[49],stage2_12[65],stage2_11[107]}
   );
   gpc615_5 gpc6171 (
      {stage1_11[222], stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226]},
      {stage1_12[142]},
      {stage1_13[81], stage1_13[82], stage1_13[83], stage1_13[84], stage1_13[85], stage1_13[86]},
      {stage2_15[31],stage2_14[32],stage2_13[50],stage2_12[66],stage2_11[108]}
   );
   gpc615_5 gpc6172 (
      {stage1_11[227], stage1_11[228], stage1_11[229], stage1_11[230], stage1_11[231]},
      {stage1_12[143]},
      {stage1_13[87], stage1_13[88], stage1_13[89], stage1_13[90], stage1_13[91], stage1_13[92]},
      {stage2_15[32],stage2_14[33],stage2_13[51],stage2_12[67],stage2_11[109]}
   );
   gpc615_5 gpc6173 (
      {stage1_11[232], stage1_11[233], stage1_11[234], stage1_11[235], stage1_11[236]},
      {stage1_12[144]},
      {stage1_13[93], stage1_13[94], stage1_13[95], stage1_13[96], stage1_13[97], stage1_13[98]},
      {stage2_15[33],stage2_14[34],stage2_13[52],stage2_12[68],stage2_11[110]}
   );
   gpc615_5 gpc6174 (
      {stage1_11[237], stage1_11[238], stage1_11[239], stage1_11[240], stage1_11[241]},
      {stage1_12[145]},
      {stage1_13[99], stage1_13[100], stage1_13[101], stage1_13[102], stage1_13[103], stage1_13[104]},
      {stage2_15[34],stage2_14[35],stage2_13[53],stage2_12[69],stage2_11[111]}
   );
   gpc615_5 gpc6175 (
      {stage1_11[242], stage1_11[243], stage1_11[244], stage1_11[245], stage1_11[246]},
      {stage1_12[146]},
      {stage1_13[105], stage1_13[106], stage1_13[107], stage1_13[108], stage1_13[109], stage1_13[110]},
      {stage2_15[35],stage2_14[36],stage2_13[54],stage2_12[70],stage2_11[112]}
   );
   gpc615_5 gpc6176 (
      {stage1_11[247], stage1_11[248], stage1_11[249], stage1_11[250], stage1_11[251]},
      {stage1_12[147]},
      {stage1_13[111], stage1_13[112], stage1_13[113], stage1_13[114], stage1_13[115], stage1_13[116]},
      {stage2_15[36],stage2_14[37],stage2_13[55],stage2_12[71],stage2_11[113]}
   );
   gpc615_5 gpc6177 (
      {stage1_11[252], stage1_11[253], stage1_11[254], stage1_11[255], stage1_11[256]},
      {stage1_12[148]},
      {stage1_13[117], stage1_13[118], stage1_13[119], stage1_13[120], stage1_13[121], stage1_13[122]},
      {stage2_15[37],stage2_14[38],stage2_13[56],stage2_12[72],stage2_11[114]}
   );
   gpc615_5 gpc6178 (
      {stage1_11[257], stage1_11[258], stage1_11[259], stage1_11[260], stage1_11[261]},
      {stage1_12[149]},
      {stage1_13[123], stage1_13[124], stage1_13[125], stage1_13[126], stage1_13[127], stage1_13[128]},
      {stage2_15[38],stage2_14[39],stage2_13[57],stage2_12[73],stage2_11[115]}
   );
   gpc615_5 gpc6179 (
      {stage1_11[262], stage1_11[263], stage1_11[264], stage1_11[265], stage1_11[266]},
      {stage1_12[150]},
      {stage1_13[129], stage1_13[130], stage1_13[131], stage1_13[132], stage1_13[133], stage1_13[134]},
      {stage2_15[39],stage2_14[40],stage2_13[58],stage2_12[74],stage2_11[116]}
   );
   gpc615_5 gpc6180 (
      {stage1_11[267], stage1_11[268], stage1_11[269], stage1_11[270], stage1_11[271]},
      {stage1_12[151]},
      {stage1_13[135], stage1_13[136], stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140]},
      {stage2_15[40],stage2_14[41],stage2_13[59],stage2_12[75],stage2_11[117]}
   );
   gpc615_5 gpc6181 (
      {stage1_11[272], stage1_11[273], stage1_11[274], stage1_11[275], stage1_11[276]},
      {stage1_12[152]},
      {stage1_13[141], stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage2_15[41],stage2_14[42],stage2_13[60],stage2_12[76],stage2_11[118]}
   );
   gpc615_5 gpc6182 (
      {stage1_11[277], stage1_11[278], stage1_11[279], stage1_11[280], stage1_11[281]},
      {stage1_12[153]},
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151], stage1_13[152]},
      {stage2_15[42],stage2_14[43],stage2_13[61],stage2_12[77],stage2_11[119]}
   );
   gpc615_5 gpc6183 (
      {stage1_11[282], stage1_11[283], stage1_11[284], stage1_11[285], stage1_11[286]},
      {stage1_12[154]},
      {stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158]},
      {stage2_15[43],stage2_14[44],stage2_13[62],stage2_12[78],stage2_11[120]}
   );
   gpc615_5 gpc6184 (
      {stage1_11[287], stage1_11[288], stage1_11[289], stage1_11[290], stage1_11[291]},
      {stage1_12[155]},
      {stage1_13[159], stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage2_15[44],stage2_14[45],stage2_13[63],stage2_12[79],stage2_11[121]}
   );
   gpc615_5 gpc6185 (
      {stage1_11[292], stage1_11[293], stage1_11[294], stage1_11[295], stage1_11[296]},
      {stage1_12[156]},
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170]},
      {stage2_15[45],stage2_14[46],stage2_13[64],stage2_12[80],stage2_11[122]}
   );
   gpc615_5 gpc6186 (
      {stage1_11[297], stage1_11[298], stage1_11[299], stage1_11[300], stage1_11[301]},
      {stage1_12[157]},
      {stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage2_15[46],stage2_14[47],stage2_13[65],stage2_12[81],stage2_11[123]}
   );
   gpc615_5 gpc6187 (
      {stage1_11[302], stage1_11[303], stage1_11[304], stage1_11[305], stage1_11[306]},
      {stage1_12[158]},
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181], stage1_13[182]},
      {stage2_15[47],stage2_14[48],stage2_13[66],stage2_12[82],stage2_11[124]}
   );
   gpc606_5 gpc6188 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26]},
      {stage2_16[0],stage2_15[48],stage2_14[49],stage2_13[67],stage2_12[83]}
   );
   gpc606_5 gpc6189 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31], stage1_14[32]},
      {stage2_16[1],stage2_15[49],stage2_14[50],stage2_13[68],stage2_12[84]}
   );
   gpc606_5 gpc6190 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37], stage1_14[38]},
      {stage2_16[2],stage2_15[50],stage2_14[51],stage2_13[69],stage2_12[85]}
   );
   gpc1163_5 gpc6191 (
      {stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[0],stage2_16[3],stage2_15[51],stage2_14[52]}
   );
   gpc1163_5 gpc6192 (
      {stage1_14[42], stage1_14[43], stage1_14[44]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[1]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[1],stage2_16[4],stage2_15[52],stage2_14[53]}
   );
   gpc1163_5 gpc6193 (
      {stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[2]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[2],stage2_16[5],stage2_15[53],stage2_14[54]}
   );
   gpc1163_5 gpc6194 (
      {stage1_14[48], stage1_14[49], stage1_14[50]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[3]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[3],stage2_16[6],stage2_15[54],stage2_14[55]}
   );
   gpc1163_5 gpc6195 (
      {stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[4]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[4],stage2_16[7],stage2_15[55],stage2_14[56]}
   );
   gpc1163_5 gpc6196 (
      {stage1_14[54], stage1_14[55], stage1_14[56]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[5]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[5],stage2_16[8],stage2_15[56],stage2_14[57]}
   );
   gpc1163_5 gpc6197 (
      {stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage1_16[6]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[6],stage2_16[9],stage2_15[57],stage2_14[58]}
   );
   gpc1163_5 gpc6198 (
      {stage1_14[60], stage1_14[61], stage1_14[62]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[7]},
      {stage1_17[7]},
      {stage2_18[7],stage2_17[7],stage2_16[10],stage2_15[58],stage2_14[59]}
   );
   gpc1163_5 gpc6199 (
      {stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[8]},
      {stage1_17[8]},
      {stage2_18[8],stage2_17[8],stage2_16[11],stage2_15[59],stage2_14[60]}
   );
   gpc1163_5 gpc6200 (
      {stage1_14[66], stage1_14[67], stage1_14[68]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage1_16[9]},
      {stage1_17[9]},
      {stage2_18[9],stage2_17[9],stage2_16[12],stage2_15[60],stage2_14[61]}
   );
   gpc1163_5 gpc6201 (
      {stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_16[10]},
      {stage1_17[10]},
      {stage2_18[10],stage2_17[10],stage2_16[13],stage2_15[61],stage2_14[62]}
   );
   gpc1163_5 gpc6202 (
      {stage1_14[72], stage1_14[73], stage1_14[74]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage1_16[11]},
      {stage1_17[11]},
      {stage2_18[11],stage2_17[11],stage2_16[14],stage2_15[62],stage2_14[63]}
   );
   gpc1163_5 gpc6203 (
      {stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[12]},
      {stage1_17[12]},
      {stage2_18[12],stage2_17[12],stage2_16[15],stage2_15[63],stage2_14[64]}
   );
   gpc1163_5 gpc6204 (
      {stage1_14[78], stage1_14[79], stage1_14[80]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[13]},
      {stage1_17[13]},
      {stage2_18[13],stage2_17[13],stage2_16[16],stage2_15[64],stage2_14[65]}
   );
   gpc1163_5 gpc6205 (
      {stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage1_16[14]},
      {stage1_17[14]},
      {stage2_18[14],stage2_17[14],stage2_16[17],stage2_15[65],stage2_14[66]}
   );
   gpc1163_5 gpc6206 (
      {stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage1_16[15]},
      {stage1_17[15]},
      {stage2_18[15],stage2_17[15],stage2_16[18],stage2_15[66],stage2_14[67]}
   );
   gpc1163_5 gpc6207 (
      {stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage1_16[16]},
      {stage1_17[16]},
      {stage2_18[16],stage2_17[16],stage2_16[19],stage2_15[67],stage2_14[68]}
   );
   gpc1163_5 gpc6208 (
      {stage1_14[90], stage1_14[91], stage1_14[92]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[17]},
      {stage1_17[17]},
      {stage2_18[17],stage2_17[17],stage2_16[20],stage2_15[68],stage2_14[69]}
   );
   gpc1163_5 gpc6209 (
      {stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage1_16[18]},
      {stage1_17[18]},
      {stage2_18[18],stage2_17[18],stage2_16[21],stage2_15[69],stage2_14[70]}
   );
   gpc1163_5 gpc6210 (
      {stage1_14[96], stage1_14[97], stage1_14[98]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage1_16[19]},
      {stage1_17[19]},
      {stage2_18[19],stage2_17[19],stage2_16[22],stage2_15[70],stage2_14[71]}
   );
   gpc1163_5 gpc6211 (
      {stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage1_16[20]},
      {stage1_17[20]},
      {stage2_18[20],stage2_17[20],stage2_16[23],stage2_15[71],stage2_14[72]}
   );
   gpc1163_5 gpc6212 (
      {stage1_14[102], stage1_14[103], stage1_14[104]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage1_16[21]},
      {stage1_17[21]},
      {stage2_18[21],stage2_17[21],stage2_16[24],stage2_15[72],stage2_14[73]}
   );
   gpc1163_5 gpc6213 (
      {stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage1_16[22]},
      {stage1_17[22]},
      {stage2_18[22],stage2_17[22],stage2_16[25],stage2_15[73],stage2_14[74]}
   );
   gpc1163_5 gpc6214 (
      {stage1_14[108], stage1_14[109], stage1_14[110]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage1_16[23]},
      {stage1_17[23]},
      {stage2_18[23],stage2_17[23],stage2_16[26],stage2_15[74],stage2_14[75]}
   );
   gpc1163_5 gpc6215 (
      {stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage1_16[24]},
      {stage1_17[24]},
      {stage2_18[24],stage2_17[24],stage2_16[27],stage2_15[75],stage2_14[76]}
   );
   gpc1163_5 gpc6216 (
      {stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage1_16[25]},
      {stage1_17[25]},
      {stage2_18[25],stage2_17[25],stage2_16[28],stage2_15[76],stage2_14[77]}
   );
   gpc1163_5 gpc6217 (
      {stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[26]},
      {stage1_17[26]},
      {stage2_18[26],stage2_17[26],stage2_16[29],stage2_15[77],stage2_14[78]}
   );
   gpc1163_5 gpc6218 (
      {stage1_14[120], stage1_14[121], stage1_14[122]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage1_16[27]},
      {stage1_17[27]},
      {stage2_18[27],stage2_17[27],stage2_16[30],stage2_15[78],stage2_14[79]}
   );
   gpc1163_5 gpc6219 (
      {stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage1_16[28]},
      {stage1_17[28]},
      {stage2_18[28],stage2_17[28],stage2_16[31],stage2_15[79],stage2_14[80]}
   );
   gpc1163_5 gpc6220 (
      {stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage1_16[29]},
      {stage1_17[29]},
      {stage2_18[29],stage2_17[29],stage2_16[32],stage2_15[80],stage2_14[81]}
   );
   gpc1163_5 gpc6221 (
      {stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage1_16[30]},
      {stage1_17[30]},
      {stage2_18[30],stage2_17[30],stage2_16[33],stage2_15[81],stage2_14[82]}
   );
   gpc1163_5 gpc6222 (
      {stage1_14[132], stage1_14[133], stage1_14[134]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[31]},
      {stage1_17[31]},
      {stage2_18[31],stage2_17[31],stage2_16[34],stage2_15[82],stage2_14[83]}
   );
   gpc606_5 gpc6223 (
      {stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140]},
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage2_18[32],stage2_17[32],stage2_16[35],stage2_15[83],stage2_14[84]}
   );
   gpc606_5 gpc6224 (
      {stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage2_18[33],stage2_17[33],stage2_16[36],stage2_15[84],stage2_14[85]}
   );
   gpc606_5 gpc6225 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152]},
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage2_18[34],stage2_17[34],stage2_16[37],stage2_15[85],stage2_14[86]}
   );
   gpc606_5 gpc6226 (
      {stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage2_18[35],stage2_17[35],stage2_16[38],stage2_15[86],stage2_14[87]}
   );
   gpc606_5 gpc6227 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163], stage1_14[164]},
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage2_18[36],stage2_17[36],stage2_16[39],stage2_15[87],stage2_14[88]}
   );
   gpc606_5 gpc6228 (
      {stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170]},
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage2_18[37],stage2_17[37],stage2_16[40],stage2_15[88],stage2_14[89]}
   );
   gpc615_5 gpc6229 (
      {stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_15[192]},
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage2_18[38],stage2_17[38],stage2_16[41],stage2_15[89],stage2_14[90]}
   );
   gpc615_5 gpc6230 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180]},
      {stage1_15[193]},
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage2_18[39],stage2_17[39],stage2_16[42],stage2_15[90],stage2_14[91]}
   );
   gpc615_5 gpc6231 (
      {stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage1_15[194]},
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage2_18[40],stage2_17[40],stage2_16[43],stage2_15[91],stage2_14[92]}
   );
   gpc615_5 gpc6232 (
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190]},
      {stage1_15[195]},
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage2_18[41],stage2_17[41],stage2_16[44],stage2_15[92],stage2_14[93]}
   );
   gpc615_5 gpc6233 (
      {stage1_14[191], stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195]},
      {stage1_15[196]},
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage2_18[42],stage2_17[42],stage2_16[45],stage2_15[93],stage2_14[94]}
   );
   gpc615_5 gpc6234 (
      {stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200]},
      {stage1_15[197]},
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage2_18[43],stage2_17[43],stage2_16[46],stage2_15[94],stage2_14[95]}
   );
   gpc615_5 gpc6235 (
      {stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_15[198]},
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage2_18[44],stage2_17[44],stage2_16[47],stage2_15[95],stage2_14[96]}
   );
   gpc615_5 gpc6236 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[199]},
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage2_18[45],stage2_17[45],stage2_16[48],stage2_15[96],stage2_14[97]}
   );
   gpc615_5 gpc6237 (
      {stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage1_15[200]},
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage2_18[46],stage2_17[46],stage2_16[49],stage2_15[97],stage2_14[98]}
   );
   gpc615_5 gpc6238 (
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220]},
      {stage1_15[201]},
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage2_18[47],stage2_17[47],stage2_16[50],stage2_15[98],stage2_14[99]}
   );
   gpc615_5 gpc6239 (
      {stage1_14[221], stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225]},
      {stage1_15[202]},
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage2_18[48],stage2_17[48],stage2_16[51],stage2_15[99],stage2_14[100]}
   );
   gpc615_5 gpc6240 (
      {stage1_14[226], stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230]},
      {stage1_15[203]},
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage2_18[49],stage2_17[49],stage2_16[52],stage2_15[100],stage2_14[101]}
   );
   gpc615_5 gpc6241 (
      {stage1_14[231], stage1_14[232], stage1_14[233], stage1_14[234], stage1_14[235]},
      {stage1_15[204]},
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage2_18[50],stage2_17[50],stage2_16[53],stage2_15[101],stage2_14[102]}
   );
   gpc615_5 gpc6242 (
      {stage1_14[236], stage1_14[237], stage1_14[238], stage1_14[239], stage1_14[240]},
      {stage1_15[205]},
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage2_18[51],stage2_17[51],stage2_16[54],stage2_15[102],stage2_14[103]}
   );
   gpc615_5 gpc6243 (
      {stage1_14[241], stage1_14[242], stage1_14[243], stage1_14[244], stage1_14[245]},
      {stage1_15[206]},
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage2_18[52],stage2_17[52],stage2_16[55],stage2_15[103],stage2_14[104]}
   );
   gpc1406_5 gpc6244 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211], stage1_15[212]},
      {stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[53],stage2_17[53],stage2_16[56],stage2_15[104]}
   );
   gpc1406_5 gpc6245 (
      {stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216], stage1_15[217], stage1_15[218]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39]},
      {stage1_18[1]},
      {stage2_19[1],stage2_18[54],stage2_17[54],stage2_16[57],stage2_15[105]}
   );
   gpc606_5 gpc6246 (
      {stage1_15[219], stage1_15[220], stage1_15[221], stage1_15[222], stage1_15[223], stage1_15[224]},
      {stage1_17[40], stage1_17[41], stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45]},
      {stage2_19[2],stage2_18[55],stage2_17[55],stage2_16[58],stage2_15[106]}
   );
   gpc606_5 gpc6247 (
      {stage1_15[225], stage1_15[226], stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230]},
      {stage1_17[46], stage1_17[47], stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51]},
      {stage2_19[3],stage2_18[56],stage2_17[56],stage2_16[59],stage2_15[107]}
   );
   gpc606_5 gpc6248 (
      {stage1_15[231], stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_17[52], stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage2_19[4],stage2_18[57],stage2_17[57],stage2_16[60],stage2_15[108]}
   );
   gpc606_5 gpc6249 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241], stage1_15[242]},
      {stage1_17[58], stage1_17[59], stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63]},
      {stage2_19[5],stage2_18[58],stage2_17[58],stage2_16[61],stage2_15[109]}
   );
   gpc606_5 gpc6250 (
      {stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246], stage1_15[247], stage1_15[248]},
      {stage1_17[64], stage1_17[65], stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69]},
      {stage2_19[6],stage2_18[59],stage2_17[59],stage2_16[62],stage2_15[110]}
   );
   gpc606_5 gpc6251 (
      {stage1_15[249], stage1_15[250], stage1_15[251], stage1_15[252], stage1_15[253], stage1_15[254]},
      {stage1_17[70], stage1_17[71], stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75]},
      {stage2_19[7],stage2_18[60],stage2_17[60],stage2_16[63],stage2_15[111]}
   );
   gpc606_5 gpc6252 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6], stage1_18[7]},
      {stage2_20[0],stage2_19[8],stage2_18[61],stage2_17[61],stage2_16[64]}
   );
   gpc606_5 gpc6253 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12], stage1_18[13]},
      {stage2_20[1],stage2_19[9],stage2_18[62],stage2_17[62],stage2_16[65]}
   );
   gpc606_5 gpc6254 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18], stage1_18[19]},
      {stage2_20[2],stage2_19[10],stage2_18[63],stage2_17[63],stage2_16[66]}
   );
   gpc606_5 gpc6255 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180], stage1_16[181]},
      {stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25]},
      {stage2_20[3],stage2_19[11],stage2_18[64],stage2_17[64],stage2_16[67]}
   );
   gpc606_5 gpc6256 (
      {stage1_17[76], stage1_17[77], stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[4],stage2_19[12],stage2_18[65],stage2_17[65]}
   );
   gpc606_5 gpc6257 (
      {stage1_17[82], stage1_17[83], stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[5],stage2_19[13],stage2_18[66],stage2_17[66]}
   );
   gpc606_5 gpc6258 (
      {stage1_17[88], stage1_17[89], stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[6],stage2_19[14],stage2_18[67],stage2_17[67]}
   );
   gpc606_5 gpc6259 (
      {stage1_17[94], stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[7],stage2_19[15],stage2_18[68],stage2_17[68]}
   );
   gpc606_5 gpc6260 (
      {stage1_17[100], stage1_17[101], stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[8],stage2_19[16],stage2_18[69],stage2_17[69]}
   );
   gpc606_5 gpc6261 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[9],stage2_19[17],stage2_18[70],stage2_17[70]}
   );
   gpc606_5 gpc6262 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[10],stage2_19[18],stage2_18[71],stage2_17[71]}
   );
   gpc606_5 gpc6263 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[11],stage2_19[19],stage2_18[72],stage2_17[72]}
   );
   gpc606_5 gpc6264 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[12],stage2_19[20],stage2_18[73],stage2_17[73]}
   );
   gpc606_5 gpc6265 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[13],stage2_19[21],stage2_18[74],stage2_17[74]}
   );
   gpc606_5 gpc6266 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[14],stage2_19[22],stage2_18[75],stage2_17[75]}
   );
   gpc606_5 gpc6267 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[15],stage2_19[23],stage2_18[76],stage2_17[76]}
   );
   gpc606_5 gpc6268 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[16],stage2_19[24],stage2_18[77],stage2_17[77]}
   );
   gpc606_5 gpc6269 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[17],stage2_19[25],stage2_18[78],stage2_17[78]}
   );
   gpc606_5 gpc6270 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[18],stage2_19[26],stage2_18[79],stage2_17[79]}
   );
   gpc606_5 gpc6271 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[19],stage2_19[27],stage2_18[80],stage2_17[80]}
   );
   gpc606_5 gpc6272 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[20],stage2_19[28],stage2_18[81],stage2_17[81]}
   );
   gpc606_5 gpc6273 (
      {stage1_17[178], stage1_17[179], stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[21],stage2_19[29],stage2_18[82],stage2_17[82]}
   );
   gpc606_5 gpc6274 (
      {stage1_17[184], stage1_17[185], stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[22],stage2_19[30],stage2_18[83],stage2_17[83]}
   );
   gpc606_5 gpc6275 (
      {stage1_17[190], stage1_17[191], stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[23],stage2_19[31],stage2_18[84],stage2_17[84]}
   );
   gpc606_5 gpc6276 (
      {stage1_17[196], stage1_17[197], stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[24],stage2_19[32],stage2_18[85],stage2_17[85]}
   );
   gpc606_5 gpc6277 (
      {stage1_17[202], stage1_17[203], stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[25],stage2_19[33],stage2_18[86],stage2_17[86]}
   );
   gpc606_5 gpc6278 (
      {stage1_17[208], stage1_17[209], stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[26],stage2_19[34],stage2_18[87],stage2_17[87]}
   );
   gpc606_5 gpc6279 (
      {stage1_17[214], stage1_17[215], stage1_17[216], stage1_17[217], 1'b0, 1'b0},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[27],stage2_19[35],stage2_18[88],stage2_17[88]}
   );
   gpc606_5 gpc6280 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[28],stage2_19[36],stage2_18[89],stage2_17[89]}
   );
   gpc606_5 gpc6281 (
      {stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[25],stage2_20[29],stage2_19[37],stage2_18[90]}
   );
   gpc606_5 gpc6282 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36], stage1_18[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[26],stage2_20[30],stage2_19[38],stage2_18[91]}
   );
   gpc606_5 gpc6283 (
      {stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42], stage1_18[43]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[27],stage2_20[31],stage2_19[39],stage2_18[92]}
   );
   gpc606_5 gpc6284 (
      {stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48], stage1_18[49]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[28],stage2_20[32],stage2_19[40],stage2_18[93]}
   );
   gpc606_5 gpc6285 (
      {stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54], stage1_18[55]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[29],stage2_20[33],stage2_19[41],stage2_18[94]}
   );
   gpc606_5 gpc6286 (
      {stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[30],stage2_20[34],stage2_19[42],stage2_18[95]}
   );
   gpc606_5 gpc6287 (
      {stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[31],stage2_20[35],stage2_19[43],stage2_18[96]}
   );
   gpc606_5 gpc6288 (
      {stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[32],stage2_20[36],stage2_19[44],stage2_18[97]}
   );
   gpc615_5 gpc6289 (
      {stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77], stage1_18[78]},
      {stage1_19[150]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[33],stage2_20[37],stage2_19[45],stage2_18[98]}
   );
   gpc615_5 gpc6290 (
      {stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_19[151]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[34],stage2_20[38],stage2_19[46],stage2_18[99]}
   );
   gpc615_5 gpc6291 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[152]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[35],stage2_20[39],stage2_19[47],stage2_18[100]}
   );
   gpc615_5 gpc6292 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[153]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[36],stage2_20[40],stage2_19[48],stage2_18[101]}
   );
   gpc615_5 gpc6293 (
      {stage1_18[94], stage1_18[95], stage1_18[96], stage1_18[97], stage1_18[98]},
      {stage1_19[154]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[37],stage2_20[41],stage2_19[49],stage2_18[102]}
   );
   gpc615_5 gpc6294 (
      {stage1_18[99], stage1_18[100], stage1_18[101], stage1_18[102], stage1_18[103]},
      {stage1_19[155]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[38],stage2_20[42],stage2_19[50],stage2_18[103]}
   );
   gpc615_5 gpc6295 (
      {stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107], stage1_18[108]},
      {stage1_19[156]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[39],stage2_20[43],stage2_19[51],stage2_18[104]}
   );
   gpc615_5 gpc6296 (
      {stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_19[157]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[40],stage2_20[44],stage2_19[52],stage2_18[105]}
   );
   gpc615_5 gpc6297 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118]},
      {stage1_19[158]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[41],stage2_20[45],stage2_19[53],stage2_18[106]}
   );
   gpc615_5 gpc6298 (
      {stage1_18[119], stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123]},
      {stage1_19[159]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[42],stage2_20[46],stage2_19[54],stage2_18[107]}
   );
   gpc615_5 gpc6299 (
      {stage1_18[124], stage1_18[125], stage1_18[126], stage1_18[127], stage1_18[128]},
      {stage1_19[160]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[43],stage2_20[47],stage2_19[55],stage2_18[108]}
   );
   gpc615_5 gpc6300 (
      {stage1_18[129], stage1_18[130], stage1_18[131], stage1_18[132], stage1_18[133]},
      {stage1_19[161]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[44],stage2_20[48],stage2_19[56],stage2_18[109]}
   );
   gpc615_5 gpc6301 (
      {stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137], stage1_18[138]},
      {stage1_19[162]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[45],stage2_20[49],stage2_19[57],stage2_18[110]}
   );
   gpc615_5 gpc6302 (
      {stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_19[163]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[46],stage2_20[50],stage2_19[58],stage2_18[111]}
   );
   gpc615_5 gpc6303 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148]},
      {stage1_19[164]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[47],stage2_20[51],stage2_19[59],stage2_18[112]}
   );
   gpc615_5 gpc6304 (
      {stage1_18[149], stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153]},
      {stage1_19[165]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[48],stage2_20[52],stage2_19[60],stage2_18[113]}
   );
   gpc615_5 gpc6305 (
      {stage1_18[154], stage1_18[155], stage1_18[156], stage1_18[157], stage1_18[158]},
      {stage1_19[166]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[49],stage2_20[53],stage2_19[61],stage2_18[114]}
   );
   gpc615_5 gpc6306 (
      {stage1_18[159], stage1_18[160], stage1_18[161], stage1_18[162], stage1_18[163]},
      {stage1_19[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[50],stage2_20[54],stage2_19[62],stage2_18[115]}
   );
   gpc615_5 gpc6307 (
      {stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167], stage1_18[168]},
      {stage1_19[168]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[51],stage2_20[55],stage2_19[63],stage2_18[116]}
   );
   gpc615_5 gpc6308 (
      {stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_19[169]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[52],stage2_20[56],stage2_19[64],stage2_18[117]}
   );
   gpc615_5 gpc6309 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[170]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[53],stage2_20[57],stage2_19[65],stage2_18[118]}
   );
   gpc615_5 gpc6310 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[171]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[54],stage2_20[58],stage2_19[66],stage2_18[119]}
   );
   gpc615_5 gpc6311 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[172]},
      {stage1_20[180], stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185]},
      {stage2_22[30],stage2_21[55],stage2_20[59],stage2_19[67],stage2_18[120]}
   );
   gpc615_5 gpc6312 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[173]},
      {stage1_20[186], stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage2_22[31],stage2_21[56],stage2_20[60],stage2_19[68],stage2_18[121]}
   );
   gpc615_5 gpc6313 (
      {stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197], stage1_18[198]},
      {stage1_19[174]},
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197]},
      {stage2_22[32],stage2_21[57],stage2_20[61],stage2_19[69],stage2_18[122]}
   );
   gpc615_5 gpc6314 (
      {stage1_18[199], stage1_18[200], stage1_18[201], stage1_18[202], stage1_18[203]},
      {stage1_19[175]},
      {stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203]},
      {stage2_22[33],stage2_21[58],stage2_20[62],stage2_19[70],stage2_18[123]}
   );
   gpc615_5 gpc6315 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[204]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[34],stage2_21[59],stage2_20[63],stage2_19[71]}
   );
   gpc615_5 gpc6316 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[205]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[35],stage2_21[60],stage2_20[64],stage2_19[72]}
   );
   gpc615_5 gpc6317 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[206]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[36],stage2_21[61],stage2_20[65],stage2_19[73]}
   );
   gpc615_5 gpc6318 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[207]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[37],stage2_21[62],stage2_20[66],stage2_19[74]}
   );
   gpc615_5 gpc6319 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[208]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[38],stage2_21[63],stage2_20[67],stage2_19[75]}
   );
   gpc606_5 gpc6320 (
      {stage1_20[209], stage1_20[210], stage1_20[211], stage1_20[212], stage1_20[213], stage1_20[214]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[39],stage2_21[64],stage2_20[68]}
   );
   gpc606_5 gpc6321 (
      {stage1_20[215], stage1_20[216], stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[40],stage2_21[65],stage2_20[69]}
   );
   gpc606_5 gpc6322 (
      {stage1_20[221], stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[41],stage2_21[66],stage2_20[70]}
   );
   gpc606_5 gpc6323 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[3],stage2_23[8],stage2_22[42],stage2_21[67]}
   );
   gpc606_5 gpc6324 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[4],stage2_23[9],stage2_22[43],stage2_21[68]}
   );
   gpc606_5 gpc6325 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[5],stage2_23[10],stage2_22[44],stage2_21[69]}
   );
   gpc606_5 gpc6326 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[6],stage2_23[11],stage2_22[45],stage2_21[70]}
   );
   gpc606_5 gpc6327 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[7],stage2_23[12],stage2_22[46],stage2_21[71]}
   );
   gpc606_5 gpc6328 (
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[8],stage2_23[13],stage2_22[47],stage2_21[72]}
   );
   gpc606_5 gpc6329 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[9],stage2_23[14],stage2_22[48],stage2_21[73]}
   );
   gpc606_5 gpc6330 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[10],stage2_23[15],stage2_22[49],stage2_21[74]}
   );
   gpc606_5 gpc6331 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[11],stage2_23[16],stage2_22[50],stage2_21[75]}
   );
   gpc606_5 gpc6332 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[12],stage2_23[17],stage2_22[51],stage2_21[76]}
   );
   gpc606_5 gpc6333 (
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[13],stage2_23[18],stage2_22[52],stage2_21[77]}
   );
   gpc606_5 gpc6334 (
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[14],stage2_23[19],stage2_22[53],stage2_21[78]}
   );
   gpc606_5 gpc6335 (
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[15],stage2_23[20],stage2_22[54],stage2_21[79]}
   );
   gpc606_5 gpc6336 (
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[16],stage2_23[21],stage2_22[55],stage2_21[80]}
   );
   gpc606_5 gpc6337 (
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[17],stage2_23[22],stage2_22[56],stage2_21[81]}
   );
   gpc606_5 gpc6338 (
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[18],stage2_23[23],stage2_22[57],stage2_21[82]}
   );
   gpc606_5 gpc6339 (
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[19],stage2_23[24],stage2_22[58],stage2_21[83]}
   );
   gpc606_5 gpc6340 (
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[20],stage2_23[25],stage2_22[59],stage2_21[84]}
   );
   gpc606_5 gpc6341 (
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[21],stage2_23[26],stage2_22[60],stage2_21[85]}
   );
   gpc606_5 gpc6342 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[22],stage2_23[27],stage2_22[61],stage2_21[86]}
   );
   gpc606_5 gpc6343 (
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[23],stage2_23[28],stage2_22[62],stage2_21[87]}
   );
   gpc606_5 gpc6344 (
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[24],stage2_23[29],stage2_22[63],stage2_21[88]}
   );
   gpc606_5 gpc6345 (
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[25],stage2_23[30],stage2_22[64],stage2_21[89]}
   );
   gpc606_5 gpc6346 (
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[26],stage2_23[31],stage2_22[65],stage2_21[90]}
   );
   gpc606_5 gpc6347 (
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[27],stage2_23[32],stage2_22[66],stage2_21[91]}
   );
   gpc606_5 gpc6348 (
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[28],stage2_23[33],stage2_22[67],stage2_21[92]}
   );
   gpc606_5 gpc6349 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[26],stage2_24[29],stage2_23[34],stage2_22[68]}
   );
   gpc615_5 gpc6350 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[156]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[27],stage2_24[30],stage2_23[35],stage2_22[69]}
   );
   gpc615_5 gpc6351 (
      {stage1_22[29], stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33]},
      {stage1_23[157]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[28],stage2_24[31],stage2_23[36],stage2_22[70]}
   );
   gpc615_5 gpc6352 (
      {stage1_22[34], stage1_22[35], stage1_22[36], stage1_22[37], stage1_22[38]},
      {stage1_23[158]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[29],stage2_24[32],stage2_23[37],stage2_22[71]}
   );
   gpc615_5 gpc6353 (
      {stage1_22[39], stage1_22[40], stage1_22[41], stage1_22[42], stage1_22[43]},
      {stage1_23[159]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[30],stage2_24[33],stage2_23[38],stage2_22[72]}
   );
   gpc615_5 gpc6354 (
      {stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47], stage1_22[48]},
      {stage1_23[160]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[31],stage2_24[34],stage2_23[39],stage2_22[73]}
   );
   gpc615_5 gpc6355 (
      {stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_23[161]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[32],stage2_24[35],stage2_23[40],stage2_22[74]}
   );
   gpc615_5 gpc6356 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58]},
      {stage1_23[162]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[33],stage2_24[36],stage2_23[41],stage2_22[75]}
   );
   gpc615_5 gpc6357 (
      {stage1_22[59], stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63]},
      {stage1_23[163]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[34],stage2_24[37],stage2_23[42],stage2_22[76]}
   );
   gpc615_5 gpc6358 (
      {stage1_22[64], stage1_22[65], stage1_22[66], stage1_22[67], stage1_22[68]},
      {stage1_23[164]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[35],stage2_24[38],stage2_23[43],stage2_22[77]}
   );
   gpc615_5 gpc6359 (
      {stage1_22[69], stage1_22[70], stage1_22[71], stage1_22[72], stage1_22[73]},
      {stage1_23[165]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[36],stage2_24[39],stage2_23[44],stage2_22[78]}
   );
   gpc615_5 gpc6360 (
      {stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77], stage1_22[78]},
      {stage1_23[166]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[37],stage2_24[40],stage2_23[45],stage2_22[79]}
   );
   gpc615_5 gpc6361 (
      {stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage1_23[167]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[38],stage2_24[41],stage2_23[46],stage2_22[80]}
   );
   gpc615_5 gpc6362 (
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88]},
      {stage1_23[168]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[39],stage2_24[42],stage2_23[47],stage2_22[81]}
   );
   gpc615_5 gpc6363 (
      {stage1_22[89], stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93]},
      {stage1_23[169]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[40],stage2_24[43],stage2_23[48],stage2_22[82]}
   );
   gpc615_5 gpc6364 (
      {stage1_22[94], stage1_22[95], stage1_22[96], stage1_22[97], stage1_22[98]},
      {stage1_23[170]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[41],stage2_24[44],stage2_23[49],stage2_22[83]}
   );
   gpc615_5 gpc6365 (
      {stage1_22[99], stage1_22[100], stage1_22[101], stage1_22[102], stage1_22[103]},
      {stage1_23[171]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[42],stage2_24[45],stage2_23[50],stage2_22[84]}
   );
   gpc615_5 gpc6366 (
      {stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108]},
      {stage1_23[172]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[43],stage2_24[46],stage2_23[51],stage2_22[85]}
   );
   gpc615_5 gpc6367 (
      {stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage1_23[173]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[44],stage2_24[47],stage2_23[52],stage2_22[86]}
   );
   gpc615_5 gpc6368 (
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118]},
      {stage1_23[174]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[45],stage2_24[48],stage2_23[53],stage2_22[87]}
   );
   gpc615_5 gpc6369 (
      {stage1_22[119], stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123]},
      {stage1_23[175]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[46],stage2_24[49],stage2_23[54],stage2_22[88]}
   );
   gpc615_5 gpc6370 (
      {stage1_22[124], stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128]},
      {stage1_23[176]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[47],stage2_24[50],stage2_23[55],stage2_22[89]}
   );
   gpc615_5 gpc6371 (
      {stage1_22[129], stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133]},
      {stage1_23[177]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[48],stage2_24[51],stage2_23[56],stage2_22[90]}
   );
   gpc615_5 gpc6372 (
      {stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138]},
      {stage1_23[178]},
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage2_26[23],stage2_25[49],stage2_24[52],stage2_23[57],stage2_22[91]}
   );
   gpc615_5 gpc6373 (
      {stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage1_23[179]},
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage2_26[24],stage2_25[50],stage2_24[53],stage2_23[58],stage2_22[92]}
   );
   gpc615_5 gpc6374 (
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148]},
      {stage1_23[180]},
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage2_26[25],stage2_25[51],stage2_24[54],stage2_23[59],stage2_22[93]}
   );
   gpc615_5 gpc6375 (
      {stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153]},
      {stage1_23[181]},
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage2_26[26],stage2_25[52],stage2_24[55],stage2_23[60],stage2_22[94]}
   );
   gpc615_5 gpc6376 (
      {stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157], stage1_22[158]},
      {stage1_23[182]},
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage2_26[27],stage2_25[53],stage2_24[56],stage2_23[61],stage2_22[95]}
   );
   gpc615_5 gpc6377 (
      {stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162], stage1_22[163]},
      {stage1_23[183]},
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage2_26[28],stage2_25[54],stage2_24[57],stage2_23[62],stage2_22[96]}
   );
   gpc615_5 gpc6378 (
      {stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167], stage1_22[168]},
      {stage1_23[184]},
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage2_26[29],stage2_25[55],stage2_24[58],stage2_23[63],stage2_22[97]}
   );
   gpc615_5 gpc6379 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173]},
      {stage1_23[185]},
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage2_26[30],stage2_25[56],stage2_24[59],stage2_23[64],stage2_22[98]}
   );
   gpc615_5 gpc6380 (
      {stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178]},
      {stage1_23[186]},
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage2_26[31],stage2_25[57],stage2_24[60],stage2_23[65],stage2_22[99]}
   );
   gpc615_5 gpc6381 (
      {stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182], stage1_22[183]},
      {stage1_23[187]},
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage2_26[32],stage2_25[58],stage2_24[61],stage2_23[66],stage2_22[100]}
   );
   gpc615_5 gpc6382 (
      {stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187], stage1_22[188]},
      {stage1_23[188]},
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage2_26[33],stage2_25[59],stage2_24[62],stage2_23[67],stage2_22[101]}
   );
   gpc615_5 gpc6383 (
      {stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192], stage1_22[193]},
      {stage1_23[189]},
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage2_26[34],stage2_25[60],stage2_24[63],stage2_23[68],stage2_22[102]}
   );
   gpc615_5 gpc6384 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[210]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[35],stage2_25[61],stage2_24[64],stage2_23[69]}
   );
   gpc615_5 gpc6385 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[211]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[36],stage2_25[62],stage2_24[65],stage2_23[70]}
   );
   gpc615_5 gpc6386 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[212]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[37],stage2_25[63],stage2_24[66],stage2_23[71]}
   );
   gpc615_5 gpc6387 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[213]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[38],stage2_25[64],stage2_24[67],stage2_23[72]}
   );
   gpc615_5 gpc6388 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[214]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[39],stage2_25[65],stage2_24[68],stage2_23[73]}
   );
   gpc615_5 gpc6389 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[215]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[40],stage2_25[66],stage2_24[69],stage2_23[74]}
   );
   gpc615_5 gpc6390 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[216]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[41],stage2_25[67],stage2_24[70],stage2_23[75]}
   );
   gpc615_5 gpc6391 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[217]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[42],stage2_25[68],stage2_24[71],stage2_23[76]}
   );
   gpc615_5 gpc6392 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[218]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[43],stage2_25[69],stage2_24[72],stage2_23[77]}
   );
   gpc615_5 gpc6393 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[219]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[44],stage2_25[70],stage2_24[73],stage2_23[78]}
   );
   gpc615_5 gpc6394 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[220]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[45],stage2_25[71],stage2_24[74],stage2_23[79]}
   );
   gpc615_5 gpc6395 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[221]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[46],stage2_25[72],stage2_24[75],stage2_23[80]}
   );
   gpc615_5 gpc6396 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[222]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[47],stage2_25[73],stage2_24[76],stage2_23[81]}
   );
   gpc615_5 gpc6397 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[223]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[48],stage2_25[74],stage2_24[77],stage2_23[82]}
   );
   gpc615_5 gpc6398 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[224]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[49],stage2_25[75],stage2_24[78],stage2_23[83]}
   );
   gpc615_5 gpc6399 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[225]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[50],stage2_25[76],stage2_24[79],stage2_23[84]}
   );
   gpc615_5 gpc6400 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[226]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[51],stage2_25[77],stage2_24[80],stage2_23[85]}
   );
   gpc615_5 gpc6401 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[227]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[52],stage2_25[78],stage2_24[81],stage2_23[86]}
   );
   gpc615_5 gpc6402 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[228]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[53],stage2_25[79],stage2_24[82],stage2_23[87]}
   );
   gpc615_5 gpc6403 (
      {stage1_23[285], stage1_23[286], stage1_23[287], stage1_23[288], stage1_23[289]},
      {stage1_24[229]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[54],stage2_25[80],stage2_24[83],stage2_23[88]}
   );
   gpc606_5 gpc6404 (
      {stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233], stage1_24[234], 1'b0},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[20],stage2_26[55],stage2_25[81],stage2_24[84]}
   );
   gpc606_5 gpc6405 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[1],stage2_27[21],stage2_26[56],stage2_25[82]}
   );
   gpc606_5 gpc6406 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[2],stage2_27[22],stage2_26[57],stage2_25[83]}
   );
   gpc606_5 gpc6407 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[3],stage2_27[23],stage2_26[58],stage2_25[84]}
   );
   gpc606_5 gpc6408 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[4],stage2_27[24],stage2_26[59],stage2_25[85]}
   );
   gpc606_5 gpc6409 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[5],stage2_27[25],stage2_26[60],stage2_25[86]}
   );
   gpc606_5 gpc6410 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[6],stage2_27[26],stage2_26[61],stage2_25[87]}
   );
   gpc606_5 gpc6411 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[7],stage2_27[27],stage2_26[62],stage2_25[88]}
   );
   gpc606_5 gpc6412 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[8],stage2_27[28],stage2_26[63],stage2_25[89]}
   );
   gpc606_5 gpc6413 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[9],stage2_27[29],stage2_26[64],stage2_25[90]}
   );
   gpc606_5 gpc6414 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[10],stage2_27[30],stage2_26[65],stage2_25[91]}
   );
   gpc615_5 gpc6415 (
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10]},
      {stage1_27[60]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[10],stage2_28[11],stage2_27[31],stage2_26[66]}
   );
   gpc615_5 gpc6416 (
      {stage1_26[11], stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15]},
      {stage1_27[61]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[11],stage2_28[12],stage2_27[32],stage2_26[67]}
   );
   gpc615_5 gpc6417 (
      {stage1_26[16], stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20]},
      {stage1_27[62]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[12],stage2_28[13],stage2_27[33],stage2_26[68]}
   );
   gpc615_5 gpc6418 (
      {stage1_26[21], stage1_26[22], stage1_26[23], stage1_26[24], stage1_26[25]},
      {stage1_27[63]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[13],stage2_28[14],stage2_27[34],stage2_26[69]}
   );
   gpc615_5 gpc6419 (
      {stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29], stage1_26[30]},
      {stage1_27[64]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[14],stage2_28[15],stage2_27[35],stage2_26[70]}
   );
   gpc615_5 gpc6420 (
      {stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[65]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[15],stage2_28[16],stage2_27[36],stage2_26[71]}
   );
   gpc615_5 gpc6421 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40]},
      {stage1_27[66]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[16],stage2_28[17],stage2_27[37],stage2_26[72]}
   );
   gpc615_5 gpc6422 (
      {stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45]},
      {stage1_27[67]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[17],stage2_28[18],stage2_27[38],stage2_26[73]}
   );
   gpc615_5 gpc6423 (
      {stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49], stage1_26[50]},
      {stage1_27[68]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[18],stage2_28[19],stage2_27[39],stage2_26[74]}
   );
   gpc615_5 gpc6424 (
      {stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54], stage1_26[55]},
      {stage1_27[69]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[19],stage2_28[20],stage2_27[40],stage2_26[75]}
   );
   gpc615_5 gpc6425 (
      {stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59], stage1_26[60]},
      {stage1_27[70]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[20],stage2_28[21],stage2_27[41],stage2_26[76]}
   );
   gpc615_5 gpc6426 (
      {stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage1_27[71]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[21],stage2_28[22],stage2_27[42],stage2_26[77]}
   );
   gpc615_5 gpc6427 (
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70]},
      {stage1_27[72]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[22],stage2_28[23],stage2_27[43],stage2_26[78]}
   );
   gpc615_5 gpc6428 (
      {stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75]},
      {stage1_27[73]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[23],stage2_28[24],stage2_27[44],stage2_26[79]}
   );
   gpc615_5 gpc6429 (
      {stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79], stage1_26[80]},
      {stage1_27[74]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[24],stage2_28[25],stage2_27[45],stage2_26[80]}
   );
   gpc615_5 gpc6430 (
      {stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84], stage1_26[85]},
      {stage1_27[75]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[25],stage2_28[26],stage2_27[46],stage2_26[81]}
   );
   gpc615_5 gpc6431 (
      {stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89], stage1_26[90]},
      {stage1_27[76]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[26],stage2_28[27],stage2_27[47],stage2_26[82]}
   );
   gpc615_5 gpc6432 (
      {stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage1_27[77]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[27],stage2_28[28],stage2_27[48],stage2_26[83]}
   );
   gpc615_5 gpc6433 (
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100]},
      {stage1_27[78]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[28],stage2_28[29],stage2_27[49],stage2_26[84]}
   );
   gpc615_5 gpc6434 (
      {stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105]},
      {stage1_27[79]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[29],stage2_28[30],stage2_27[50],stage2_26[85]}
   );
   gpc615_5 gpc6435 (
      {stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109], stage1_26[110]},
      {stage1_27[80]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[30],stage2_28[31],stage2_27[51],stage2_26[86]}
   );
   gpc615_5 gpc6436 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[81]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[31],stage2_28[32],stage2_27[52],stage2_26[87]}
   );
   gpc615_5 gpc6437 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[82]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[32],stage2_28[33],stage2_27[53],stage2_26[88]}
   );
   gpc615_5 gpc6438 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[83]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[33],stage2_28[34],stage2_27[54],stage2_26[89]}
   );
   gpc615_5 gpc6439 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[84]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[34],stage2_28[35],stage2_27[55],stage2_26[90]}
   );
   gpc615_5 gpc6440 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[85]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[35],stage2_28[36],stage2_27[56],stage2_26[91]}
   );
   gpc615_5 gpc6441 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[86]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[36],stage2_28[37],stage2_27[57],stage2_26[92]}
   );
   gpc615_5 gpc6442 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[87]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[37],stage2_28[38],stage2_27[58],stage2_26[93]}
   );
   gpc615_5 gpc6443 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[88]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[38],stage2_28[39],stage2_27[59],stage2_26[94]}
   );
   gpc623_5 gpc6444 (
      {stage1_26[151], stage1_26[152], stage1_26[153]},
      {stage1_27[89], stage1_27[90]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[39],stage2_28[40],stage2_27[60],stage2_26[95]}
   );
   gpc615_5 gpc6445 (
      {stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage1_28[180]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[30],stage2_29[40],stage2_28[41],stage2_27[61]}
   );
   gpc615_5 gpc6446 (
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100]},
      {stage1_28[181]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[31],stage2_29[41],stage2_28[42],stage2_27[62]}
   );
   gpc615_5 gpc6447 (
      {stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105]},
      {stage1_28[182]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[32],stage2_29[42],stage2_28[43],stage2_27[63]}
   );
   gpc615_5 gpc6448 (
      {stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109], stage1_27[110]},
      {stage1_28[183]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[33],stage2_29[43],stage2_28[44],stage2_27[64]}
   );
   gpc615_5 gpc6449 (
      {stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114], stage1_27[115]},
      {stage1_28[184]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[34],stage2_29[44],stage2_28[45],stage2_27[65]}
   );
   gpc615_5 gpc6450 (
      {stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119], stage1_27[120]},
      {stage1_28[185]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[35],stage2_29[45],stage2_28[46],stage2_27[66]}
   );
   gpc615_5 gpc6451 (
      {stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage1_28[186]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[36],stage2_29[46],stage2_28[47],stage2_27[67]}
   );
   gpc615_5 gpc6452 (
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130]},
      {stage1_28[187]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[37],stage2_29[47],stage2_28[48],stage2_27[68]}
   );
   gpc615_5 gpc6453 (
      {stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135]},
      {stage1_28[188]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[38],stage2_29[48],stage2_28[49],stage2_27[69]}
   );
   gpc615_5 gpc6454 (
      {stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139], stage1_27[140]},
      {stage1_28[189]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[39],stage2_29[49],stage2_28[50],stage2_27[70]}
   );
   gpc615_5 gpc6455 (
      {stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144], stage1_27[145]},
      {stage1_28[190]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[40],stage2_29[50],stage2_28[51],stage2_27[71]}
   );
   gpc615_5 gpc6456 (
      {stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149], stage1_27[150]},
      {stage1_28[191]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[41],stage2_29[51],stage2_28[52],stage2_27[72]}
   );
   gpc615_5 gpc6457 (
      {stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage1_28[192]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[42],stage2_29[52],stage2_28[53],stage2_27[73]}
   );
   gpc615_5 gpc6458 (
      {stage1_27[156], stage1_27[157], stage1_27[158], stage1_27[159], stage1_27[160]},
      {stage1_28[193]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[43],stage2_29[53],stage2_28[54],stage2_27[74]}
   );
   gpc615_5 gpc6459 (
      {stage1_27[161], stage1_27[162], stage1_27[163], stage1_27[164], stage1_27[165]},
      {stage1_28[194]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[44],stage2_29[54],stage2_28[55],stage2_27[75]}
   );
   gpc615_5 gpc6460 (
      {stage1_27[166], stage1_27[167], stage1_27[168], stage1_27[169], stage1_27[170]},
      {stage1_28[195]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[45],stage2_29[55],stage2_28[56],stage2_27[76]}
   );
   gpc615_5 gpc6461 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[196]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[46],stage2_29[56],stage2_28[57],stage2_27[77]}
   );
   gpc615_5 gpc6462 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[197]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[47],stage2_29[57],stage2_28[58],stage2_27[78]}
   );
   gpc615_5 gpc6463 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[198]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[48],stage2_29[58],stage2_28[59],stage2_27[79]}
   );
   gpc615_5 gpc6464 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[199]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[49],stage2_29[59],stage2_28[60],stage2_27[80]}
   );
   gpc615_5 gpc6465 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[200]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[50],stage2_29[60],stage2_28[61],stage2_27[81]}
   );
   gpc615_5 gpc6466 (
      {stage1_27[196], stage1_27[197], stage1_27[198], stage1_27[199], stage1_27[200]},
      {stage1_28[201]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[51],stage2_29[61],stage2_28[62],stage2_27[82]}
   );
   gpc615_5 gpc6467 (
      {stage1_27[201], stage1_27[202], stage1_27[203], stage1_27[204], stage1_27[205]},
      {stage1_28[202]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[52],stage2_29[62],stage2_28[63],stage2_27[83]}
   );
   gpc615_5 gpc6468 (
      {stage1_27[206], stage1_27[207], stage1_27[208], stage1_27[209], stage1_27[210]},
      {stage1_28[203]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[53],stage2_29[63],stage2_28[64],stage2_27[84]}
   );
   gpc606_5 gpc6469 (
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[24],stage2_30[54],stage2_29[64],stage2_28[65]}
   );
   gpc606_5 gpc6470 (
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[25],stage2_30[55],stage2_29[65],stage2_28[66]}
   );
   gpc606_5 gpc6471 (
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[26],stage2_30[56],stage2_29[66],stage2_28[67]}
   );
   gpc606_5 gpc6472 (
      {stage1_28[222], stage1_28[223], stage1_28[224], stage1_28[225], stage1_28[226], stage1_28[227]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[27],stage2_30[57],stage2_29[67],stage2_28[68]}
   );
   gpc606_5 gpc6473 (
      {stage1_28[228], stage1_28[229], stage1_28[230], stage1_28[231], stage1_28[232], stage1_28[233]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[28],stage2_30[58],stage2_29[68],stage2_28[69]}
   );
   gpc606_5 gpc6474 (
      {stage1_28[234], stage1_28[235], stage1_28[236], stage1_28[237], stage1_28[238], stage1_28[239]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[29],stage2_30[59],stage2_29[69],stage2_28[70]}
   );
   gpc606_5 gpc6475 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[6],stage2_31[30],stage2_30[60],stage2_29[70]}
   );
   gpc606_5 gpc6476 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[7],stage2_31[31],stage2_30[61],stage2_29[71]}
   );
   gpc606_5 gpc6477 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[8],stage2_31[32],stage2_30[62],stage2_29[72]}
   );
   gpc606_5 gpc6478 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[9],stage2_31[33],stage2_30[63],stage2_29[73]}
   );
   gpc606_5 gpc6479 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[10],stage2_31[34],stage2_30[64],stage2_29[74]}
   );
   gpc606_5 gpc6480 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[11],stage2_31[35],stage2_30[65],stage2_29[75]}
   );
   gpc606_5 gpc6481 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[12],stage2_31[36],stage2_30[66],stage2_29[76]}
   );
   gpc2135_5 gpc6482 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40]},
      {stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_32[0]},
      {stage1_33[0], stage1_33[1]},
      {stage2_34[0],stage2_33[7],stage2_32[13],stage2_31[37],stage2_30[67]}
   );
   gpc207_4 gpc6483 (
      {stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[1], stage1_32[2]},
      {stage2_33[8],stage2_32[14],stage2_31[38],stage2_30[68]}
   );
   gpc207_4 gpc6484 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_32[3], stage1_32[4]},
      {stage2_33[9],stage2_32[15],stage2_31[39],stage2_30[69]}
   );
   gpc207_4 gpc6485 (
      {stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_32[5], stage1_32[6]},
      {stage2_33[10],stage2_32[16],stage2_31[40],stage2_30[70]}
   );
   gpc207_4 gpc6486 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66], stage1_30[67], stage1_30[68]},
      {stage1_32[7], stage1_32[8]},
      {stage2_33[11],stage2_32[17],stage2_31[41],stage2_30[71]}
   );
   gpc207_4 gpc6487 (
      {stage1_30[69], stage1_30[70], stage1_30[71], stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75]},
      {stage1_32[9], stage1_32[10]},
      {stage2_33[12],stage2_32[18],stage2_31[42],stage2_30[72]}
   );
   gpc606_5 gpc6488 (
      {stage1_30[76], stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16]},
      {stage2_34[1],stage2_33[13],stage2_32[19],stage2_31[43],stage2_30[73]}
   );
   gpc606_5 gpc6489 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87]},
      {stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22]},
      {stage2_34[2],stage2_33[14],stage2_32[20],stage2_31[44],stage2_30[74]}
   );
   gpc606_5 gpc6490 (
      {stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93]},
      {stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28]},
      {stage2_34[3],stage2_33[15],stage2_32[21],stage2_31[45],stage2_30[75]}
   );
   gpc606_5 gpc6491 (
      {stage1_30[94], stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34]},
      {stage2_34[4],stage2_33[16],stage2_32[22],stage2_31[46],stage2_30[76]}
   );
   gpc606_5 gpc6492 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105]},
      {stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40]},
      {stage2_34[5],stage2_33[17],stage2_32[23],stage2_31[47],stage2_30[77]}
   );
   gpc606_5 gpc6493 (
      {stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111]},
      {stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46]},
      {stage2_34[6],stage2_33[18],stage2_32[24],stage2_31[48],stage2_30[78]}
   );
   gpc606_5 gpc6494 (
      {stage1_30[112], stage1_30[113], stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117]},
      {stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52]},
      {stage2_34[7],stage2_33[19],stage2_32[25],stage2_31[49],stage2_30[79]}
   );
   gpc606_5 gpc6495 (
      {stage1_30[118], stage1_30[119], stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123]},
      {stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58]},
      {stage2_34[8],stage2_33[20],stage2_32[26],stage2_31[50],stage2_30[80]}
   );
   gpc606_5 gpc6496 (
      {stage1_30[124], stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64]},
      {stage2_34[9],stage2_33[21],stage2_32[27],stage2_31[51],stage2_30[81]}
   );
   gpc606_5 gpc6497 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135]},
      {stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70]},
      {stage2_34[10],stage2_33[22],stage2_32[28],stage2_31[52],stage2_30[82]}
   );
   gpc606_5 gpc6498 (
      {stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141]},
      {stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76]},
      {stage2_34[11],stage2_33[23],stage2_32[29],stage2_31[53],stage2_30[83]}
   );
   gpc606_5 gpc6499 (
      {stage1_30[142], stage1_30[143], stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147]},
      {stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82]},
      {stage2_34[12],stage2_33[24],stage2_32[30],stage2_31[54],stage2_30[84]}
   );
   gpc606_5 gpc6500 (
      {stage1_30[148], stage1_30[149], stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153]},
      {stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88]},
      {stage2_34[13],stage2_33[25],stage2_32[31],stage2_31[55],stage2_30[85]}
   );
   gpc606_5 gpc6501 (
      {stage1_30[154], stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94]},
      {stage2_34[14],stage2_33[26],stage2_32[32],stage2_31[56],stage2_30[86]}
   );
   gpc606_5 gpc6502 (
      {stage1_30[160], stage1_30[161], stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165]},
      {stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100]},
      {stage2_34[15],stage2_33[27],stage2_32[33],stage2_31[57],stage2_30[87]}
   );
   gpc606_5 gpc6503 (
      {stage1_30[166], stage1_30[167], stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171]},
      {stage1_32[101], stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106]},
      {stage2_34[16],stage2_33[28],stage2_32[34],stage2_31[58],stage2_30[88]}
   );
   gpc606_5 gpc6504 (
      {stage1_30[172], stage1_30[173], stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177]},
      {stage1_32[107], stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112]},
      {stage2_34[17],stage2_33[29],stage2_32[35],stage2_31[59],stage2_30[89]}
   );
   gpc606_5 gpc6505 (
      {stage1_30[178], stage1_30[179], stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183]},
      {stage1_32[113], stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118]},
      {stage2_34[18],stage2_33[30],stage2_32[36],stage2_31[60],stage2_30[90]}
   );
   gpc606_5 gpc6506 (
      {stage1_30[184], stage1_30[185], stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189]},
      {stage1_32[119], stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124]},
      {stage2_34[19],stage2_33[31],stage2_32[37],stage2_31[61],stage2_30[91]}
   );
   gpc606_5 gpc6507 (
      {stage1_30[190], stage1_30[191], stage1_30[192], stage1_30[193], stage1_30[194], stage1_30[195]},
      {stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130]},
      {stage2_34[20],stage2_33[32],stage2_32[38],stage2_31[62],stage2_30[92]}
   );
   gpc606_5 gpc6508 (
      {stage1_30[196], stage1_30[197], stage1_30[198], stage1_30[199], stage1_30[200], stage1_30[201]},
      {stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136]},
      {stage2_34[21],stage2_33[33],stage2_32[39],stage2_31[63],stage2_30[93]}
   );
   gpc606_5 gpc6509 (
      {stage1_30[202], stage1_30[203], stage1_30[204], stage1_30[205], stage1_30[206], stage1_30[207]},
      {stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140], stage1_32[141], stage1_32[142]},
      {stage2_34[22],stage2_33[34],stage2_32[40],stage2_31[64],stage2_30[94]}
   );
   gpc606_5 gpc6510 (
      {stage1_30[208], stage1_30[209], stage1_30[210], stage1_30[211], stage1_30[212], stage1_30[213]},
      {stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146], stage1_32[147], stage1_32[148]},
      {stage2_34[23],stage2_33[35],stage2_32[41],stage2_31[65],stage2_30[95]}
   );
   gpc606_5 gpc6511 (
      {stage1_30[214], stage1_30[215], stage1_30[216], stage1_30[217], stage1_30[218], stage1_30[219]},
      {stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152], stage1_32[153], stage1_32[154]},
      {stage2_34[24],stage2_33[36],stage2_32[42],stage2_31[66],stage2_30[96]}
   );
   gpc606_5 gpc6512 (
      {stage1_30[220], stage1_30[221], stage1_30[222], stage1_30[223], stage1_30[224], stage1_30[225]},
      {stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158], stage1_32[159], stage1_32[160]},
      {stage2_34[25],stage2_33[37],stage2_32[43],stage2_31[67],stage2_30[97]}
   );
   gpc606_5 gpc6513 (
      {stage1_30[226], stage1_30[227], stage1_30[228], stage1_30[229], stage1_30[230], stage1_30[231]},
      {stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164], stage1_32[165], stage1_32[166]},
      {stage2_34[26],stage2_33[38],stage2_32[44],stage2_31[68],stage2_30[98]}
   );
   gpc615_5 gpc6514 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49]},
      {stage1_32[167]},
      {stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6], stage1_33[7]},
      {stage2_35[0],stage2_34[27],stage2_33[39],stage2_32[45],stage2_31[69]}
   );
   gpc615_5 gpc6515 (
      {stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54]},
      {stage1_32[168]},
      {stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12], stage1_33[13]},
      {stage2_35[1],stage2_34[28],stage2_33[40],stage2_32[46],stage2_31[70]}
   );
   gpc615_5 gpc6516 (
      {stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage1_32[169]},
      {stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18], stage1_33[19]},
      {stage2_35[2],stage2_34[29],stage2_33[41],stage2_32[47],stage2_31[71]}
   );
   gpc615_5 gpc6517 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64]},
      {stage1_32[170]},
      {stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24], stage1_33[25]},
      {stage2_35[3],stage2_34[30],stage2_33[42],stage2_32[48],stage2_31[72]}
   );
   gpc615_5 gpc6518 (
      {stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69]},
      {stage1_32[171]},
      {stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30], stage1_33[31]},
      {stage2_35[4],stage2_34[31],stage2_33[43],stage2_32[49],stage2_31[73]}
   );
   gpc615_5 gpc6519 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[172]},
      {stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36], stage1_33[37]},
      {stage2_35[5],stage2_34[32],stage2_33[44],stage2_32[50],stage2_31[74]}
   );
   gpc615_5 gpc6520 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79]},
      {stage1_32[173]},
      {stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42], stage1_33[43]},
      {stage2_35[6],stage2_34[33],stage2_33[45],stage2_32[51],stage2_31[75]}
   );
   gpc615_5 gpc6521 (
      {stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84]},
      {stage1_32[174]},
      {stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48], stage1_33[49]},
      {stage2_35[7],stage2_34[34],stage2_33[46],stage2_32[52],stage2_31[76]}
   );
   gpc615_5 gpc6522 (
      {stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_32[175]},
      {stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54], stage1_33[55]},
      {stage2_35[8],stage2_34[35],stage2_33[47],stage2_32[53],stage2_31[77]}
   );
   gpc615_5 gpc6523 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94]},
      {stage1_32[176]},
      {stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60], stage1_33[61]},
      {stage2_35[9],stage2_34[36],stage2_33[48],stage2_32[54],stage2_31[78]}
   );
   gpc615_5 gpc6524 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99]},
      {stage1_32[177]},
      {stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66], stage1_33[67]},
      {stage2_35[10],stage2_34[37],stage2_33[49],stage2_32[55],stage2_31[79]}
   );
   gpc615_5 gpc6525 (
      {stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_32[178]},
      {stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72], stage1_33[73]},
      {stage2_35[11],stage2_34[38],stage2_33[50],stage2_32[56],stage2_31[80]}
   );
   gpc615_5 gpc6526 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[179]},
      {stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78], stage1_33[79]},
      {stage2_35[12],stage2_34[39],stage2_33[51],stage2_32[57],stage2_31[81]}
   );
   gpc615_5 gpc6527 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[180]},
      {stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84], stage1_33[85]},
      {stage2_35[13],stage2_34[40],stage2_33[52],stage2_32[58],stage2_31[82]}
   );
   gpc615_5 gpc6528 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[181]},
      {stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90], stage1_33[91]},
      {stage2_35[14],stage2_34[41],stage2_33[53],stage2_32[59],stage2_31[83]}
   );
   gpc615_5 gpc6529 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[182]},
      {stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96], stage1_33[97]},
      {stage2_35[15],stage2_34[42],stage2_33[54],stage2_32[60],stage2_31[84]}
   );
   gpc615_5 gpc6530 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[183]},
      {stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102], stage1_33[103]},
      {stage2_35[16],stage2_34[43],stage2_33[55],stage2_32[61],stage2_31[85]}
   );
   gpc615_5 gpc6531 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[184]},
      {stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108], stage1_33[109]},
      {stage2_35[17],stage2_34[44],stage2_33[56],stage2_32[62],stage2_31[86]}
   );
   gpc615_5 gpc6532 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[185]},
      {stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114], stage1_33[115]},
      {stage2_35[18],stage2_34[45],stage2_33[57],stage2_32[63],stage2_31[87]}
   );
   gpc615_5 gpc6533 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[186]},
      {stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120], stage1_33[121]},
      {stage2_35[19],stage2_34[46],stage2_33[58],stage2_32[64],stage2_31[88]}
   );
   gpc615_5 gpc6534 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[187]},
      {stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126], stage1_33[127]},
      {stage2_35[20],stage2_34[47],stage2_33[59],stage2_32[65],stage2_31[89]}
   );
   gpc615_5 gpc6535 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[188]},
      {stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132], stage1_33[133]},
      {stage2_35[21],stage2_34[48],stage2_33[60],stage2_32[66],stage2_31[90]}
   );
   gpc615_5 gpc6536 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[189]},
      {stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138], stage1_33[139]},
      {stage2_35[22],stage2_34[49],stage2_33[61],stage2_32[67],stage2_31[91]}
   );
   gpc615_5 gpc6537 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[190]},
      {stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144], stage1_33[145]},
      {stage2_35[23],stage2_34[50],stage2_33[62],stage2_32[68],stage2_31[92]}
   );
   gpc615_5 gpc6538 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[191]},
      {stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150], stage1_33[151]},
      {stage2_35[24],stage2_34[51],stage2_33[63],stage2_32[69],stage2_31[93]}
   );
   gpc615_5 gpc6539 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[192]},
      {stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156], stage1_33[157]},
      {stage2_35[25],stage2_34[52],stage2_33[64],stage2_32[70],stage2_31[94]}
   );
   gpc615_5 gpc6540 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[193]},
      {stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162], stage1_33[163]},
      {stage2_35[26],stage2_34[53],stage2_33[65],stage2_32[71],stage2_31[95]}
   );
   gpc606_5 gpc6541 (
      {stage1_32[194], stage1_32[195], stage1_32[196], stage1_32[197], stage1_32[198], stage1_32[199]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[27],stage2_34[54],stage2_33[66],stage2_32[72]}
   );
   gpc606_5 gpc6542 (
      {stage1_32[200], stage1_32[201], stage1_32[202], stage1_32[203], stage1_32[204], stage1_32[205]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[28],stage2_34[55],stage2_33[67],stage2_32[73]}
   );
   gpc606_5 gpc6543 (
      {stage1_32[206], stage1_32[207], stage1_32[208], stage1_32[209], stage1_32[210], stage1_32[211]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[29],stage2_34[56],stage2_33[68],stage2_32[74]}
   );
   gpc606_5 gpc6544 (
      {stage1_32[212], stage1_32[213], stage1_32[214], stage1_32[215], stage1_32[216], stage1_32[217]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[30],stage2_34[57],stage2_33[69],stage2_32[75]}
   );
   gpc606_5 gpc6545 (
      {stage1_32[218], stage1_32[219], stage1_32[220], stage1_32[221], stage1_32[222], stage1_32[223]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[31],stage2_34[58],stage2_33[70],stage2_32[76]}
   );
   gpc606_5 gpc6546 (
      {stage1_32[224], stage1_32[225], stage1_32[226], stage1_32[227], stage1_32[228], stage1_32[229]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[32],stage2_34[59],stage2_33[71],stage2_32[77]}
   );
   gpc606_5 gpc6547 (
      {stage1_32[230], stage1_32[231], stage1_32[232], stage1_32[233], stage1_32[234], stage1_32[235]},
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage2_36[6],stage2_35[33],stage2_34[60],stage2_33[72],stage2_32[78]}
   );
   gpc606_5 gpc6548 (
      {stage1_32[236], stage1_32[237], stage1_32[238], stage1_32[239], stage1_32[240], stage1_32[241]},
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage2_36[7],stage2_35[34],stage2_34[61],stage2_33[73],stage2_32[79]}
   );
   gpc606_5 gpc6549 (
      {stage1_32[242], stage1_32[243], stage1_32[244], stage1_32[245], stage1_32[246], stage1_32[247]},
      {stage1_34[48], stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53]},
      {stage2_36[8],stage2_35[35],stage2_34[62],stage2_33[74],stage2_32[80]}
   );
   gpc606_5 gpc6550 (
      {stage1_32[248], stage1_32[249], stage1_32[250], stage1_32[251], stage1_32[252], stage1_32[253]},
      {stage1_34[54], stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59]},
      {stage2_36[9],stage2_35[36],stage2_34[63],stage2_33[75],stage2_32[81]}
   );
   gpc606_5 gpc6551 (
      {stage1_32[254], stage1_32[255], stage1_32[256], stage1_32[257], stage1_32[258], stage1_32[259]},
      {stage1_34[60], stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage2_36[10],stage2_35[37],stage2_34[64],stage2_33[76],stage2_32[82]}
   );
   gpc606_5 gpc6552 (
      {stage1_32[260], stage1_32[261], stage1_32[262], stage1_32[263], stage1_32[264], stage1_32[265]},
      {stage1_34[66], stage1_34[67], stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71]},
      {stage2_36[11],stage2_35[38],stage2_34[65],stage2_33[77],stage2_32[83]}
   );
   gpc606_5 gpc6553 (
      {stage1_32[266], stage1_32[267], stage1_32[268], stage1_32[269], stage1_32[270], stage1_32[271]},
      {stage1_34[72], stage1_34[73], stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77]},
      {stage2_36[12],stage2_35[39],stage2_34[66],stage2_33[78],stage2_32[84]}
   );
   gpc606_5 gpc6554 (
      {stage1_32[272], stage1_32[273], stage1_32[274], stage1_32[275], stage1_32[276], stage1_32[277]},
      {stage1_34[78], stage1_34[79], stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83]},
      {stage2_36[13],stage2_35[40],stage2_34[67],stage2_33[79],stage2_32[85]}
   );
   gpc606_5 gpc6555 (
      {stage1_32[278], stage1_32[279], stage1_32[280], stage1_32[281], stage1_32[282], stage1_32[283]},
      {stage1_34[84], stage1_34[85], stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89]},
      {stage2_36[14],stage2_35[41],stage2_34[68],stage2_33[80],stage2_32[86]}
   );
   gpc606_5 gpc6556 (
      {stage1_32[284], stage1_32[285], stage1_32[286], stage1_32[287], stage1_32[288], stage1_32[289]},
      {stage1_34[90], stage1_34[91], stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95]},
      {stage2_36[15],stage2_35[42],stage2_34[69],stage2_33[81],stage2_32[87]}
   );
   gpc606_5 gpc6557 (
      {stage1_32[290], stage1_32[291], stage1_32[292], stage1_32[293], stage1_32[294], stage1_32[295]},
      {stage1_34[96], stage1_34[97], stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101]},
      {stage2_36[16],stage2_35[43],stage2_34[70],stage2_33[82],stage2_32[88]}
   );
   gpc606_5 gpc6558 (
      {stage1_32[296], stage1_32[297], stage1_32[298], stage1_32[299], stage1_32[300], stage1_32[301]},
      {stage1_34[102], stage1_34[103], stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107]},
      {stage2_36[17],stage2_35[44],stage2_34[71],stage2_33[83],stage2_32[89]}
   );
   gpc606_5 gpc6559 (
      {stage1_32[302], stage1_32[303], stage1_32[304], stage1_32[305], stage1_32[306], stage1_32[307]},
      {stage1_34[108], stage1_34[109], stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113]},
      {stage2_36[18],stage2_35[45],stage2_34[72],stage2_33[84],stage2_32[90]}
   );
   gpc606_5 gpc6560 (
      {stage1_32[308], stage1_32[309], stage1_32[310], stage1_32[311], stage1_32[312], stage1_32[313]},
      {stage1_34[114], stage1_34[115], stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119]},
      {stage2_36[19],stage2_35[46],stage2_34[73],stage2_33[85],stage2_32[91]}
   );
   gpc606_5 gpc6561 (
      {stage1_32[314], stage1_32[315], stage1_32[316], stage1_32[317], stage1_32[318], stage1_32[319]},
      {stage1_34[120], stage1_34[121], stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125]},
      {stage2_36[20],stage2_35[47],stage2_34[74],stage2_33[86],stage2_32[92]}
   );
   gpc606_5 gpc6562 (
      {stage1_32[320], stage1_32[321], stage1_32[322], stage1_32[323], stage1_32[324], stage1_32[325]},
      {stage1_34[126], stage1_34[127], stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131]},
      {stage2_36[21],stage2_35[48],stage2_34[75],stage2_33[87],stage2_32[93]}
   );
   gpc606_5 gpc6563 (
      {stage1_32[326], stage1_32[327], stage1_32[328], stage1_32[329], stage1_32[330], stage1_32[331]},
      {stage1_34[132], stage1_34[133], stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137]},
      {stage2_36[22],stage2_35[49],stage2_34[76],stage2_33[88],stage2_32[94]}
   );
   gpc606_5 gpc6564 (
      {stage1_32[332], stage1_32[333], stage1_32[334], stage1_32[335], stage1_32[336], stage1_32[337]},
      {stage1_34[138], stage1_34[139], stage1_34[140], stage1_34[141], stage1_34[142], stage1_34[143]},
      {stage2_36[23],stage2_35[50],stage2_34[77],stage2_33[89],stage2_32[95]}
   );
   gpc606_5 gpc6565 (
      {stage1_32[338], stage1_32[339], stage1_32[340], stage1_32[341], stage1_32[342], stage1_32[343]},
      {stage1_34[144], stage1_34[145], stage1_34[146], stage1_34[147], stage1_34[148], stage1_34[149]},
      {stage2_36[24],stage2_35[51],stage2_34[78],stage2_33[90],stage2_32[96]}
   );
   gpc606_5 gpc6566 (
      {stage1_32[344], stage1_32[345], stage1_32[346], stage1_32[347], stage1_32[348], stage1_32[349]},
      {stage1_34[150], stage1_34[151], stage1_34[152], stage1_34[153], stage1_34[154], stage1_34[155]},
      {stage2_36[25],stage2_35[52],stage2_34[79],stage2_33[91],stage2_32[97]}
   );
   gpc606_5 gpc6567 (
      {stage1_32[350], stage1_32[351], stage1_32[352], stage1_32[353], stage1_32[354], stage1_32[355]},
      {stage1_34[156], stage1_34[157], stage1_34[158], stage1_34[159], stage1_34[160], stage1_34[161]},
      {stage2_36[26],stage2_35[53],stage2_34[80],stage2_33[92],stage2_32[98]}
   );
   gpc606_5 gpc6568 (
      {stage1_32[356], stage1_32[357], stage1_32[358], stage1_32[359], stage1_32[360], stage1_32[361]},
      {stage1_34[162], stage1_34[163], stage1_34[164], stage1_34[165], stage1_34[166], stage1_34[167]},
      {stage2_36[27],stage2_35[54],stage2_34[81],stage2_33[93],stage2_32[99]}
   );
   gpc606_5 gpc6569 (
      {stage1_32[362], stage1_32[363], stage1_32[364], stage1_32[365], stage1_32[366], stage1_32[367]},
      {stage1_34[168], stage1_34[169], stage1_34[170], stage1_34[171], stage1_34[172], stage1_34[173]},
      {stage2_36[28],stage2_35[55],stage2_34[82],stage2_33[94],stage2_32[100]}
   );
   gpc606_5 gpc6570 (
      {stage1_32[368], stage1_32[369], stage1_32[370], stage1_32[371], stage1_32[372], stage1_32[373]},
      {stage1_34[174], stage1_34[175], stage1_34[176], stage1_34[177], stage1_34[178], stage1_34[179]},
      {stage2_36[29],stage2_35[56],stage2_34[83],stage2_33[95],stage2_32[101]}
   );
   gpc606_5 gpc6571 (
      {stage1_32[374], stage1_32[375], stage1_32[376], stage1_32[377], stage1_32[378], stage1_32[379]},
      {stage1_34[180], stage1_34[181], stage1_34[182], stage1_34[183], stage1_34[184], stage1_34[185]},
      {stage2_36[30],stage2_35[57],stage2_34[84],stage2_33[96],stage2_32[102]}
   );
   gpc606_5 gpc6572 (
      {stage1_32[380], stage1_32[381], stage1_32[382], stage1_32[383], stage1_32[384], stage1_32[385]},
      {stage1_34[186], stage1_34[187], stage1_34[188], stage1_34[189], stage1_34[190], stage1_34[191]},
      {stage2_36[31],stage2_35[58],stage2_34[85],stage2_33[97],stage2_32[103]}
   );
   gpc606_5 gpc6573 (
      {stage1_32[386], stage1_32[387], stage1_32[388], stage1_32[389], stage1_32[390], stage1_32[391]},
      {stage1_34[192], stage1_34[193], stage1_34[194], stage1_34[195], stage1_34[196], stage1_34[197]},
      {stage2_36[32],stage2_35[59],stage2_34[86],stage2_33[98],stage2_32[104]}
   );
   gpc606_5 gpc6574 (
      {stage1_32[392], stage1_32[393], stage1_32[394], stage1_32[395], stage1_32[396], stage1_32[397]},
      {stage1_34[198], stage1_34[199], stage1_34[200], stage1_34[201], stage1_34[202], stage1_34[203]},
      {stage2_36[33],stage2_35[60],stage2_34[87],stage2_33[99],stage2_32[105]}
   );
   gpc606_5 gpc6575 (
      {stage1_32[398], stage1_32[399], stage1_32[400], stage1_32[401], stage1_32[402], stage1_32[403]},
      {stage1_34[204], stage1_34[205], stage1_34[206], stage1_34[207], stage1_34[208], stage1_34[209]},
      {stage2_36[34],stage2_35[61],stage2_34[88],stage2_33[100],stage2_32[106]}
   );
   gpc606_5 gpc6576 (
      {stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168], stage1_33[169]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[35],stage2_35[62],stage2_34[89],stage2_33[101]}
   );
   gpc606_5 gpc6577 (
      {stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174], stage1_33[175]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[36],stage2_35[63],stage2_34[90],stage2_33[102]}
   );
   gpc606_5 gpc6578 (
      {stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180], stage1_33[181]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[37],stage2_35[64],stage2_34[91],stage2_33[103]}
   );
   gpc606_5 gpc6579 (
      {stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186], stage1_33[187]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[38],stage2_35[65],stage2_34[92],stage2_33[104]}
   );
   gpc606_5 gpc6580 (
      {stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192], stage1_33[193]},
      {stage1_35[24], stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29]},
      {stage2_37[4],stage2_36[39],stage2_35[66],stage2_34[93],stage2_33[105]}
   );
   gpc606_5 gpc6581 (
      {stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198], stage1_33[199]},
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage2_37[5],stage2_36[40],stage2_35[67],stage2_34[94],stage2_33[106]}
   );
   gpc615_5 gpc6582 (
      {stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage1_34[210]},
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage2_37[6],stage2_36[41],stage2_35[68],stage2_34[95],stage2_33[107]}
   );
   gpc615_5 gpc6583 (
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209]},
      {stage1_34[211]},
      {stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage2_37[7],stage2_36[42],stage2_35[69],stage2_34[96],stage2_33[108]}
   );
   gpc606_5 gpc6584 (
      {stage1_34[212], stage1_34[213], stage1_34[214], stage1_34[215], stage1_34[216], stage1_34[217]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[8],stage2_36[43],stage2_35[70],stage2_34[97]}
   );
   gpc606_5 gpc6585 (
      {stage1_34[218], stage1_34[219], stage1_34[220], stage1_34[221], stage1_34[222], stage1_34[223]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[9],stage2_36[44],stage2_35[71],stage2_34[98]}
   );
   gpc606_5 gpc6586 (
      {stage1_34[224], stage1_34[225], stage1_34[226], stage1_34[227], stage1_34[228], stage1_34[229]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[10],stage2_36[45],stage2_35[72],stage2_34[99]}
   );
   gpc606_5 gpc6587 (
      {stage1_34[230], stage1_34[231], stage1_34[232], stage1_34[233], stage1_34[234], stage1_34[235]},
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23]},
      {stage2_38[3],stage2_37[11],stage2_36[46],stage2_35[73],stage2_34[100]}
   );
   gpc606_5 gpc6588 (
      {stage1_34[236], stage1_34[237], stage1_34[238], stage1_34[239], stage1_34[240], stage1_34[241]},
      {stage1_36[24], stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29]},
      {stage2_38[4],stage2_37[12],stage2_36[47],stage2_35[74],stage2_34[101]}
   );
   gpc615_5 gpc6589 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[30]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[5],stage2_37[13],stage2_36[48],stage2_35[75]}
   );
   gpc615_5 gpc6590 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[31]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[6],stage2_37[14],stage2_36[49],stage2_35[76]}
   );
   gpc615_5 gpc6591 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[32]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[7],stage2_37[15],stage2_36[50],stage2_35[77]}
   );
   gpc615_5 gpc6592 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[33]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[8],stage2_37[16],stage2_36[51],stage2_35[78]}
   );
   gpc615_5 gpc6593 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[34]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[9],stage2_37[17],stage2_36[52],stage2_35[79]}
   );
   gpc615_5 gpc6594 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[35]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[10],stage2_37[18],stage2_36[53],stage2_35[80]}
   );
   gpc615_5 gpc6595 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[36]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[11],stage2_37[19],stage2_36[54],stage2_35[81]}
   );
   gpc615_5 gpc6596 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[37]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[12],stage2_37[20],stage2_36[55],stage2_35[82]}
   );
   gpc615_5 gpc6597 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[38]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[13],stage2_37[21],stage2_36[56],stage2_35[83]}
   );
   gpc615_5 gpc6598 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[39]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[14],stage2_37[22],stage2_36[57],stage2_35[84]}
   );
   gpc615_5 gpc6599 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[40]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[15],stage2_37[23],stage2_36[58],stage2_35[85]}
   );
   gpc615_5 gpc6600 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[41]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[16],stage2_37[24],stage2_36[59],stage2_35[86]}
   );
   gpc615_5 gpc6601 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[42]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[17],stage2_37[25],stage2_36[60],stage2_35[87]}
   );
   gpc615_5 gpc6602 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[43]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[18],stage2_37[26],stage2_36[61],stage2_35[88]}
   );
   gpc615_5 gpc6603 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[44]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[19],stage2_37[27],stage2_36[62],stage2_35[89]}
   );
   gpc615_5 gpc6604 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[45]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[20],stage2_37[28],stage2_36[63],stage2_35[90]}
   );
   gpc615_5 gpc6605 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[46]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[21],stage2_37[29],stage2_36[64],stage2_35[91]}
   );
   gpc615_5 gpc6606 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[47]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[22],stage2_37[30],stage2_36[65],stage2_35[92]}
   );
   gpc615_5 gpc6607 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[48]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[23],stage2_37[31],stage2_36[66],stage2_35[93]}
   );
   gpc615_5 gpc6608 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[49]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[24],stage2_37[32],stage2_36[67],stage2_35[94]}
   );
   gpc615_5 gpc6609 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[50]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[25],stage2_37[33],stage2_36[68],stage2_35[95]}
   );
   gpc615_5 gpc6610 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[51]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[26],stage2_37[34],stage2_36[69],stage2_35[96]}
   );
   gpc615_5 gpc6611 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[52]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[27],stage2_37[35],stage2_36[70],stage2_35[97]}
   );
   gpc615_5 gpc6612 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[53]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[28],stage2_37[36],stage2_36[71],stage2_35[98]}
   );
   gpc615_5 gpc6613 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[54]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[29],stage2_37[37],stage2_36[72],stage2_35[99]}
   );
   gpc1163_5 gpc6614 (
      {stage1_36[55], stage1_36[56], stage1_36[57]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage1_38[0]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[25],stage2_38[30],stage2_37[38],stage2_36[73]}
   );
   gpc606_5 gpc6615 (
      {stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61], stage1_36[62], stage1_36[63]},
      {stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6]},
      {stage2_40[1],stage2_39[26],stage2_38[31],stage2_37[39],stage2_36[74]}
   );
   gpc606_5 gpc6616 (
      {stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67], stage1_36[68], stage1_36[69]},
      {stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12]},
      {stage2_40[2],stage2_39[27],stage2_38[32],stage2_37[40],stage2_36[75]}
   );
   gpc606_5 gpc6617 (
      {stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73], stage1_36[74], stage1_36[75]},
      {stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18]},
      {stage2_40[3],stage2_39[28],stage2_38[33],stage2_37[41],stage2_36[76]}
   );
   gpc606_5 gpc6618 (
      {stage1_36[76], stage1_36[77], stage1_36[78], stage1_36[79], stage1_36[80], stage1_36[81]},
      {stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24]},
      {stage2_40[4],stage2_39[29],stage2_38[34],stage2_37[42],stage2_36[77]}
   );
   gpc606_5 gpc6619 (
      {stage1_36[82], stage1_36[83], stage1_36[84], stage1_36[85], stage1_36[86], stage1_36[87]},
      {stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30]},
      {stage2_40[5],stage2_39[30],stage2_38[35],stage2_37[43],stage2_36[78]}
   );
   gpc606_5 gpc6620 (
      {stage1_36[88], stage1_36[89], stage1_36[90], stage1_36[91], stage1_36[92], stage1_36[93]},
      {stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36]},
      {stage2_40[6],stage2_39[31],stage2_38[36],stage2_37[44],stage2_36[79]}
   );
   gpc606_5 gpc6621 (
      {stage1_36[94], stage1_36[95], stage1_36[96], stage1_36[97], stage1_36[98], stage1_36[99]},
      {stage1_38[37], stage1_38[38], stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42]},
      {stage2_40[7],stage2_39[32],stage2_38[37],stage2_37[45],stage2_36[80]}
   );
   gpc606_5 gpc6622 (
      {stage1_36[100], stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105]},
      {stage1_38[43], stage1_38[44], stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48]},
      {stage2_40[8],stage2_39[33],stage2_38[38],stage2_37[46],stage2_36[81]}
   );
   gpc606_5 gpc6623 (
      {stage1_36[106], stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111]},
      {stage1_38[49], stage1_38[50], stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54]},
      {stage2_40[9],stage2_39[34],stage2_38[39],stage2_37[47],stage2_36[82]}
   );
   gpc606_5 gpc6624 (
      {stage1_36[112], stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117]},
      {stage1_38[55], stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage2_40[10],stage2_39[35],stage2_38[40],stage2_37[48],stage2_36[83]}
   );
   gpc606_5 gpc6625 (
      {stage1_36[118], stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123]},
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65], stage1_38[66]},
      {stage2_40[11],stage2_39[36],stage2_38[41],stage2_37[49],stage2_36[84]}
   );
   gpc606_5 gpc6626 (
      {stage1_36[124], stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129]},
      {stage1_38[67], stage1_38[68], stage1_38[69], stage1_38[70], stage1_38[71], stage1_38[72]},
      {stage2_40[12],stage2_39[37],stage2_38[42],stage2_37[50],stage2_36[85]}
   );
   gpc606_5 gpc6627 (
      {stage1_36[130], stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135]},
      {stage1_38[73], stage1_38[74], stage1_38[75], stage1_38[76], stage1_38[77], stage1_38[78]},
      {stage2_40[13],stage2_39[38],stage2_38[43],stage2_37[51],stage2_36[86]}
   );
   gpc606_5 gpc6628 (
      {stage1_36[136], stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141]},
      {stage1_38[79], stage1_38[80], stage1_38[81], stage1_38[82], stage1_38[83], stage1_38[84]},
      {stage2_40[14],stage2_39[39],stage2_38[44],stage2_37[52],stage2_36[87]}
   );
   gpc606_5 gpc6629 (
      {stage1_36[142], stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147]},
      {stage1_38[85], stage1_38[86], stage1_38[87], stage1_38[88], stage1_38[89], stage1_38[90]},
      {stage2_40[15],stage2_39[40],stage2_38[45],stage2_37[53],stage2_36[88]}
   );
   gpc606_5 gpc6630 (
      {stage1_36[148], stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153]},
      {stage1_38[91], stage1_38[92], stage1_38[93], stage1_38[94], stage1_38[95], stage1_38[96]},
      {stage2_40[16],stage2_39[41],stage2_38[46],stage2_37[54],stage2_36[89]}
   );
   gpc606_5 gpc6631 (
      {stage1_36[154], stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159]},
      {stage1_38[97], stage1_38[98], stage1_38[99], stage1_38[100], stage1_38[101], stage1_38[102]},
      {stage2_40[17],stage2_39[42],stage2_38[47],stage2_37[55],stage2_36[90]}
   );
   gpc606_5 gpc6632 (
      {stage1_36[160], stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165]},
      {stage1_38[103], stage1_38[104], stage1_38[105], stage1_38[106], stage1_38[107], stage1_38[108]},
      {stage2_40[18],stage2_39[43],stage2_38[48],stage2_37[56],stage2_36[91]}
   );
   gpc606_5 gpc6633 (
      {stage1_36[166], stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171]},
      {stage1_38[109], stage1_38[110], stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114]},
      {stage2_40[19],stage2_39[44],stage2_38[49],stage2_37[57],stage2_36[92]}
   );
   gpc606_5 gpc6634 (
      {stage1_36[172], stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177]},
      {stage1_38[115], stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage2_40[20],stage2_39[45],stage2_38[50],stage2_37[58],stage2_36[93]}
   );
   gpc606_5 gpc6635 (
      {stage1_36[178], stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183]},
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125], stage1_38[126]},
      {stage2_40[21],stage2_39[46],stage2_38[51],stage2_37[59],stage2_36[94]}
   );
   gpc606_5 gpc6636 (
      {stage1_36[184], stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189]},
      {stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130], stage1_38[131], stage1_38[132]},
      {stage2_40[22],stage2_39[47],stage2_38[52],stage2_37[60],stage2_36[95]}
   );
   gpc606_5 gpc6637 (
      {stage1_36[190], stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195]},
      {stage1_38[133], stage1_38[134], stage1_38[135], stage1_38[136], stage1_38[137], stage1_38[138]},
      {stage2_40[23],stage2_39[48],stage2_38[53],stage2_37[61],stage2_36[96]}
   );
   gpc606_5 gpc6638 (
      {stage1_36[196], stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201]},
      {stage1_38[139], stage1_38[140], stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144]},
      {stage2_40[24],stage2_39[49],stage2_38[54],stage2_37[62],stage2_36[97]}
   );
   gpc606_5 gpc6639 (
      {stage1_36[202], stage1_36[203], stage1_36[204], stage1_36[205], stage1_36[206], stage1_36[207]},
      {stage1_38[145], stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage2_40[25],stage2_39[50],stage2_38[55],stage2_37[63],stage2_36[98]}
   );
   gpc606_5 gpc6640 (
      {stage1_36[208], stage1_36[209], stage1_36[210], stage1_36[211], stage1_36[212], stage1_36[213]},
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155], stage1_38[156]},
      {stage2_40[26],stage2_39[51],stage2_38[56],stage2_37[64],stage2_36[99]}
   );
   gpc606_5 gpc6641 (
      {stage1_36[214], stage1_36[215], stage1_36[216], stage1_36[217], stage1_36[218], stage1_36[219]},
      {stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160], stage1_38[161], stage1_38[162]},
      {stage2_40[27],stage2_39[52],stage2_38[57],stage2_37[65],stage2_36[100]}
   );
   gpc606_5 gpc6642 (
      {stage1_36[220], stage1_36[221], stage1_36[222], stage1_36[223], stage1_36[224], stage1_36[225]},
      {stage1_38[163], stage1_38[164], stage1_38[165], stage1_38[166], stage1_38[167], stage1_38[168]},
      {stage2_40[28],stage2_39[53],stage2_38[58],stage2_37[66],stage2_36[101]}
   );
   gpc606_5 gpc6643 (
      {stage1_36[226], stage1_36[227], stage1_36[228], stage1_36[229], stage1_36[230], stage1_36[231]},
      {stage1_38[169], stage1_38[170], stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174]},
      {stage2_40[29],stage2_39[54],stage2_38[59],stage2_37[67],stage2_36[102]}
   );
   gpc606_5 gpc6644 (
      {stage1_36[232], stage1_36[233], stage1_36[234], stage1_36[235], stage1_36[236], stage1_36[237]},
      {stage1_38[175], stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage2_40[30],stage2_39[55],stage2_38[60],stage2_37[68],stage2_36[103]}
   );
   gpc606_5 gpc6645 (
      {stage1_36[238], stage1_36[239], stage1_36[240], stage1_36[241], stage1_36[242], stage1_36[243]},
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185], stage1_38[186]},
      {stage2_40[31],stage2_39[56],stage2_38[61],stage2_37[69],stage2_36[104]}
   );
   gpc606_5 gpc6646 (
      {stage1_36[244], stage1_36[245], stage1_36[246], stage1_36[247], stage1_36[248], stage1_36[249]},
      {stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190], stage1_38[191], stage1_38[192]},
      {stage2_40[32],stage2_39[57],stage2_38[62],stage2_37[70],stage2_36[105]}
   );
   gpc606_5 gpc6647 (
      {stage1_36[250], stage1_36[251], stage1_36[252], stage1_36[253], stage1_36[254], stage1_36[255]},
      {stage1_38[193], stage1_38[194], stage1_38[195], stage1_38[196], stage1_38[197], stage1_38[198]},
      {stage2_40[33],stage2_39[58],stage2_38[63],stage2_37[71],stage2_36[106]}
   );
   gpc606_5 gpc6648 (
      {stage1_36[256], stage1_36[257], stage1_36[258], stage1_36[259], stage1_36[260], stage1_36[261]},
      {stage1_38[199], stage1_38[200], stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204]},
      {stage2_40[34],stage2_39[59],stage2_38[64],stage2_37[72],stage2_36[107]}
   );
   gpc606_5 gpc6649 (
      {stage1_36[262], stage1_36[263], stage1_36[264], stage1_36[265], stage1_36[266], stage1_36[267]},
      {stage1_38[205], stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage2_40[35],stage2_39[60],stage2_38[65],stage2_37[73],stage2_36[108]}
   );
   gpc606_5 gpc6650 (
      {stage1_36[268], stage1_36[269], stage1_36[270], stage1_36[271], stage1_36[272], stage1_36[273]},
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215], stage1_38[216]},
      {stage2_40[36],stage2_39[61],stage2_38[66],stage2_37[74],stage2_36[109]}
   );
   gpc606_5 gpc6651 (
      {stage1_36[274], stage1_36[275], stage1_36[276], stage1_36[277], stage1_36[278], stage1_36[279]},
      {stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220], stage1_38[221], stage1_38[222]},
      {stage2_40[37],stage2_39[62],stage2_38[67],stage2_37[75],stage2_36[110]}
   );
   gpc606_5 gpc6652 (
      {stage1_36[280], stage1_36[281], stage1_36[282], stage1_36[283], stage1_36[284], stage1_36[285]},
      {stage1_38[223], stage1_38[224], stage1_38[225], stage1_38[226], stage1_38[227], stage1_38[228]},
      {stage2_40[38],stage2_39[63],stage2_38[68],stage2_37[76],stage2_36[111]}
   );
   gpc606_5 gpc6653 (
      {stage1_36[286], stage1_36[287], stage1_36[288], stage1_36[289], stage1_36[290], stage1_36[291]},
      {stage1_38[229], stage1_38[230], stage1_38[231], stage1_38[232], stage1_38[233], stage1_38[234]},
      {stage2_40[39],stage2_39[64],stage2_38[69],stage2_37[77],stage2_36[112]}
   );
   gpc606_5 gpc6654 (
      {stage1_36[292], stage1_36[293], stage1_36[294], stage1_36[295], stage1_36[296], stage1_36[297]},
      {stage1_38[235], stage1_38[236], stage1_38[237], stage1_38[238], stage1_38[239], stage1_38[240]},
      {stage2_40[40],stage2_39[65],stage2_38[70],stage2_37[78],stage2_36[113]}
   );
   gpc606_5 gpc6655 (
      {stage1_36[298], stage1_36[299], stage1_36[300], stage1_36[301], stage1_36[302], stage1_36[303]},
      {stage1_38[241], stage1_38[242], stage1_38[243], stage1_38[244], stage1_38[245], stage1_38[246]},
      {stage2_40[41],stage2_39[66],stage2_38[71],stage2_37[79],stage2_36[114]}
   );
   gpc606_5 gpc6656 (
      {stage1_36[304], stage1_36[305], stage1_36[306], stage1_36[307], stage1_36[308], stage1_36[309]},
      {stage1_38[247], stage1_38[248], stage1_38[249], stage1_38[250], stage1_38[251], stage1_38[252]},
      {stage2_40[42],stage2_39[67],stage2_38[72],stage2_37[80],stage2_36[115]}
   );
   gpc606_5 gpc6657 (
      {stage1_36[310], stage1_36[311], stage1_36[312], stage1_36[313], stage1_36[314], stage1_36[315]},
      {stage1_38[253], stage1_38[254], stage1_38[255], stage1_38[256], stage1_38[257], stage1_38[258]},
      {stage2_40[43],stage2_39[68],stage2_38[73],stage2_37[81],stage2_36[116]}
   );
   gpc615_5 gpc6658 (
      {stage1_36[316], stage1_36[317], stage1_36[318], stage1_36[319], stage1_36[320]},
      {stage1_37[156]},
      {stage1_38[259], stage1_38[260], stage1_38[261], stage1_38[262], stage1_38[263], stage1_38[264]},
      {stage2_40[44],stage2_39[69],stage2_38[74],stage2_37[82],stage2_36[117]}
   );
   gpc615_5 gpc6659 (
      {stage1_36[321], stage1_36[322], stage1_36[323], stage1_36[324], stage1_36[325]},
      {stage1_37[157]},
      {stage1_38[265], stage1_38[266], stage1_38[267], stage1_38[268], stage1_38[269], stage1_38[270]},
      {stage2_40[45],stage2_39[70],stage2_38[75],stage2_37[83],stage2_36[118]}
   );
   gpc615_5 gpc6660 (
      {stage1_36[326], stage1_36[327], stage1_36[328], stage1_36[329], stage1_36[330]},
      {stage1_37[158]},
      {stage1_38[271], stage1_38[272], stage1_38[273], stage1_38[274], stage1_38[275], stage1_38[276]},
      {stage2_40[46],stage2_39[71],stage2_38[76],stage2_37[84],stage2_36[119]}
   );
   gpc606_5 gpc6661 (
      {stage1_37[159], stage1_37[160], stage1_37[161], stage1_37[162], stage1_37[163], stage1_37[164]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[47],stage2_39[72],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc6662 (
      {stage1_37[165], stage1_37[166], stage1_37[167], stage1_37[168], stage1_37[169], stage1_37[170]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[48],stage2_39[73],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc6663 (
      {stage1_37[171], stage1_37[172], stage1_37[173], stage1_37[174], stage1_37[175], stage1_37[176]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[49],stage2_39[74],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc6664 (
      {stage1_37[177], stage1_37[178], stage1_37[179], stage1_37[180], stage1_37[181], stage1_37[182]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[50],stage2_39[75],stage2_38[80],stage2_37[88]}
   );
   gpc606_5 gpc6665 (
      {stage1_37[183], stage1_37[184], stage1_37[185], stage1_37[186], stage1_37[187], stage1_37[188]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[51],stage2_39[76],stage2_38[81],stage2_37[89]}
   );
   gpc606_5 gpc6666 (
      {stage1_37[189], stage1_37[190], stage1_37[191], stage1_37[192], stage1_37[193], stage1_37[194]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[52],stage2_39[77],stage2_38[82],stage2_37[90]}
   );
   gpc606_5 gpc6667 (
      {stage1_37[195], stage1_37[196], stage1_37[197], stage1_37[198], stage1_37[199], stage1_37[200]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[53],stage2_39[78],stage2_38[83],stage2_37[91]}
   );
   gpc606_5 gpc6668 (
      {stage1_37[201], stage1_37[202], stage1_37[203], stage1_37[204], stage1_37[205], stage1_37[206]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[54],stage2_39[79],stage2_38[84],stage2_37[92]}
   );
   gpc606_5 gpc6669 (
      {stage1_37[207], stage1_37[208], stage1_37[209], stage1_37[210], stage1_37[211], stage1_37[212]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[55],stage2_39[80],stage2_38[85],stage2_37[93]}
   );
   gpc606_5 gpc6670 (
      {stage1_37[213], stage1_37[214], stage1_37[215], stage1_37[216], stage1_37[217], stage1_37[218]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[56],stage2_39[81],stage2_38[86],stage2_37[94]}
   );
   gpc606_5 gpc6671 (
      {stage1_37[219], stage1_37[220], stage1_37[221], stage1_37[222], stage1_37[223], stage1_37[224]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[57],stage2_39[82],stage2_38[87],stage2_37[95]}
   );
   gpc606_5 gpc6672 (
      {stage1_37[225], stage1_37[226], stage1_37[227], stage1_37[228], stage1_37[229], stage1_37[230]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[58],stage2_39[83],stage2_38[88],stage2_37[96]}
   );
   gpc606_5 gpc6673 (
      {stage1_37[231], stage1_37[232], stage1_37[233], stage1_37[234], stage1_37[235], stage1_37[236]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[59],stage2_39[84],stage2_38[89],stage2_37[97]}
   );
   gpc606_5 gpc6674 (
      {stage1_37[237], stage1_37[238], stage1_37[239], stage1_37[240], stage1_37[241], stage1_37[242]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[60],stage2_39[85],stage2_38[90],stage2_37[98]}
   );
   gpc606_5 gpc6675 (
      {stage1_37[243], stage1_37[244], stage1_37[245], stage1_37[246], stage1_37[247], stage1_37[248]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[61],stage2_39[86],stage2_38[91],stage2_37[99]}
   );
   gpc606_5 gpc6676 (
      {stage1_37[249], stage1_37[250], stage1_37[251], stage1_37[252], stage1_37[253], stage1_37[254]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[62],stage2_39[87],stage2_38[92],stage2_37[100]}
   );
   gpc606_5 gpc6677 (
      {stage1_37[255], stage1_37[256], stage1_37[257], stage1_37[258], stage1_37[259], stage1_37[260]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[63],stage2_39[88],stage2_38[93],stage2_37[101]}
   );
   gpc606_5 gpc6678 (
      {stage1_37[261], stage1_37[262], stage1_37[263], stage1_37[264], stage1_37[265], stage1_37[266]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[64],stage2_39[89],stage2_38[94],stage2_37[102]}
   );
   gpc606_5 gpc6679 (
      {stage1_37[267], stage1_37[268], stage1_37[269], stage1_37[270], stage1_37[271], stage1_37[272]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[65],stage2_39[90],stage2_38[95],stage2_37[103]}
   );
   gpc606_5 gpc6680 (
      {stage1_37[273], stage1_37[274], stage1_37[275], stage1_37[276], stage1_37[277], stage1_37[278]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[66],stage2_39[91],stage2_38[96],stage2_37[104]}
   );
   gpc606_5 gpc6681 (
      {stage1_37[279], stage1_37[280], stage1_37[281], stage1_37[282], stage1_37[283], stage1_37[284]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[67],stage2_39[92],stage2_38[97],stage2_37[105]}
   );
   gpc606_5 gpc6682 (
      {stage1_37[285], stage1_37[286], stage1_37[287], stage1_37[288], stage1_37[289], stage1_37[290]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[68],stage2_39[93],stage2_38[98],stage2_37[106]}
   );
   gpc606_5 gpc6683 (
      {stage1_37[291], stage1_37[292], stage1_37[293], stage1_37[294], stage1_37[295], stage1_37[296]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[69],stage2_39[94],stage2_38[99],stage2_37[107]}
   );
   gpc606_5 gpc6684 (
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[0],stage2_41[23],stage2_40[70],stage2_39[95]}
   );
   gpc606_5 gpc6685 (
      {stage1_39[145], stage1_39[146], stage1_39[147], stage1_39[148], stage1_39[149], stage1_39[150]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage2_43[1],stage2_42[1],stage2_41[24],stage2_40[71],stage2_39[96]}
   );
   gpc606_5 gpc6686 (
      {stage1_39[151], stage1_39[152], stage1_39[153], stage1_39[154], stage1_39[155], stage1_39[156]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage2_43[2],stage2_42[2],stage2_41[25],stage2_40[72],stage2_39[97]}
   );
   gpc606_5 gpc6687 (
      {stage1_39[157], stage1_39[158], stage1_39[159], stage1_39[160], stage1_39[161], stage1_39[162]},
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage2_43[3],stage2_42[3],stage2_41[26],stage2_40[73],stage2_39[98]}
   );
   gpc606_5 gpc6688 (
      {stage1_39[163], stage1_39[164], stage1_39[165], stage1_39[166], stage1_39[167], stage1_39[168]},
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage2_43[4],stage2_42[4],stage2_41[27],stage2_40[74],stage2_39[99]}
   );
   gpc615_5 gpc6689 (
      {stage1_39[169], stage1_39[170], stage1_39[171], stage1_39[172], stage1_39[173]},
      {stage1_40[0]},
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage2_43[5],stage2_42[5],stage2_41[28],stage2_40[75],stage2_39[100]}
   );
   gpc615_5 gpc6690 (
      {stage1_39[174], stage1_39[175], stage1_39[176], stage1_39[177], stage1_39[178]},
      {stage1_40[1]},
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage2_43[6],stage2_42[6],stage2_41[29],stage2_40[76],stage2_39[101]}
   );
   gpc615_5 gpc6691 (
      {stage1_39[179], stage1_39[180], stage1_39[181], stage1_39[182], stage1_39[183]},
      {stage1_40[2]},
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage2_43[7],stage2_42[7],stage2_41[30],stage2_40[77],stage2_39[102]}
   );
   gpc615_5 gpc6692 (
      {stage1_39[184], stage1_39[185], stage1_39[186], stage1_39[187], stage1_39[188]},
      {stage1_40[3]},
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52], stage1_41[53]},
      {stage2_43[8],stage2_42[8],stage2_41[31],stage2_40[78],stage2_39[103]}
   );
   gpc615_5 gpc6693 (
      {stage1_39[189], stage1_39[190], stage1_39[191], stage1_39[192], stage1_39[193]},
      {stage1_40[4]},
      {stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57], stage1_41[58], stage1_41[59]},
      {stage2_43[9],stage2_42[9],stage2_41[32],stage2_40[79],stage2_39[104]}
   );
   gpc606_5 gpc6694 (
      {stage1_40[5], stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[10],stage2_42[10],stage2_41[33],stage2_40[80]}
   );
   gpc606_5 gpc6695 (
      {stage1_40[11], stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[11],stage2_42[11],stage2_41[34],stage2_40[81]}
   );
   gpc606_5 gpc6696 (
      {stage1_40[17], stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[12],stage2_42[12],stage2_41[35],stage2_40[82]}
   );
   gpc606_5 gpc6697 (
      {stage1_40[23], stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[13],stage2_42[13],stage2_41[36],stage2_40[83]}
   );
   gpc606_5 gpc6698 (
      {stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[14],stage2_42[14],stage2_41[37],stage2_40[84]}
   );
   gpc606_5 gpc6699 (
      {stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[15],stage2_42[15],stage2_41[38],stage2_40[85]}
   );
   gpc606_5 gpc6700 (
      {stage1_40[41], stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[16],stage2_42[16],stage2_41[39],stage2_40[86]}
   );
   gpc606_5 gpc6701 (
      {stage1_40[47], stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[17],stage2_42[17],stage2_41[40],stage2_40[87]}
   );
   gpc606_5 gpc6702 (
      {stage1_40[53], stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[18],stage2_42[18],stage2_41[41],stage2_40[88]}
   );
   gpc606_5 gpc6703 (
      {stage1_40[59], stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[19],stage2_42[19],stage2_41[42],stage2_40[89]}
   );
   gpc606_5 gpc6704 (
      {stage1_40[65], stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[20],stage2_42[20],stage2_41[43],stage2_40[90]}
   );
   gpc606_5 gpc6705 (
      {stage1_40[71], stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[21],stage2_42[21],stage2_41[44],stage2_40[91]}
   );
   gpc606_5 gpc6706 (
      {stage1_40[77], stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[22],stage2_42[22],stage2_41[45],stage2_40[92]}
   );
   gpc606_5 gpc6707 (
      {stage1_40[83], stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[23],stage2_42[23],stage2_41[46],stage2_40[93]}
   );
   gpc606_5 gpc6708 (
      {stage1_40[89], stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[24],stage2_42[24],stage2_41[47],stage2_40[94]}
   );
   gpc606_5 gpc6709 (
      {stage1_40[95], stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[25],stage2_42[25],stage2_41[48],stage2_40[95]}
   );
   gpc606_5 gpc6710 (
      {stage1_40[101], stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[26],stage2_42[26],stage2_41[49],stage2_40[96]}
   );
   gpc606_5 gpc6711 (
      {stage1_40[107], stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[27],stage2_42[27],stage2_41[50],stage2_40[97]}
   );
   gpc606_5 gpc6712 (
      {stage1_40[113], stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[28],stage2_42[28],stage2_41[51],stage2_40[98]}
   );
   gpc606_5 gpc6713 (
      {stage1_40[119], stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[29],stage2_42[29],stage2_41[52],stage2_40[99]}
   );
   gpc606_5 gpc6714 (
      {stage1_40[125], stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[30],stage2_42[30],stage2_41[53],stage2_40[100]}
   );
   gpc606_5 gpc6715 (
      {stage1_40[131], stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[31],stage2_42[31],stage2_41[54],stage2_40[101]}
   );
   gpc606_5 gpc6716 (
      {stage1_40[137], stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[32],stage2_42[32],stage2_41[55],stage2_40[102]}
   );
   gpc606_5 gpc6717 (
      {stage1_40[143], stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148]},
      {stage1_42[138], stage1_42[139], stage1_42[140], stage1_42[141], stage1_42[142], stage1_42[143]},
      {stage2_44[23],stage2_43[33],stage2_42[33],stage2_41[56],stage2_40[103]}
   );
   gpc606_5 gpc6718 (
      {stage1_40[149], stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154]},
      {stage1_42[144], stage1_42[145], stage1_42[146], stage1_42[147], stage1_42[148], stage1_42[149]},
      {stage2_44[24],stage2_43[34],stage2_42[34],stage2_41[57],stage2_40[104]}
   );
   gpc606_5 gpc6719 (
      {stage1_40[155], stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160]},
      {stage1_42[150], stage1_42[151], stage1_42[152], stage1_42[153], stage1_42[154], stage1_42[155]},
      {stage2_44[25],stage2_43[35],stage2_42[35],stage2_41[58],stage2_40[105]}
   );
   gpc606_5 gpc6720 (
      {stage1_40[161], stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166]},
      {stage1_42[156], stage1_42[157], stage1_42[158], stage1_42[159], stage1_42[160], stage1_42[161]},
      {stage2_44[26],stage2_43[36],stage2_42[36],stage2_41[59],stage2_40[106]}
   );
   gpc606_5 gpc6721 (
      {stage1_40[167], stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172]},
      {stage1_42[162], stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage2_44[27],stage2_43[37],stage2_42[37],stage2_41[60],stage2_40[107]}
   );
   gpc606_5 gpc6722 (
      {stage1_40[173], stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178]},
      {stage1_42[168], stage1_42[169], stage1_42[170], stage1_42[171], stage1_42[172], stage1_42[173]},
      {stage2_44[28],stage2_43[38],stage2_42[38],stage2_41[61],stage2_40[108]}
   );
   gpc606_5 gpc6723 (
      {stage1_40[179], stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184]},
      {stage1_42[174], stage1_42[175], stage1_42[176], stage1_42[177], stage1_42[178], stage1_42[179]},
      {stage2_44[29],stage2_43[39],stage2_42[39],stage2_41[62],stage2_40[109]}
   );
   gpc606_5 gpc6724 (
      {stage1_40[185], stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190]},
      {stage1_42[180], stage1_42[181], stage1_42[182], stage1_42[183], stage1_42[184], stage1_42[185]},
      {stage2_44[30],stage2_43[40],stage2_42[40],stage2_41[63],stage2_40[110]}
   );
   gpc606_5 gpc6725 (
      {stage1_40[191], stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196]},
      {stage1_42[186], stage1_42[187], stage1_42[188], stage1_42[189], stage1_42[190], stage1_42[191]},
      {stage2_44[31],stage2_43[41],stage2_42[41],stage2_41[64],stage2_40[111]}
   );
   gpc606_5 gpc6726 (
      {stage1_40[197], stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202]},
      {stage1_42[192], stage1_42[193], stage1_42[194], stage1_42[195], stage1_42[196], stage1_42[197]},
      {stage2_44[32],stage2_43[42],stage2_42[42],stage2_41[65],stage2_40[112]}
   );
   gpc606_5 gpc6727 (
      {stage1_41[60], stage1_41[61], stage1_41[62], stage1_41[63], stage1_41[64], stage1_41[65]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[33],stage2_43[43],stage2_42[43],stage2_41[66]}
   );
   gpc606_5 gpc6728 (
      {stage1_41[66], stage1_41[67], stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[34],stage2_43[44],stage2_42[44],stage2_41[67]}
   );
   gpc606_5 gpc6729 (
      {stage1_41[72], stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[35],stage2_43[45],stage2_42[45],stage2_41[68]}
   );
   gpc606_5 gpc6730 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82], stage1_41[83]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[36],stage2_43[46],stage2_42[46],stage2_41[69]}
   );
   gpc606_5 gpc6731 (
      {stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87], stage1_41[88], stage1_41[89]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[37],stage2_43[47],stage2_42[47],stage2_41[70]}
   );
   gpc606_5 gpc6732 (
      {stage1_41[90], stage1_41[91], stage1_41[92], stage1_41[93], stage1_41[94], stage1_41[95]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[38],stage2_43[48],stage2_42[48],stage2_41[71]}
   );
   gpc606_5 gpc6733 (
      {stage1_41[96], stage1_41[97], stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[39],stage2_43[49],stage2_42[49],stage2_41[72]}
   );
   gpc606_5 gpc6734 (
      {stage1_41[102], stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[40],stage2_43[50],stage2_42[50],stage2_41[73]}
   );
   gpc606_5 gpc6735 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112], stage1_41[113]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[41],stage2_43[51],stage2_42[51],stage2_41[74]}
   );
   gpc606_5 gpc6736 (
      {stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117], stage1_41[118], stage1_41[119]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[42],stage2_43[52],stage2_42[52],stage2_41[75]}
   );
   gpc606_5 gpc6737 (
      {stage1_41[120], stage1_41[121], stage1_41[122], stage1_41[123], stage1_41[124], stage1_41[125]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[43],stage2_43[53],stage2_42[53],stage2_41[76]}
   );
   gpc606_5 gpc6738 (
      {stage1_41[126], stage1_41[127], stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[44],stage2_43[54],stage2_42[54],stage2_41[77]}
   );
   gpc606_5 gpc6739 (
      {stage1_41[132], stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[45],stage2_43[55],stage2_42[55],stage2_41[78]}
   );
   gpc606_5 gpc6740 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142], stage1_41[143]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[46],stage2_43[56],stage2_42[56],stage2_41[79]}
   );
   gpc606_5 gpc6741 (
      {stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147], stage1_41[148], stage1_41[149]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[47],stage2_43[57],stage2_42[57],stage2_41[80]}
   );
   gpc606_5 gpc6742 (
      {stage1_41[150], stage1_41[151], stage1_41[152], stage1_41[153], stage1_41[154], stage1_41[155]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[48],stage2_43[58],stage2_42[58],stage2_41[81]}
   );
   gpc606_5 gpc6743 (
      {stage1_41[156], stage1_41[157], stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[49],stage2_43[59],stage2_42[59],stage2_41[82]}
   );
   gpc606_5 gpc6744 (
      {stage1_41[162], stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[50],stage2_43[60],stage2_42[60],stage2_41[83]}
   );
   gpc606_5 gpc6745 (
      {stage1_41[168], stage1_41[169], stage1_41[170], stage1_41[171], stage1_41[172], stage1_41[173]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[51],stage2_43[61],stage2_42[61],stage2_41[84]}
   );
   gpc606_5 gpc6746 (
      {stage1_41[174], stage1_41[175], stage1_41[176], stage1_41[177], stage1_41[178], stage1_41[179]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[52],stage2_43[62],stage2_42[62],stage2_41[85]}
   );
   gpc606_5 gpc6747 (
      {stage1_41[180], stage1_41[181], stage1_41[182], stage1_41[183], stage1_41[184], stage1_41[185]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[53],stage2_43[63],stage2_42[63],stage2_41[86]}
   );
   gpc606_5 gpc6748 (
      {stage1_41[186], stage1_41[187], stage1_41[188], stage1_41[189], stage1_41[190], stage1_41[191]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[54],stage2_43[64],stage2_42[64],stage2_41[87]}
   );
   gpc606_5 gpc6749 (
      {stage1_41[192], stage1_41[193], stage1_41[194], stage1_41[195], stage1_41[196], stage1_41[197]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[55],stage2_43[65],stage2_42[65],stage2_41[88]}
   );
   gpc606_5 gpc6750 (
      {stage1_41[198], stage1_41[199], stage1_41[200], stage1_41[201], stage1_41[202], stage1_41[203]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[56],stage2_43[66],stage2_42[66],stage2_41[89]}
   );
   gpc606_5 gpc6751 (
      {stage1_41[204], stage1_41[205], stage1_41[206], stage1_41[207], stage1_41[208], stage1_41[209]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[57],stage2_43[67],stage2_42[67],stage2_41[90]}
   );
   gpc606_5 gpc6752 (
      {stage1_41[210], stage1_41[211], stage1_41[212], stage1_41[213], stage1_41[214], stage1_41[215]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[58],stage2_43[68],stage2_42[68],stage2_41[91]}
   );
   gpc606_5 gpc6753 (
      {stage1_41[216], stage1_41[217], stage1_41[218], stage1_41[219], stage1_41[220], stage1_41[221]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[59],stage2_43[69],stage2_42[69],stage2_41[92]}
   );
   gpc606_5 gpc6754 (
      {stage1_41[222], stage1_41[223], stage1_41[224], stage1_41[225], stage1_41[226], stage1_41[227]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[60],stage2_43[70],stage2_42[70],stage2_41[93]}
   );
   gpc606_5 gpc6755 (
      {stage1_41[228], stage1_41[229], stage1_41[230], stage1_41[231], stage1_41[232], stage1_41[233]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[61],stage2_43[71],stage2_42[71],stage2_41[94]}
   );
   gpc606_5 gpc6756 (
      {stage1_41[234], stage1_41[235], stage1_41[236], stage1_41[237], stage1_41[238], stage1_41[239]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[62],stage2_43[72],stage2_42[72],stage2_41[95]}
   );
   gpc606_5 gpc6757 (
      {stage1_41[240], stage1_41[241], stage1_41[242], stage1_41[243], stage1_41[244], stage1_41[245]},
      {stage1_43[180], stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage2_45[30],stage2_44[63],stage2_43[73],stage2_42[73],stage2_41[96]}
   );
   gpc606_5 gpc6758 (
      {stage1_41[246], stage1_41[247], stage1_41[248], stage1_41[249], stage1_41[250], stage1_41[251]},
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190], stage1_43[191]},
      {stage2_45[31],stage2_44[64],stage2_43[74],stage2_42[74],stage2_41[97]}
   );
   gpc615_5 gpc6759 (
      {stage1_42[198], stage1_42[199], stage1_42[200], stage1_42[201], stage1_42[202]},
      {stage1_43[192]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[32],stage2_44[65],stage2_43[75],stage2_42[75]}
   );
   gpc615_5 gpc6760 (
      {stage1_42[203], stage1_42[204], stage1_42[205], stage1_42[206], stage1_42[207]},
      {stage1_43[193]},
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage2_46[1],stage2_45[33],stage2_44[66],stage2_43[76],stage2_42[76]}
   );
   gpc615_5 gpc6761 (
      {stage1_42[208], stage1_42[209], stage1_42[210], stage1_42[211], stage1_42[212]},
      {stage1_43[194]},
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage2_46[2],stage2_45[34],stage2_44[67],stage2_43[77],stage2_42[77]}
   );
   gpc615_5 gpc6762 (
      {stage1_42[213], stage1_42[214], stage1_42[215], stage1_42[216], stage1_42[217]},
      {stage1_43[195]},
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage2_46[3],stage2_45[35],stage2_44[68],stage2_43[78],stage2_42[78]}
   );
   gpc615_5 gpc6763 (
      {stage1_42[218], stage1_42[219], stage1_42[220], stage1_42[221], stage1_42[222]},
      {stage1_43[196]},
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage2_46[4],stage2_45[36],stage2_44[69],stage2_43[79],stage2_42[79]}
   );
   gpc615_5 gpc6764 (
      {stage1_42[223], stage1_42[224], stage1_42[225], stage1_42[226], stage1_42[227]},
      {stage1_43[197]},
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage2_46[5],stage2_45[37],stage2_44[70],stage2_43[80],stage2_42[80]}
   );
   gpc1415_5 gpc6765 (
      {stage1_43[198], stage1_43[199], stage1_43[200], stage1_43[201], stage1_43[202]},
      {stage1_44[36]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3]},
      {stage1_46[0]},
      {stage2_47[0],stage2_46[6],stage2_45[38],stage2_44[71],stage2_43[81]}
   );
   gpc1415_5 gpc6766 (
      {stage1_43[203], stage1_43[204], stage1_43[205], stage1_43[206], stage1_43[207]},
      {stage1_44[37]},
      {stage1_45[4], stage1_45[5], stage1_45[6], stage1_45[7]},
      {stage1_46[1]},
      {stage2_47[1],stage2_46[7],stage2_45[39],stage2_44[72],stage2_43[82]}
   );
   gpc1415_5 gpc6767 (
      {stage1_43[208], stage1_43[209], stage1_43[210], stage1_43[211], stage1_43[212]},
      {stage1_44[38]},
      {stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage1_46[2]},
      {stage2_47[2],stage2_46[8],stage2_45[40],stage2_44[73],stage2_43[83]}
   );
   gpc1415_5 gpc6768 (
      {stage1_43[213], stage1_43[214], stage1_43[215], stage1_43[216], stage1_43[217]},
      {stage1_44[39]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15]},
      {stage1_46[3]},
      {stage2_47[3],stage2_46[9],stage2_45[41],stage2_44[74],stage2_43[84]}
   );
   gpc606_5 gpc6769 (
      {stage1_44[40], stage1_44[41], stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45]},
      {stage1_46[4], stage1_46[5], stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9]},
      {stage2_48[0],stage2_47[4],stage2_46[10],stage2_45[42],stage2_44[75]}
   );
   gpc606_5 gpc6770 (
      {stage1_44[46], stage1_44[47], stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51]},
      {stage1_46[10], stage1_46[11], stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15]},
      {stage2_48[1],stage2_47[5],stage2_46[11],stage2_45[43],stage2_44[76]}
   );
   gpc606_5 gpc6771 (
      {stage1_44[52], stage1_44[53], stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57]},
      {stage1_46[16], stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage2_48[2],stage2_47[6],stage2_46[12],stage2_45[44],stage2_44[77]}
   );
   gpc606_5 gpc6772 (
      {stage1_44[58], stage1_44[59], stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63]},
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27]},
      {stage2_48[3],stage2_47[7],stage2_46[13],stage2_45[45],stage2_44[78]}
   );
   gpc606_5 gpc6773 (
      {stage1_44[64], stage1_44[65], stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69]},
      {stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33]},
      {stage2_48[4],stage2_47[8],stage2_46[14],stage2_45[46],stage2_44[79]}
   );
   gpc606_5 gpc6774 (
      {stage1_44[70], stage1_44[71], stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75]},
      {stage1_46[34], stage1_46[35], stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39]},
      {stage2_48[5],stage2_47[9],stage2_46[15],stage2_45[47],stage2_44[80]}
   );
   gpc606_5 gpc6775 (
      {stage1_44[76], stage1_44[77], stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81]},
      {stage1_46[40], stage1_46[41], stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45]},
      {stage2_48[6],stage2_47[10],stage2_46[16],stage2_45[48],stage2_44[81]}
   );
   gpc606_5 gpc6776 (
      {stage1_44[82], stage1_44[83], stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87]},
      {stage1_46[46], stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage2_48[7],stage2_47[11],stage2_46[17],stage2_45[49],stage2_44[82]}
   );
   gpc606_5 gpc6777 (
      {stage1_44[88], stage1_44[89], stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93]},
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57]},
      {stage2_48[8],stage2_47[12],stage2_46[18],stage2_45[50],stage2_44[83]}
   );
   gpc606_5 gpc6778 (
      {stage1_44[94], stage1_44[95], stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99]},
      {stage1_46[58], stage1_46[59], stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63]},
      {stage2_48[9],stage2_47[13],stage2_46[19],stage2_45[51],stage2_44[84]}
   );
   gpc606_5 gpc6779 (
      {stage1_44[100], stage1_44[101], stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105]},
      {stage1_46[64], stage1_46[65], stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69]},
      {stage2_48[10],stage2_47[14],stage2_46[20],stage2_45[52],stage2_44[85]}
   );
   gpc606_5 gpc6780 (
      {stage1_44[106], stage1_44[107], stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111]},
      {stage1_46[70], stage1_46[71], stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75]},
      {stage2_48[11],stage2_47[15],stage2_46[21],stage2_45[53],stage2_44[86]}
   );
   gpc606_5 gpc6781 (
      {stage1_44[112], stage1_44[113], stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117]},
      {stage1_46[76], stage1_46[77], stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81]},
      {stage2_48[12],stage2_47[16],stage2_46[22],stage2_45[54],stage2_44[87]}
   );
   gpc606_5 gpc6782 (
      {stage1_44[118], stage1_44[119], stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123]},
      {stage1_46[82], stage1_46[83], stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87]},
      {stage2_48[13],stage2_47[17],stage2_46[23],stage2_45[55],stage2_44[88]}
   );
   gpc615_5 gpc6783 (
      {stage1_44[124], stage1_44[125], stage1_44[126], stage1_44[127], stage1_44[128]},
      {stage1_45[16]},
      {stage1_46[88], stage1_46[89], stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93]},
      {stage2_48[14],stage2_47[18],stage2_46[24],stage2_45[56],stage2_44[89]}
   );
   gpc615_5 gpc6784 (
      {stage1_44[129], stage1_44[130], stage1_44[131], stage1_44[132], stage1_44[133]},
      {stage1_45[17]},
      {stage1_46[94], stage1_46[95], stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99]},
      {stage2_48[15],stage2_47[19],stage2_46[25],stage2_45[57],stage2_44[90]}
   );
   gpc615_5 gpc6785 (
      {stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137], stage1_44[138]},
      {stage1_45[18]},
      {stage1_46[100], stage1_46[101], stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105]},
      {stage2_48[16],stage2_47[20],stage2_46[26],stage2_45[58],stage2_44[91]}
   );
   gpc615_5 gpc6786 (
      {stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_45[19]},
      {stage1_46[106], stage1_46[107], stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111]},
      {stage2_48[17],stage2_47[21],stage2_46[27],stage2_45[59],stage2_44[92]}
   );
   gpc615_5 gpc6787 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148]},
      {stage1_45[20]},
      {stage1_46[112], stage1_46[113], stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117]},
      {stage2_48[18],stage2_47[22],stage2_46[28],stage2_45[60],stage2_44[93]}
   );
   gpc615_5 gpc6788 (
      {stage1_44[149], stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153]},
      {stage1_45[21]},
      {stage1_46[118], stage1_46[119], stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123]},
      {stage2_48[19],stage2_47[23],stage2_46[29],stage2_45[61],stage2_44[94]}
   );
   gpc615_5 gpc6789 (
      {stage1_44[154], stage1_44[155], stage1_44[156], stage1_44[157], stage1_44[158]},
      {stage1_45[22]},
      {stage1_46[124], stage1_46[125], stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129]},
      {stage2_48[20],stage2_47[24],stage2_46[30],stage2_45[62],stage2_44[95]}
   );
   gpc615_5 gpc6790 (
      {stage1_44[159], stage1_44[160], stage1_44[161], stage1_44[162], stage1_44[163]},
      {stage1_45[23]},
      {stage1_46[130], stage1_46[131], stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135]},
      {stage2_48[21],stage2_47[25],stage2_46[31],stage2_45[63],stage2_44[96]}
   );
   gpc615_5 gpc6791 (
      {stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167], stage1_44[168]},
      {stage1_45[24]},
      {stage1_46[136], stage1_46[137], stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141]},
      {stage2_48[22],stage2_47[26],stage2_46[32],stage2_45[64],stage2_44[97]}
   );
   gpc615_5 gpc6792 (
      {stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_45[25]},
      {stage1_46[142], stage1_46[143], stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147]},
      {stage2_48[23],stage2_47[27],stage2_46[33],stage2_45[65],stage2_44[98]}
   );
   gpc615_5 gpc6793 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178]},
      {stage1_45[26]},
      {stage1_46[148], stage1_46[149], stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153]},
      {stage2_48[24],stage2_47[28],stage2_46[34],stage2_45[66],stage2_44[99]}
   );
   gpc615_5 gpc6794 (
      {stage1_44[179], stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183]},
      {stage1_45[27]},
      {stage1_46[154], stage1_46[155], stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159]},
      {stage2_48[25],stage2_47[29],stage2_46[35],stage2_45[67],stage2_44[100]}
   );
   gpc615_5 gpc6795 (
      {stage1_44[184], stage1_44[185], stage1_44[186], stage1_44[187], stage1_44[188]},
      {stage1_45[28]},
      {stage1_46[160], stage1_46[161], stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165]},
      {stage2_48[26],stage2_47[30],stage2_46[36],stage2_45[68],stage2_44[101]}
   );
   gpc615_5 gpc6796 (
      {stage1_44[189], stage1_44[190], stage1_44[191], stage1_44[192], stage1_44[193]},
      {stage1_45[29]},
      {stage1_46[166], stage1_46[167], stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171]},
      {stage2_48[27],stage2_47[31],stage2_46[37],stage2_45[69],stage2_44[102]}
   );
   gpc615_5 gpc6797 (
      {stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197], stage1_44[198]},
      {stage1_45[30]},
      {stage1_46[172], stage1_46[173], stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177]},
      {stage2_48[28],stage2_47[32],stage2_46[38],stage2_45[70],stage2_44[103]}
   );
   gpc615_5 gpc6798 (
      {stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_45[31]},
      {stage1_46[178], stage1_46[179], stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183]},
      {stage2_48[29],stage2_47[33],stage2_46[39],stage2_45[71],stage2_44[104]}
   );
   gpc615_5 gpc6799 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208]},
      {stage1_45[32]},
      {stage1_46[184], stage1_46[185], stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189]},
      {stage2_48[30],stage2_47[34],stage2_46[40],stage2_45[72],stage2_44[105]}
   );
   gpc615_5 gpc6800 (
      {stage1_44[209], stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213]},
      {stage1_45[33]},
      {stage1_46[190], stage1_46[191], stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195]},
      {stage2_48[31],stage2_47[35],stage2_46[41],stage2_45[73],stage2_44[106]}
   );
   gpc615_5 gpc6801 (
      {stage1_44[214], stage1_44[215], stage1_44[216], stage1_44[217], stage1_44[218]},
      {stage1_45[34]},
      {stage1_46[196], stage1_46[197], stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201]},
      {stage2_48[32],stage2_47[36],stage2_46[42],stage2_45[74],stage2_44[107]}
   );
   gpc615_5 gpc6802 (
      {stage1_44[219], stage1_44[220], stage1_44[221], stage1_44[222], stage1_44[223]},
      {stage1_45[35]},
      {stage1_46[202], stage1_46[203], stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207]},
      {stage2_48[33],stage2_47[37],stage2_46[43],stage2_45[75],stage2_44[108]}
   );
   gpc615_5 gpc6803 (
      {stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227], stage1_44[228]},
      {stage1_45[36]},
      {stage1_46[208], stage1_46[209], stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213]},
      {stage2_48[34],stage2_47[38],stage2_46[44],stage2_45[76],stage2_44[109]}
   );
   gpc615_5 gpc6804 (
      {stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_45[37]},
      {stage1_46[214], stage1_46[215], stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219]},
      {stage2_48[35],stage2_47[39],stage2_46[45],stage2_45[77],stage2_44[110]}
   );
   gpc615_5 gpc6805 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238]},
      {stage1_45[38]},
      {stage1_46[220], stage1_46[221], stage1_46[222], stage1_46[223], stage1_46[224], stage1_46[225]},
      {stage2_48[36],stage2_47[40],stage2_46[46],stage2_45[78],stage2_44[111]}
   );
   gpc615_5 gpc6806 (
      {stage1_44[239], stage1_44[240], stage1_44[241], stage1_44[242], stage1_44[243]},
      {stage1_45[39]},
      {stage1_46[226], stage1_46[227], stage1_46[228], stage1_46[229], stage1_46[230], stage1_46[231]},
      {stage2_48[37],stage2_47[41],stage2_46[47],stage2_45[79],stage2_44[112]}
   );
   gpc606_5 gpc6807 (
      {stage1_45[40], stage1_45[41], stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[38],stage2_47[42],stage2_46[48],stage2_45[80]}
   );
   gpc606_5 gpc6808 (
      {stage1_45[46], stage1_45[47], stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[39],stage2_47[43],stage2_46[49],stage2_45[81]}
   );
   gpc606_5 gpc6809 (
      {stage1_45[52], stage1_45[53], stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[40],stage2_47[44],stage2_46[50],stage2_45[82]}
   );
   gpc606_5 gpc6810 (
      {stage1_45[58], stage1_45[59], stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[41],stage2_47[45],stage2_46[51],stage2_45[83]}
   );
   gpc606_5 gpc6811 (
      {stage1_45[64], stage1_45[65], stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[42],stage2_47[46],stage2_46[52],stage2_45[84]}
   );
   gpc606_5 gpc6812 (
      {stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[43],stage2_47[47],stage2_46[53],stage2_45[85]}
   );
   gpc606_5 gpc6813 (
      {stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[44],stage2_47[48],stage2_46[54],stage2_45[86]}
   );
   gpc606_5 gpc6814 (
      {stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[45],stage2_47[49],stage2_46[55],stage2_45[87]}
   );
   gpc606_5 gpc6815 (
      {stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[46],stage2_47[50],stage2_46[56],stage2_45[88]}
   );
   gpc606_5 gpc6816 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98], stage1_45[99]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[47],stage2_47[51],stage2_46[57],stage2_45[89]}
   );
   gpc606_5 gpc6817 (
      {stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103], stage1_45[104], stage1_45[105]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[48],stage2_47[52],stage2_46[58],stage2_45[90]}
   );
   gpc606_5 gpc6818 (
      {stage1_45[106], stage1_45[107], stage1_45[108], stage1_45[109], stage1_45[110], stage1_45[111]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[49],stage2_47[53],stage2_46[59],stage2_45[91]}
   );
   gpc606_5 gpc6819 (
      {stage1_45[112], stage1_45[113], stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[50],stage2_47[54],stage2_46[60],stage2_45[92]}
   );
   gpc606_5 gpc6820 (
      {stage1_45[118], stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[51],stage2_47[55],stage2_46[61],stage2_45[93]}
   );
   gpc606_5 gpc6821 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128], stage1_45[129]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[52],stage2_47[56],stage2_46[62],stage2_45[94]}
   );
   gpc606_5 gpc6822 (
      {stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133], stage1_45[134], stage1_45[135]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[53],stage2_47[57],stage2_46[63],stage2_45[95]}
   );
   gpc606_5 gpc6823 (
      {stage1_45[136], stage1_45[137], stage1_45[138], stage1_45[139], stage1_45[140], stage1_45[141]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[54],stage2_47[58],stage2_46[64],stage2_45[96]}
   );
   gpc615_5 gpc6824 (
      {stage1_45[142], stage1_45[143], stage1_45[144], stage1_45[145], stage1_45[146]},
      {stage1_46[232]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[55],stage2_47[59],stage2_46[65],stage2_45[97]}
   );
   gpc615_5 gpc6825 (
      {stage1_45[147], stage1_45[148], stage1_45[149], stage1_45[150], stage1_45[151]},
      {stage1_46[233]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[56],stage2_47[60],stage2_46[66],stage2_45[98]}
   );
   gpc615_5 gpc6826 (
      {stage1_45[152], stage1_45[153], stage1_45[154], stage1_45[155], stage1_45[156]},
      {stage1_46[234]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[57],stage2_47[61],stage2_46[67],stage2_45[99]}
   );
   gpc615_5 gpc6827 (
      {stage1_46[235], stage1_46[236], stage1_46[237], stage1_46[238], stage1_46[239]},
      {stage1_47[120]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[20],stage2_48[58],stage2_47[62],stage2_46[68]}
   );
   gpc615_5 gpc6828 (
      {stage1_46[240], stage1_46[241], stage1_46[242], stage1_46[243], stage1_46[244]},
      {stage1_47[121]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[21],stage2_48[59],stage2_47[63],stage2_46[69]}
   );
   gpc615_5 gpc6829 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[122]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[22],stage2_48[60],stage2_47[64],stage2_46[70]}
   );
   gpc615_5 gpc6830 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[123]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[23],stage2_48[61],stage2_47[65],stage2_46[71]}
   );
   gpc615_5 gpc6831 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[124]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[24],stage2_48[62],stage2_47[66],stage2_46[72]}
   );
   gpc615_5 gpc6832 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[125]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[25],stage2_48[63],stage2_47[67],stage2_46[73]}
   );
   gpc615_5 gpc6833 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[126]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[26],stage2_48[64],stage2_47[68],stage2_46[74]}
   );
   gpc615_5 gpc6834 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[127]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[27],stage2_48[65],stage2_47[69],stage2_46[75]}
   );
   gpc615_5 gpc6835 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[128]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[28],stage2_48[66],stage2_47[70],stage2_46[76]}
   );
   gpc615_5 gpc6836 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[129]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[29],stage2_48[67],stage2_47[71],stage2_46[77]}
   );
   gpc615_5 gpc6837 (
      {stage1_47[130], stage1_47[131], stage1_47[132], stage1_47[133], stage1_47[134]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[30],stage2_48[68],stage2_47[72]}
   );
   gpc615_5 gpc6838 (
      {stage1_47[135], stage1_47[136], stage1_47[137], stage1_47[138], stage1_47[139]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[31],stage2_48[69],stage2_47[73]}
   );
   gpc615_5 gpc6839 (
      {stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143], stage1_47[144]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[32],stage2_48[70],stage2_47[74]}
   );
   gpc615_5 gpc6840 (
      {stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[33],stage2_48[71],stage2_47[75]}
   );
   gpc615_5 gpc6841 (
      {stage1_47[150], stage1_47[151], stage1_47[152], stage1_47[153], stage1_47[154]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[34],stage2_48[72],stage2_47[76]}
   );
   gpc615_5 gpc6842 (
      {stage1_47[155], stage1_47[156], stage1_47[157], stage1_47[158], stage1_47[159]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[35],stage2_48[73],stage2_47[77]}
   );
   gpc615_5 gpc6843 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[36],stage2_48[74],stage2_47[78]}
   );
   gpc615_5 gpc6844 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[37],stage2_48[75],stage2_47[79]}
   );
   gpc615_5 gpc6845 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[38],stage2_48[76],stage2_47[80]}
   );
   gpc615_5 gpc6846 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[39],stage2_48[77],stage2_47[81]}
   );
   gpc615_5 gpc6847 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[40],stage2_48[78],stage2_47[82]}
   );
   gpc615_5 gpc6848 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[41],stage2_48[79],stage2_47[83]}
   );
   gpc615_5 gpc6849 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[42],stage2_48[80],stage2_47[84]}
   );
   gpc615_5 gpc6850 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[43],stage2_48[81],stage2_47[85]}
   );
   gpc615_5 gpc6851 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[74]},
      {stage1_49[84], stage1_49[85], stage1_49[86], stage1_49[87], stage1_49[88], stage1_49[89]},
      {stage2_51[14],stage2_50[24],stage2_49[44],stage2_48[82],stage2_47[86]}
   );
   gpc615_5 gpc6852 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[75]},
      {stage1_49[90], stage1_49[91], stage1_49[92], stage1_49[93], stage1_49[94], stage1_49[95]},
      {stage2_51[15],stage2_50[25],stage2_49[45],stage2_48[83],stage2_47[87]}
   );
   gpc615_5 gpc6853 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[76]},
      {stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99], stage1_49[100], stage1_49[101]},
      {stage2_51[16],stage2_50[26],stage2_49[46],stage2_48[84],stage2_47[88]}
   );
   gpc615_5 gpc6854 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[77]},
      {stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105], stage1_49[106], stage1_49[107]},
      {stage2_51[17],stage2_50[27],stage2_49[47],stage2_48[85],stage2_47[89]}
   );
   gpc615_5 gpc6855 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[78]},
      {stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111], stage1_49[112], stage1_49[113]},
      {stage2_51[18],stage2_50[28],stage2_49[48],stage2_48[86],stage2_47[90]}
   );
   gpc615_5 gpc6856 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[79]},
      {stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117], stage1_49[118], stage1_49[119]},
      {stage2_51[19],stage2_50[29],stage2_49[49],stage2_48[87],stage2_47[91]}
   );
   gpc615_5 gpc6857 (
      {stage1_47[230], stage1_47[231], stage1_47[232], stage1_47[233], stage1_47[234]},
      {stage1_48[80]},
      {stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123], stage1_49[124], stage1_49[125]},
      {stage2_51[20],stage2_50[30],stage2_49[50],stage2_48[88],stage2_47[92]}
   );
   gpc615_5 gpc6858 (
      {stage1_47[235], stage1_47[236], stage1_47[237], stage1_47[238], stage1_47[239]},
      {stage1_48[81]},
      {stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129], stage1_49[130], stage1_49[131]},
      {stage2_51[21],stage2_50[31],stage2_49[51],stage2_48[89],stage2_47[93]}
   );
   gpc615_5 gpc6859 (
      {stage1_47[240], stage1_47[241], stage1_47[242], stage1_47[243], stage1_47[244]},
      {stage1_48[82]},
      {stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135], stage1_49[136], stage1_49[137]},
      {stage2_51[22],stage2_50[32],stage2_49[52],stage2_48[90],stage2_47[94]}
   );
   gpc615_5 gpc6860 (
      {stage1_47[245], stage1_47[246], stage1_47[247], stage1_47[248], stage1_47[249]},
      {stage1_48[83]},
      {stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141], stage1_49[142], stage1_49[143]},
      {stage2_51[23],stage2_50[33],stage2_49[53],stage2_48[91],stage2_47[95]}
   );
   gpc615_5 gpc6861 (
      {stage1_47[250], stage1_47[251], stage1_47[252], stage1_47[253], stage1_47[254]},
      {stage1_48[84]},
      {stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147], stage1_49[148], stage1_49[149]},
      {stage2_51[24],stage2_50[34],stage2_49[54],stage2_48[92],stage2_47[96]}
   );
   gpc615_5 gpc6862 (
      {stage1_47[255], stage1_47[256], stage1_47[257], stage1_47[258], stage1_47[259]},
      {stage1_48[85]},
      {stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153], stage1_49[154], stage1_49[155]},
      {stage2_51[25],stage2_50[35],stage2_49[55],stage2_48[93],stage2_47[97]}
   );
   gpc615_5 gpc6863 (
      {stage1_47[260], stage1_47[261], stage1_47[262], stage1_47[263], stage1_47[264]},
      {stage1_48[86]},
      {stage1_49[156], stage1_49[157], stage1_49[158], stage1_49[159], stage1_49[160], stage1_49[161]},
      {stage2_51[26],stage2_50[36],stage2_49[56],stage2_48[94],stage2_47[98]}
   );
   gpc615_5 gpc6864 (
      {stage1_47[265], stage1_47[266], stage1_47[267], stage1_47[268], stage1_47[269]},
      {stage1_48[87]},
      {stage1_49[162], stage1_49[163], stage1_49[164], stage1_49[165], stage1_49[166], stage1_49[167]},
      {stage2_51[27],stage2_50[37],stage2_49[57],stage2_48[95],stage2_47[99]}
   );
   gpc606_5 gpc6865 (
      {stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91], stage1_48[92], stage1_48[93]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[28],stage2_50[38],stage2_49[58],stage2_48[96]}
   );
   gpc606_5 gpc6866 (
      {stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97], stage1_48[98], stage1_48[99]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[29],stage2_50[39],stage2_49[59],stage2_48[97]}
   );
   gpc606_5 gpc6867 (
      {stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103], stage1_48[104], stage1_48[105]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[30],stage2_50[40],stage2_49[60],stage2_48[98]}
   );
   gpc606_5 gpc6868 (
      {stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109], stage1_48[110], stage1_48[111]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[31],stage2_50[41],stage2_49[61],stage2_48[99]}
   );
   gpc606_5 gpc6869 (
      {stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115], stage1_48[116], stage1_48[117]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[32],stage2_50[42],stage2_49[62],stage2_48[100]}
   );
   gpc606_5 gpc6870 (
      {stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121], stage1_48[122], stage1_48[123]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[33],stage2_50[43],stage2_49[63],stage2_48[101]}
   );
   gpc606_5 gpc6871 (
      {stage1_48[124], stage1_48[125], stage1_48[126], stage1_48[127], stage1_48[128], stage1_48[129]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[34],stage2_50[44],stage2_49[64],stage2_48[102]}
   );
   gpc606_5 gpc6872 (
      {stage1_48[130], stage1_48[131], stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[35],stage2_50[45],stage2_49[65],stage2_48[103]}
   );
   gpc606_5 gpc6873 (
      {stage1_48[136], stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[36],stage2_50[46],stage2_49[66],stage2_48[104]}
   );
   gpc606_5 gpc6874 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146], stage1_48[147]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[37],stage2_50[47],stage2_49[67],stage2_48[105]}
   );
   gpc606_5 gpc6875 (
      {stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151], stage1_48[152], stage1_48[153]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[38],stage2_50[48],stage2_49[68],stage2_48[106]}
   );
   gpc606_5 gpc6876 (
      {stage1_48[154], stage1_48[155], stage1_48[156], stage1_48[157], stage1_48[158], stage1_48[159]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[39],stage2_50[49],stage2_49[69],stage2_48[107]}
   );
   gpc606_5 gpc6877 (
      {stage1_48[160], stage1_48[161], stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[40],stage2_50[50],stage2_49[70],stage2_48[108]}
   );
   gpc606_5 gpc6878 (
      {stage1_49[168], stage1_49[169], stage1_49[170], stage1_49[171], stage1_49[172], stage1_49[173]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[13],stage2_51[41],stage2_50[51],stage2_49[71]}
   );
   gpc606_5 gpc6879 (
      {stage1_49[174], stage1_49[175], stage1_49[176], stage1_49[177], stage1_49[178], stage1_49[179]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[14],stage2_51[42],stage2_50[52],stage2_49[72]}
   );
   gpc606_5 gpc6880 (
      {stage1_49[180], stage1_49[181], stage1_49[182], stage1_49[183], stage1_49[184], stage1_49[185]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[15],stage2_51[43],stage2_50[53],stage2_49[73]}
   );
   gpc606_5 gpc6881 (
      {stage1_49[186], stage1_49[187], stage1_49[188], stage1_49[189], stage1_49[190], stage1_49[191]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[16],stage2_51[44],stage2_50[54],stage2_49[74]}
   );
   gpc606_5 gpc6882 (
      {stage1_49[192], stage1_49[193], stage1_49[194], stage1_49[195], stage1_49[196], stage1_49[197]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[17],stage2_51[45],stage2_50[55],stage2_49[75]}
   );
   gpc615_5 gpc6883 (
      {stage1_49[198], stage1_49[199], stage1_49[200], stage1_49[201], stage1_49[202]},
      {stage1_50[78]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[18],stage2_51[46],stage2_50[56],stage2_49[76]}
   );
   gpc1163_5 gpc6884 (
      {stage1_50[79], stage1_50[80], stage1_50[81]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage1_52[0]},
      {stage1_53[0]},
      {stage2_54[0],stage2_53[6],stage2_52[19],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc6885 (
      {stage1_50[82], stage1_50[83], stage1_50[84]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage1_52[1]},
      {stage1_53[1]},
      {stage2_54[1],stage2_53[7],stage2_52[20],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc6886 (
      {stage1_50[85], stage1_50[86], stage1_50[87]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage1_52[2]},
      {stage1_53[2]},
      {stage2_54[2],stage2_53[8],stage2_52[21],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc6887 (
      {stage1_50[88], stage1_50[89], stage1_50[90]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage1_52[3]},
      {stage1_53[3]},
      {stage2_54[3],stage2_53[9],stage2_52[22],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc6888 (
      {stage1_50[91], stage1_50[92], stage1_50[93]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage1_52[4]},
      {stage1_53[4]},
      {stage2_54[4],stage2_53[10],stage2_52[23],stage2_51[51],stage2_50[61]}
   );
   gpc615_5 gpc6889 (
      {stage1_50[94], stage1_50[95], stage1_50[96], stage1_50[97], stage1_50[98]},
      {stage1_51[66]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[11],stage2_52[24],stage2_51[52],stage2_50[62]}
   );
   gpc615_5 gpc6890 (
      {stage1_50[99], stage1_50[100], stage1_50[101], stage1_50[102], stage1_50[103]},
      {stage1_51[67]},
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage2_54[6],stage2_53[12],stage2_52[25],stage2_51[53],stage2_50[63]}
   );
   gpc615_5 gpc6891 (
      {stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107], stage1_50[108]},
      {stage1_51[68]},
      {stage1_52[17], stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22]},
      {stage2_54[7],stage2_53[13],stage2_52[26],stage2_51[54],stage2_50[64]}
   );
   gpc615_5 gpc6892 (
      {stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112], stage1_50[113]},
      {stage1_51[69]},
      {stage1_52[23], stage1_52[24], stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28]},
      {stage2_54[8],stage2_53[14],stage2_52[27],stage2_51[55],stage2_50[65]}
   );
   gpc615_5 gpc6893 (
      {stage1_50[114], stage1_50[115], stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[70]},
      {stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34]},
      {stage2_54[9],stage2_53[15],stage2_52[28],stage2_51[56],stage2_50[66]}
   );
   gpc615_5 gpc6894 (
      {stage1_50[119], stage1_50[120], stage1_50[121], stage1_50[122], stage1_50[123]},
      {stage1_51[71]},
      {stage1_52[35], stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40]},
      {stage2_54[10],stage2_53[16],stage2_52[29],stage2_51[57],stage2_50[67]}
   );
   gpc615_5 gpc6895 (
      {stage1_50[124], stage1_50[125], stage1_50[126], stage1_50[127], stage1_50[128]},
      {stage1_51[72]},
      {stage1_52[41], stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46]},
      {stage2_54[11],stage2_53[17],stage2_52[30],stage2_51[58],stage2_50[68]}
   );
   gpc615_5 gpc6896 (
      {stage1_50[129], stage1_50[130], stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[73]},
      {stage1_52[47], stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52]},
      {stage2_54[12],stage2_53[18],stage2_52[31],stage2_51[59],stage2_50[69]}
   );
   gpc606_5 gpc6897 (
      {stage1_51[74], stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79]},
      {stage1_53[5], stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10]},
      {stage2_55[0],stage2_54[13],stage2_53[19],stage2_52[32],stage2_51[60]}
   );
   gpc606_5 gpc6898 (
      {stage1_51[80], stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85]},
      {stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16]},
      {stage2_55[1],stage2_54[14],stage2_53[20],stage2_52[33],stage2_51[61]}
   );
   gpc606_5 gpc6899 (
      {stage1_51[86], stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91]},
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22]},
      {stage2_55[2],stage2_54[15],stage2_53[21],stage2_52[34],stage2_51[62]}
   );
   gpc606_5 gpc6900 (
      {stage1_51[92], stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97]},
      {stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28]},
      {stage2_55[3],stage2_54[16],stage2_53[22],stage2_52[35],stage2_51[63]}
   );
   gpc606_5 gpc6901 (
      {stage1_51[98], stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103]},
      {stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage2_55[4],stage2_54[17],stage2_53[23],stage2_52[36],stage2_51[64]}
   );
   gpc606_5 gpc6902 (
      {stage1_51[104], stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109]},
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40]},
      {stage2_55[5],stage2_54[18],stage2_53[24],stage2_52[37],stage2_51[65]}
   );
   gpc606_5 gpc6903 (
      {stage1_51[110], stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115]},
      {stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46]},
      {stage2_55[6],stage2_54[19],stage2_53[25],stage2_52[38],stage2_51[66]}
   );
   gpc606_5 gpc6904 (
      {stage1_51[116], stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121]},
      {stage1_53[47], stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52]},
      {stage2_55[7],stage2_54[20],stage2_53[26],stage2_52[39],stage2_51[67]}
   );
   gpc606_5 gpc6905 (
      {stage1_51[122], stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127]},
      {stage1_53[53], stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58]},
      {stage2_55[8],stage2_54[21],stage2_53[27],stage2_52[40],stage2_51[68]}
   );
   gpc606_5 gpc6906 (
      {stage1_51[128], stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133]},
      {stage1_53[59], stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64]},
      {stage2_55[9],stage2_54[22],stage2_53[28],stage2_52[41],stage2_51[69]}
   );
   gpc606_5 gpc6907 (
      {stage1_51[134], stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139]},
      {stage1_53[65], stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70]},
      {stage2_55[10],stage2_54[23],stage2_53[29],stage2_52[42],stage2_51[70]}
   );
   gpc606_5 gpc6908 (
      {stage1_51[140], stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145]},
      {stage1_53[71], stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76]},
      {stage2_55[11],stage2_54[24],stage2_53[30],stage2_52[43],stage2_51[71]}
   );
   gpc606_5 gpc6909 (
      {stage1_51[146], stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151]},
      {stage1_53[77], stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82]},
      {stage2_55[12],stage2_54[25],stage2_53[31],stage2_52[44],stage2_51[72]}
   );
   gpc606_5 gpc6910 (
      {stage1_51[152], stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157]},
      {stage1_53[83], stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88]},
      {stage2_55[13],stage2_54[26],stage2_53[32],stage2_52[45],stage2_51[73]}
   );
   gpc606_5 gpc6911 (
      {stage1_51[158], stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163]},
      {stage1_53[89], stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94]},
      {stage2_55[14],stage2_54[27],stage2_53[33],stage2_52[46],stage2_51[74]}
   );
   gpc606_5 gpc6912 (
      {stage1_51[164], stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169]},
      {stage1_53[95], stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100]},
      {stage2_55[15],stage2_54[28],stage2_53[34],stage2_52[47],stage2_51[75]}
   );
   gpc606_5 gpc6913 (
      {stage1_51[170], stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175]},
      {stage1_53[101], stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106]},
      {stage2_55[16],stage2_54[29],stage2_53[35],stage2_52[48],stage2_51[76]}
   );
   gpc606_5 gpc6914 (
      {stage1_51[176], stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181]},
      {stage1_53[107], stage1_53[108], stage1_53[109], stage1_53[110], stage1_53[111], stage1_53[112]},
      {stage2_55[17],stage2_54[30],stage2_53[36],stage2_52[49],stage2_51[77]}
   );
   gpc606_5 gpc6915 (
      {stage1_51[182], stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187]},
      {stage1_53[113], stage1_53[114], stage1_53[115], stage1_53[116], stage1_53[117], stage1_53[118]},
      {stage2_55[18],stage2_54[31],stage2_53[37],stage2_52[50],stage2_51[78]}
   );
   gpc606_5 gpc6916 (
      {stage1_51[188], stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193]},
      {stage1_53[119], stage1_53[120], stage1_53[121], stage1_53[122], stage1_53[123], stage1_53[124]},
      {stage2_55[19],stage2_54[32],stage2_53[38],stage2_52[51],stage2_51[79]}
   );
   gpc606_5 gpc6917 (
      {stage1_51[194], stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199]},
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129], stage1_53[130]},
      {stage2_55[20],stage2_54[33],stage2_53[39],stage2_52[52],stage2_51[80]}
   );
   gpc606_5 gpc6918 (
      {stage1_51[200], stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_53[131], stage1_53[132], stage1_53[133], stage1_53[134], stage1_53[135], stage1_53[136]},
      {stage2_55[21],stage2_54[34],stage2_53[40],stage2_52[53],stage2_51[81]}
   );
   gpc606_5 gpc6919 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210], stage1_51[211]},
      {stage1_53[137], stage1_53[138], stage1_53[139], stage1_53[140], stage1_53[141], stage1_53[142]},
      {stage2_55[22],stage2_54[35],stage2_53[41],stage2_52[54],stage2_51[82]}
   );
   gpc606_5 gpc6920 (
      {stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215], stage1_51[216], stage1_51[217]},
      {stage1_53[143], stage1_53[144], stage1_53[145], stage1_53[146], stage1_53[147], stage1_53[148]},
      {stage2_55[23],stage2_54[36],stage2_53[42],stage2_52[55],stage2_51[83]}
   );
   gpc606_5 gpc6921 (
      {stage1_51[218], stage1_51[219], stage1_51[220], stage1_51[221], stage1_51[222], stage1_51[223]},
      {stage1_53[149], stage1_53[150], stage1_53[151], stage1_53[152], stage1_53[153], stage1_53[154]},
      {stage2_55[24],stage2_54[37],stage2_53[43],stage2_52[56],stage2_51[84]}
   );
   gpc606_5 gpc6922 (
      {stage1_52[53], stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[25],stage2_54[38],stage2_53[44],stage2_52[57]}
   );
   gpc606_5 gpc6923 (
      {stage1_52[59], stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[26],stage2_54[39],stage2_53[45],stage2_52[58]}
   );
   gpc606_5 gpc6924 (
      {stage1_52[65], stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[27],stage2_54[40],stage2_53[46],stage2_52[59]}
   );
   gpc606_5 gpc6925 (
      {stage1_52[71], stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[28],stage2_54[41],stage2_53[47],stage2_52[60]}
   );
   gpc606_5 gpc6926 (
      {stage1_52[77], stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[29],stage2_54[42],stage2_53[48],stage2_52[61]}
   );
   gpc606_5 gpc6927 (
      {stage1_52[83], stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[30],stage2_54[43],stage2_53[49],stage2_52[62]}
   );
   gpc606_5 gpc6928 (
      {stage1_52[89], stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[31],stage2_54[44],stage2_53[50],stage2_52[63]}
   );
   gpc606_5 gpc6929 (
      {stage1_52[95], stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[32],stage2_54[45],stage2_53[51],stage2_52[64]}
   );
   gpc606_5 gpc6930 (
      {stage1_52[101], stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[33],stage2_54[46],stage2_53[52],stage2_52[65]}
   );
   gpc606_5 gpc6931 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111], stage1_52[112]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[34],stage2_54[47],stage2_53[53],stage2_52[66]}
   );
   gpc606_5 gpc6932 (
      {stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116], stage1_52[117], stage1_52[118]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[35],stage2_54[48],stage2_53[54],stage2_52[67]}
   );
   gpc606_5 gpc6933 (
      {stage1_52[119], stage1_52[120], stage1_52[121], stage1_52[122], stage1_52[123], stage1_52[124]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[36],stage2_54[49],stage2_53[55],stage2_52[68]}
   );
   gpc606_5 gpc6934 (
      {stage1_52[125], stage1_52[126], stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[37],stage2_54[50],stage2_53[56],stage2_52[69]}
   );
   gpc606_5 gpc6935 (
      {stage1_52[131], stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[38],stage2_54[51],stage2_53[57],stage2_52[70]}
   );
   gpc606_5 gpc6936 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141], stage1_52[142]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[39],stage2_54[52],stage2_53[58],stage2_52[71]}
   );
   gpc606_5 gpc6937 (
      {stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146], stage1_52[147], stage1_52[148]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[40],stage2_54[53],stage2_53[59],stage2_52[72]}
   );
   gpc606_5 gpc6938 (
      {stage1_52[149], stage1_52[150], stage1_52[151], stage1_52[152], stage1_52[153], stage1_52[154]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[41],stage2_54[54],stage2_53[60],stage2_52[73]}
   );
   gpc606_5 gpc6939 (
      {stage1_52[155], stage1_52[156], stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[42],stage2_54[55],stage2_53[61],stage2_52[74]}
   );
   gpc606_5 gpc6940 (
      {stage1_52[161], stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[43],stage2_54[56],stage2_53[62],stage2_52[75]}
   );
   gpc606_5 gpc6941 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171], stage1_52[172]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[44],stage2_54[57],stage2_53[63],stage2_52[76]}
   );
   gpc606_5 gpc6942 (
      {stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176], stage1_52[177], stage1_52[178]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[45],stage2_54[58],stage2_53[64],stage2_52[77]}
   );
   gpc606_5 gpc6943 (
      {stage1_52[179], stage1_52[180], stage1_52[181], stage1_52[182], stage1_52[183], stage1_52[184]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[46],stage2_54[59],stage2_53[65],stage2_52[78]}
   );
   gpc606_5 gpc6944 (
      {stage1_52[185], stage1_52[186], stage1_52[187], stage1_52[188], stage1_52[189], stage1_52[190]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[47],stage2_54[60],stage2_53[66],stage2_52[79]}
   );
   gpc606_5 gpc6945 (
      {stage1_52[191], stage1_52[192], stage1_52[193], stage1_52[194], stage1_52[195], stage1_52[196]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[48],stage2_54[61],stage2_53[67],stage2_52[80]}
   );
   gpc606_5 gpc6946 (
      {stage1_52[197], stage1_52[198], stage1_52[199], stage1_52[200], stage1_52[201], stage1_52[202]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[49],stage2_54[62],stage2_53[68],stage2_52[81]}
   );
   gpc606_5 gpc6947 (
      {stage1_52[203], stage1_52[204], stage1_52[205], stage1_52[206], stage1_52[207], stage1_52[208]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[50],stage2_54[63],stage2_53[69],stage2_52[82]}
   );
   gpc606_5 gpc6948 (
      {stage1_52[209], stage1_52[210], stage1_52[211], stage1_52[212], stage1_52[213], stage1_52[214]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[51],stage2_54[64],stage2_53[70],stage2_52[83]}
   );
   gpc606_5 gpc6949 (
      {stage1_52[215], stage1_52[216], stage1_52[217], stage1_52[218], stage1_52[219], stage1_52[220]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[52],stage2_54[65],stage2_53[71],stage2_52[84]}
   );
   gpc606_5 gpc6950 (
      {stage1_52[221], stage1_52[222], stage1_52[223], stage1_52[224], stage1_52[225], stage1_52[226]},
      {stage1_54[168], stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173]},
      {stage2_56[28],stage2_55[53],stage2_54[66],stage2_53[72],stage2_52[85]}
   );
   gpc606_5 gpc6951 (
      {stage1_52[227], stage1_52[228], stage1_52[229], stage1_52[230], stage1_52[231], stage1_52[232]},
      {stage1_54[174], stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179]},
      {stage2_56[29],stage2_55[54],stage2_54[67],stage2_53[73],stage2_52[86]}
   );
   gpc606_5 gpc6952 (
      {stage1_52[233], stage1_52[234], stage1_52[235], stage1_52[236], stage1_52[237], stage1_52[238]},
      {stage1_54[180], stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185]},
      {stage2_56[30],stage2_55[55],stage2_54[68],stage2_53[74],stage2_52[87]}
   );
   gpc606_5 gpc6953 (
      {stage1_52[239], stage1_52[240], stage1_52[241], stage1_52[242], stage1_52[243], stage1_52[244]},
      {stage1_54[186], stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191]},
      {stage2_56[31],stage2_55[56],stage2_54[69],stage2_53[75],stage2_52[88]}
   );
   gpc606_5 gpc6954 (
      {stage1_52[245], stage1_52[246], stage1_52[247], stage1_52[248], stage1_52[249], stage1_52[250]},
      {stage1_54[192], stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage2_56[32],stage2_55[57],stage2_54[70],stage2_53[76],stage2_52[89]}
   );
   gpc606_5 gpc6955 (
      {stage1_52[251], stage1_52[252], stage1_52[253], stage1_52[254], stage1_52[255], stage1_52[256]},
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202], stage1_54[203]},
      {stage2_56[33],stage2_55[58],stage2_54[71],stage2_53[77],stage2_52[90]}
   );
   gpc606_5 gpc6956 (
      {stage1_52[257], stage1_52[258], stage1_52[259], stage1_52[260], stage1_52[261], stage1_52[262]},
      {stage1_54[204], stage1_54[205], stage1_54[206], stage1_54[207], stage1_54[208], stage1_54[209]},
      {stage2_56[34],stage2_55[59],stage2_54[72],stage2_53[78],stage2_52[91]}
   );
   gpc606_5 gpc6957 (
      {stage1_52[263], stage1_52[264], stage1_52[265], stage1_52[266], stage1_52[267], stage1_52[268]},
      {stage1_54[210], stage1_54[211], stage1_54[212], stage1_54[213], stage1_54[214], stage1_54[215]},
      {stage2_56[35],stage2_55[60],stage2_54[73],stage2_53[79],stage2_52[92]}
   );
   gpc606_5 gpc6958 (
      {stage1_53[155], stage1_53[156], stage1_53[157], stage1_53[158], stage1_53[159], stage1_53[160]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[36],stage2_55[61],stage2_54[74],stage2_53[80]}
   );
   gpc606_5 gpc6959 (
      {stage1_53[161], stage1_53[162], stage1_53[163], stage1_53[164], stage1_53[165], stage1_53[166]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[37],stage2_55[62],stage2_54[75],stage2_53[81]}
   );
   gpc606_5 gpc6960 (
      {stage1_53[167], stage1_53[168], stage1_53[169], stage1_53[170], stage1_53[171], stage1_53[172]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[38],stage2_55[63],stage2_54[76],stage2_53[82]}
   );
   gpc2135_5 gpc6961 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[0], stage1_56[1], stage1_56[2]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[0],stage2_57[3],stage2_56[39],stage2_55[64]}
   );
   gpc2135_5 gpc6962 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[1],stage2_57[4],stage2_56[40],stage2_55[65]}
   );
   gpc2135_5 gpc6963 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[6], stage1_56[7], stage1_56[8]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[2],stage2_57[5],stage2_56[41],stage2_55[66]}
   );
   gpc2135_5 gpc6964 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[3],stage2_57[6],stage2_56[42],stage2_55[67]}
   );
   gpc2135_5 gpc6965 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12], stage1_56[13], stage1_56[14]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[4],stage2_57[7],stage2_56[43],stage2_55[68]}
   );
   gpc2135_5 gpc6966 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[5],stage2_57[8],stage2_56[44],stage2_55[69]}
   );
   gpc2135_5 gpc6967 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[18], stage1_56[19], stage1_56[20]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[6],stage2_57[9],stage2_56[45],stage2_55[70]}
   );
   gpc2135_5 gpc6968 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[7],stage2_57[10],stage2_56[46],stage2_55[71]}
   );
   gpc2135_5 gpc6969 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[24], stage1_56[25], stage1_56[26]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[8],stage2_57[11],stage2_56[47],stage2_55[72]}
   );
   gpc2135_5 gpc6970 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[9],stage2_57[12],stage2_56[48],stage2_55[73]}
   );
   gpc2135_5 gpc6971 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[30], stage1_56[31], stage1_56[32]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[10],stage2_57[13],stage2_56[49],stage2_55[74]}
   );
   gpc2135_5 gpc6972 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[11],stage2_57[14],stage2_56[50],stage2_55[75]}
   );
   gpc2135_5 gpc6973 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[12],stage2_57[15],stage2_56[51],stage2_55[76]}
   );
   gpc2135_5 gpc6974 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[13],stage2_57[16],stage2_56[52],stage2_55[77]}
   );
   gpc2135_5 gpc6975 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[14],stage2_57[17],stage2_56[53],stage2_55[78]}
   );
   gpc2135_5 gpc6976 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[15],stage2_57[18],stage2_56[54],stage2_55[79]}
   );
   gpc2135_5 gpc6977 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[16],stage2_57[19],stage2_56[55],stage2_55[80]}
   );
   gpc2135_5 gpc6978 (
      {stage1_55[103], stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[17],stage2_57[20],stage2_56[56],stage2_55[81]}
   );
   gpc2135_5 gpc6979 (
      {stage1_55[108], stage1_55[109], stage1_55[110], stage1_55[111], stage1_55[112]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[18]},
      {stage1_58[36], stage1_58[37]},
      {stage2_59[18],stage2_58[18],stage2_57[21],stage2_56[57],stage2_55[82]}
   );
   gpc2135_5 gpc6980 (
      {stage1_55[113], stage1_55[114], stage1_55[115], stage1_55[116], stage1_55[117]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[19]},
      {stage1_58[38], stage1_58[39]},
      {stage2_59[19],stage2_58[19],stage2_57[22],stage2_56[58],stage2_55[83]}
   );
   gpc2135_5 gpc6981 (
      {stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121], stage1_55[122]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[20]},
      {stage1_58[40], stage1_58[41]},
      {stage2_59[20],stage2_58[20],stage2_57[23],stage2_56[59],stage2_55[84]}
   );
   gpc2135_5 gpc6982 (
      {stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[21]},
      {stage1_58[42], stage1_58[43]},
      {stage2_59[21],stage2_58[21],stage2_57[24],stage2_56[60],stage2_55[85]}
   );
   gpc2135_5 gpc6983 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[22]},
      {stage1_58[44], stage1_58[45]},
      {stage2_59[22],stage2_58[22],stage2_57[25],stage2_56[61],stage2_55[86]}
   );
   gpc2135_5 gpc6984 (
      {stage1_55[133], stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[23]},
      {stage1_58[46], stage1_58[47]},
      {stage2_59[23],stage2_58[23],stage2_57[26],stage2_56[62],stage2_55[87]}
   );
   gpc2135_5 gpc6985 (
      {stage1_55[138], stage1_55[139], stage1_55[140], stage1_55[141], stage1_55[142]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[24]},
      {stage1_58[48], stage1_58[49]},
      {stage2_59[24],stage2_58[24],stage2_57[27],stage2_56[63],stage2_55[88]}
   );
   gpc2135_5 gpc6986 (
      {stage1_55[143], stage1_55[144], stage1_55[145], stage1_55[146], stage1_55[147]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[25]},
      {stage1_58[50], stage1_58[51]},
      {stage2_59[25],stage2_58[25],stage2_57[28],stage2_56[64],stage2_55[89]}
   );
   gpc2135_5 gpc6987 (
      {stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151], stage1_55[152]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[26]},
      {stage1_58[52], stage1_58[53]},
      {stage2_59[26],stage2_58[26],stage2_57[29],stage2_56[65],stage2_55[90]}
   );
   gpc2135_5 gpc6988 (
      {stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[27]},
      {stage1_58[54], stage1_58[55]},
      {stage2_59[27],stage2_58[27],stage2_57[30],stage2_56[66],stage2_55[91]}
   );
   gpc2135_5 gpc6989 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[28]},
      {stage1_58[56], stage1_58[57]},
      {stage2_59[28],stage2_58[28],stage2_57[31],stage2_56[67],stage2_55[92]}
   );
   gpc2135_5 gpc6990 (
      {stage1_55[163], stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[29]},
      {stage1_58[58], stage1_58[59]},
      {stage2_59[29],stage2_58[29],stage2_57[32],stage2_56[68],stage2_55[93]}
   );
   gpc606_5 gpc6991 (
      {stage1_55[168], stage1_55[169], stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[30],stage2_58[30],stage2_57[33],stage2_56[69],stage2_55[94]}
   );
   gpc615_5 gpc6992 (
      {stage1_55[174], stage1_55[175], stage1_55[176], stage1_55[177], stage1_55[178]},
      {stage1_56[90]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[31],stage2_58[31],stage2_57[34],stage2_56[70],stage2_55[95]}
   );
   gpc615_5 gpc6993 (
      {stage1_55[179], stage1_55[180], stage1_55[181], stage1_55[182], stage1_55[183]},
      {stage1_56[91]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[32],stage2_58[32],stage2_57[35],stage2_56[71],stage2_55[96]}
   );
   gpc615_5 gpc6994 (
      {stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187], stage1_55[188]},
      {stage1_56[92]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[33],stage2_58[33],stage2_57[36],stage2_56[72],stage2_55[97]}
   );
   gpc615_5 gpc6995 (
      {stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_56[93]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[34],stage2_58[34],stage2_57[37],stage2_56[73],stage2_55[98]}
   );
   gpc615_5 gpc6996 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198]},
      {stage1_56[94]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[35],stage2_58[35],stage2_57[38],stage2_56[74],stage2_55[99]}
   );
   gpc615_5 gpc6997 (
      {stage1_55[199], stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203]},
      {stage1_56[95]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[36],stage2_58[36],stage2_57[39],stage2_56[75],stage2_55[100]}
   );
   gpc615_5 gpc6998 (
      {stage1_55[204], stage1_55[205], stage1_55[206], stage1_55[207], stage1_55[208]},
      {stage1_56[96]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[37],stage2_58[37],stage2_57[40],stage2_56[76],stage2_55[101]}
   );
   gpc615_5 gpc6999 (
      {stage1_55[209], stage1_55[210], stage1_55[211], stage1_55[212], stage1_55[213]},
      {stage1_56[97]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[38],stage2_58[38],stage2_57[41],stage2_56[77],stage2_55[102]}
   );
   gpc615_5 gpc7000 (
      {stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217], stage1_55[218]},
      {stage1_56[98]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[39],stage2_58[39],stage2_57[42],stage2_56[78],stage2_55[103]}
   );
   gpc606_5 gpc7001 (
      {stage1_56[99], stage1_56[100], stage1_56[101], stage1_56[102], stage1_56[103], stage1_56[104]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[0],stage2_59[40],stage2_58[40],stage2_57[43],stage2_56[79]}
   );
   gpc606_5 gpc7002 (
      {stage1_56[105], stage1_56[106], stage1_56[107], stage1_56[108], stage1_56[109], stage1_56[110]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[1],stage2_59[41],stage2_58[41],stage2_57[44],stage2_56[80]}
   );
   gpc606_5 gpc7003 (
      {stage1_56[111], stage1_56[112], stage1_56[113], stage1_56[114], stage1_56[115], stage1_56[116]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[2],stage2_59[42],stage2_58[42],stage2_57[45],stage2_56[81]}
   );
   gpc606_5 gpc7004 (
      {stage1_56[117], stage1_56[118], stage1_56[119], stage1_56[120], stage1_56[121], stage1_56[122]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[3],stage2_59[43],stage2_58[43],stage2_57[46],stage2_56[82]}
   );
   gpc606_5 gpc7005 (
      {stage1_56[123], stage1_56[124], stage1_56[125], stage1_56[126], stage1_56[127], stage1_56[128]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[4],stage2_59[44],stage2_58[44],stage2_57[47],stage2_56[83]}
   );
   gpc606_5 gpc7006 (
      {stage1_56[129], stage1_56[130], stage1_56[131], stage1_56[132], stage1_56[133], stage1_56[134]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[5],stage2_59[45],stage2_58[45],stage2_57[48],stage2_56[84]}
   );
   gpc606_5 gpc7007 (
      {stage1_56[135], stage1_56[136], stage1_56[137], stage1_56[138], stage1_56[139], stage1_56[140]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[6],stage2_59[46],stage2_58[46],stage2_57[49],stage2_56[85]}
   );
   gpc606_5 gpc7008 (
      {stage1_56[141], stage1_56[142], stage1_56[143], stage1_56[144], stage1_56[145], stage1_56[146]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[7],stage2_59[47],stage2_58[47],stage2_57[50],stage2_56[86]}
   );
   gpc606_5 gpc7009 (
      {stage1_56[147], stage1_56[148], stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[8],stage2_59[48],stage2_58[48],stage2_57[51],stage2_56[87]}
   );
   gpc606_5 gpc7010 (
      {stage1_56[153], stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_58[114], stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage2_60[9],stage2_59[49],stage2_58[49],stage2_57[52],stage2_56[88]}
   );
   gpc606_5 gpc7011 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163], stage1_56[164]},
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124], stage1_58[125]},
      {stage2_60[10],stage2_59[50],stage2_58[50],stage2_57[53],stage2_56[89]}
   );
   gpc606_5 gpc7012 (
      {stage1_56[165], stage1_56[166], stage1_56[167], stage1_56[168], stage1_56[169], stage1_56[170]},
      {stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129], stage1_58[130], stage1_58[131]},
      {stage2_60[11],stage2_59[51],stage2_58[51],stage2_57[54],stage2_56[90]}
   );
   gpc606_5 gpc7013 (
      {stage1_56[171], stage1_56[172], stage1_56[173], stage1_56[174], stage1_56[175], stage1_56[176]},
      {stage1_58[132], stage1_58[133], stage1_58[134], stage1_58[135], stage1_58[136], stage1_58[137]},
      {stage2_60[12],stage2_59[52],stage2_58[52],stage2_57[55],stage2_56[91]}
   );
   gpc606_5 gpc7014 (
      {stage1_56[177], stage1_56[178], stage1_56[179], stage1_56[180], stage1_56[181], stage1_56[182]},
      {stage1_58[138], stage1_58[139], stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143]},
      {stage2_60[13],stage2_59[53],stage2_58[53],stage2_57[56],stage2_56[92]}
   );
   gpc606_5 gpc7015 (
      {stage1_56[183], stage1_56[184], stage1_56[185], stage1_56[186], stage1_56[187], stage1_56[188]},
      {stage1_58[144], stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage2_60[14],stage2_59[54],stage2_58[54],stage2_57[57],stage2_56[93]}
   );
   gpc606_5 gpc7016 (
      {stage1_56[189], stage1_56[190], stage1_56[191], stage1_56[192], stage1_56[193], stage1_56[194]},
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154], stage1_58[155]},
      {stage2_60[15],stage2_59[55],stage2_58[55],stage2_57[58],stage2_56[94]}
   );
   gpc606_5 gpc7017 (
      {stage1_56[195], stage1_56[196], stage1_56[197], stage1_56[198], stage1_56[199], stage1_56[200]},
      {stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159], stage1_58[160], stage1_58[161]},
      {stage2_60[16],stage2_59[56],stage2_58[56],stage2_57[59],stage2_56[95]}
   );
   gpc606_5 gpc7018 (
      {stage1_56[201], stage1_56[202], stage1_56[203], stage1_56[204], stage1_56[205], stage1_56[206]},
      {stage1_58[162], stage1_58[163], stage1_58[164], stage1_58[165], stage1_58[166], stage1_58[167]},
      {stage2_60[17],stage2_59[57],stage2_58[57],stage2_57[60],stage2_56[96]}
   );
   gpc606_5 gpc7019 (
      {stage1_56[207], stage1_56[208], stage1_56[209], stage1_56[210], stage1_56[211], stage1_56[212]},
      {stage1_58[168], stage1_58[169], stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173]},
      {stage2_60[18],stage2_59[58],stage2_58[58],stage2_57[61],stage2_56[97]}
   );
   gpc606_5 gpc7020 (
      {stage1_56[213], stage1_56[214], stage1_56[215], stage1_56[216], stage1_56[217], stage1_56[218]},
      {stage1_58[174], stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage2_60[19],stage2_59[59],stage2_58[59],stage2_57[62],stage2_56[98]}
   );
   gpc606_5 gpc7021 (
      {stage1_56[219], stage1_56[220], stage1_56[221], stage1_56[222], stage1_56[223], stage1_56[224]},
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184], stage1_58[185]},
      {stage2_60[20],stage2_59[60],stage2_58[60],stage2_57[63],stage2_56[99]}
   );
   gpc606_5 gpc7022 (
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[21],stage2_59[61],stage2_58[61],stage2_57[64]}
   );
   gpc606_5 gpc7023 (
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[22],stage2_59[62],stage2_58[62],stage2_57[65]}
   );
   gpc606_5 gpc7024 (
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[23],stage2_59[63],stage2_58[63],stage2_57[66]}
   );
   gpc606_5 gpc7025 (
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[24],stage2_59[64],stage2_58[64],stage2_57[67]}
   );
   gpc606_5 gpc7026 (
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage2_61[4],stage2_60[25],stage2_59[65],stage2_58[65],stage2_57[68]}
   );
   gpc606_5 gpc7027 (
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage2_61[5],stage2_60[26],stage2_59[66],stage2_58[66],stage2_57[69]}
   );
   gpc606_5 gpc7028 (
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage2_61[6],stage2_60[27],stage2_59[67],stage2_58[67],stage2_57[70]}
   );
   gpc606_5 gpc7029 (
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage1_59[42], stage1_59[43], stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47]},
      {stage2_61[7],stage2_60[28],stage2_59[68],stage2_58[68],stage2_57[71]}
   );
   gpc606_5 gpc7030 (
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage1_59[48], stage1_59[49], stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53]},
      {stage2_61[8],stage2_60[29],stage2_59[69],stage2_58[69],stage2_57[72]}
   );
   gpc606_5 gpc7031 (
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage1_59[54], stage1_59[55], stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59]},
      {stage2_61[9],stage2_60[30],stage2_59[70],stage2_58[70],stage2_57[73]}
   );
   gpc606_5 gpc7032 (
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage1_59[60], stage1_59[61], stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65]},
      {stage2_61[10],stage2_60[31],stage2_59[71],stage2_58[71],stage2_57[74]}
   );
   gpc606_5 gpc7033 (
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage1_59[66], stage1_59[67], stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71]},
      {stage2_61[11],stage2_60[32],stage2_59[72],stage2_58[72],stage2_57[75]}
   );
   gpc606_5 gpc7034 (
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage1_59[72], stage1_59[73], stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77]},
      {stage2_61[12],stage2_60[33],stage2_59[73],stage2_58[73],stage2_57[76]}
   );
   gpc606_5 gpc7035 (
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage1_59[78], stage1_59[79], stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83]},
      {stage2_61[13],stage2_60[34],stage2_59[74],stage2_58[74],stage2_57[77]}
   );
   gpc606_5 gpc7036 (
      {stage1_57[174], stage1_57[175], stage1_57[176], stage1_57[177], stage1_57[178], stage1_57[179]},
      {stage1_59[84], stage1_59[85], stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89]},
      {stage2_61[14],stage2_60[35],stage2_59[75],stage2_58[75],stage2_57[78]}
   );
   gpc117_4 gpc7037 (
      {stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189], stage1_58[190], stage1_58[191], stage1_58[192]},
      {stage1_59[90]},
      {stage1_60[0]},
      {stage2_61[15],stage2_60[36],stage2_59[76],stage2_58[76]}
   );
   gpc117_4 gpc7038 (
      {stage1_58[193], stage1_58[194], stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[91]},
      {stage1_60[1]},
      {stage2_61[16],stage2_60[37],stage2_59[77],stage2_58[77]}
   );
   gpc117_4 gpc7039 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204], stage1_58[205], stage1_58[206]},
      {stage1_59[92]},
      {stage1_60[2]},
      {stage2_61[17],stage2_60[38],stage2_59[78],stage2_58[78]}
   );
   gpc117_4 gpc7040 (
      {stage1_58[207], stage1_58[208], stage1_58[209], stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213]},
      {stage1_59[93]},
      {stage1_60[3]},
      {stage2_61[18],stage2_60[39],stage2_59[79],stage2_58[79]}
   );
   gpc606_5 gpc7041 (
      {stage1_58[214], stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_60[4], stage1_60[5], stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9]},
      {stage2_62[0],stage2_61[19],stage2_60[40],stage2_59[80],stage2_58[80]}
   );
   gpc606_5 gpc7042 (
      {stage1_58[220], stage1_58[221], stage1_58[222], stage1_58[223], stage1_58[224], stage1_58[225]},
      {stage1_60[10], stage1_60[11], stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15]},
      {stage2_62[1],stage2_61[20],stage2_60[41],stage2_59[81],stage2_58[81]}
   );
   gpc606_5 gpc7043 (
      {stage1_58[226], stage1_58[227], stage1_58[228], stage1_58[229], stage1_58[230], stage1_58[231]},
      {stage1_60[16], stage1_60[17], stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21]},
      {stage2_62[2],stage2_61[21],stage2_60[42],stage2_59[82],stage2_58[82]}
   );
   gpc606_5 gpc7044 (
      {stage1_58[232], stage1_58[233], stage1_58[234], stage1_58[235], stage1_58[236], stage1_58[237]},
      {stage1_60[22], stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage2_62[3],stage2_61[22],stage2_60[43],stage2_59[83],stage2_58[83]}
   );
   gpc606_5 gpc7045 (
      {stage1_58[238], stage1_58[239], stage1_58[240], stage1_58[241], stage1_58[242], 1'b0},
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33]},
      {stage2_62[4],stage2_61[23],stage2_60[44],stage2_59[84],stage2_58[84]}
   );
   gpc606_5 gpc7046 (
      {stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97], stage1_59[98], stage1_59[99]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[24],stage2_60[45],stage2_59[85]}
   );
   gpc606_5 gpc7047 (
      {stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103], stage1_59[104], stage1_59[105]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[25],stage2_60[46],stage2_59[86]}
   );
   gpc606_5 gpc7048 (
      {stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109], stage1_59[110], stage1_59[111]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[26],stage2_60[47],stage2_59[87]}
   );
   gpc606_5 gpc7049 (
      {stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115], stage1_59[116], stage1_59[117]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[27],stage2_60[48],stage2_59[88]}
   );
   gpc606_5 gpc7050 (
      {stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121], stage1_59[122], stage1_59[123]},
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage2_63[4],stage2_62[9],stage2_61[28],stage2_60[49],stage2_59[89]}
   );
   gpc606_5 gpc7051 (
      {stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127], stage1_59[128], stage1_59[129]},
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage2_63[5],stage2_62[10],stage2_61[29],stage2_60[50],stage2_59[90]}
   );
   gpc606_5 gpc7052 (
      {stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133], stage1_59[134], stage1_59[135]},
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage2_63[6],stage2_62[11],stage2_61[30],stage2_60[51],stage2_59[91]}
   );
   gpc606_5 gpc7053 (
      {stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139], stage1_59[140], stage1_59[141]},
      {stage1_61[42], stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage2_63[7],stage2_62[12],stage2_61[31],stage2_60[52],stage2_59[92]}
   );
   gpc606_5 gpc7054 (
      {stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145], stage1_59[146], stage1_59[147]},
      {stage1_61[48], stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53]},
      {stage2_63[8],stage2_62[13],stage2_61[32],stage2_60[53],stage2_59[93]}
   );
   gpc606_5 gpc7055 (
      {stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151], stage1_59[152], stage1_59[153]},
      {stage1_61[54], stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59]},
      {stage2_63[9],stage2_62[14],stage2_61[33],stage2_60[54],stage2_59[94]}
   );
   gpc606_5 gpc7056 (
      {stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157], stage1_59[158], stage1_59[159]},
      {stage1_61[60], stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65]},
      {stage2_63[10],stage2_62[15],stage2_61[34],stage2_60[55],stage2_59[95]}
   );
   gpc606_5 gpc7057 (
      {stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163], stage1_59[164], stage1_59[165]},
      {stage1_61[66], stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71]},
      {stage2_63[11],stage2_62[16],stage2_61[35],stage2_60[56],stage2_59[96]}
   );
   gpc606_5 gpc7058 (
      {stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169], stage1_59[170], stage1_59[171]},
      {stage1_61[72], stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77]},
      {stage2_63[12],stage2_62[17],stage2_61[36],stage2_60[57],stage2_59[97]}
   );
   gpc606_5 gpc7059 (
      {stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175], stage1_59[176], stage1_59[177]},
      {stage1_61[78], stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83]},
      {stage2_63[13],stage2_62[18],stage2_61[37],stage2_60[58],stage2_59[98]}
   );
   gpc606_5 gpc7060 (
      {stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181], stage1_59[182], stage1_59[183]},
      {stage1_61[84], stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89]},
      {stage2_63[14],stage2_62[19],stage2_61[38],stage2_60[59],stage2_59[99]}
   );
   gpc606_5 gpc7061 (
      {stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187], stage1_59[188], stage1_59[189]},
      {stage1_61[90], stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95]},
      {stage2_63[15],stage2_62[20],stage2_61[39],stage2_60[60],stage2_59[100]}
   );
   gpc606_5 gpc7062 (
      {stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193], stage1_59[194], stage1_59[195]},
      {stage1_61[96], stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101]},
      {stage2_63[16],stage2_62[21],stage2_61[40],stage2_60[61],stage2_59[101]}
   );
   gpc606_5 gpc7063 (
      {stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199], stage1_59[200], stage1_59[201]},
      {stage1_61[102], stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107]},
      {stage2_63[17],stage2_62[22],stage2_61[41],stage2_60[62],stage2_59[102]}
   );
   gpc606_5 gpc7064 (
      {stage1_59[202], stage1_59[203], stage1_59[204], stage1_59[205], stage1_59[206], stage1_59[207]},
      {stage1_61[108], stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113]},
      {stage2_63[18],stage2_62[23],stage2_61[42],stage2_60[63],stage2_59[103]}
   );
   gpc606_5 gpc7065 (
      {stage1_59[208], stage1_59[209], stage1_59[210], stage1_59[211], stage1_59[212], stage1_59[213]},
      {stage1_61[114], stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119]},
      {stage2_63[19],stage2_62[24],stage2_61[43],stage2_60[64],stage2_59[104]}
   );
   gpc606_5 gpc7066 (
      {stage1_59[214], stage1_59[215], stage1_59[216], stage1_59[217], stage1_59[218], stage1_59[219]},
      {stage1_61[120], stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125]},
      {stage2_63[20],stage2_62[25],stage2_61[44],stage2_60[65],stage2_59[105]}
   );
   gpc606_5 gpc7067 (
      {stage1_59[220], stage1_59[221], stage1_59[222], stage1_59[223], stage1_59[224], stage1_59[225]},
      {stage1_61[126], stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131]},
      {stage2_63[21],stage2_62[26],stage2_61[45],stage2_60[66],stage2_59[106]}
   );
   gpc606_5 gpc7068 (
      {stage1_59[226], stage1_59[227], stage1_59[228], stage1_59[229], stage1_59[230], stage1_59[231]},
      {stage1_61[132], stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137]},
      {stage2_63[22],stage2_62[27],stage2_61[46],stage2_60[67],stage2_59[107]}
   );
   gpc606_5 gpc7069 (
      {stage1_59[232], stage1_59[233], stage1_59[234], stage1_59[235], stage1_59[236], stage1_59[237]},
      {stage1_61[138], stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143]},
      {stage2_63[23],stage2_62[28],stage2_61[47],stage2_60[68],stage2_59[108]}
   );
   gpc606_5 gpc7070 (
      {stage1_59[238], stage1_59[239], stage1_59[240], stage1_59[241], stage1_59[242], stage1_59[243]},
      {stage1_61[144], stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149]},
      {stage2_63[24],stage2_62[29],stage2_61[48],stage2_60[69],stage2_59[109]}
   );
   gpc606_5 gpc7071 (
      {stage1_59[244], stage1_59[245], stage1_59[246], stage1_59[247], stage1_59[248], stage1_59[249]},
      {stage1_61[150], stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155]},
      {stage2_63[25],stage2_62[30],stage2_61[49],stage2_60[70],stage2_59[110]}
   );
   gpc606_5 gpc7072 (
      {stage1_59[250], stage1_59[251], stage1_59[252], stage1_59[253], stage1_59[254], stage1_59[255]},
      {stage1_61[156], stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161]},
      {stage2_63[26],stage2_62[31],stage2_61[50],stage2_60[71],stage2_59[111]}
   );
   gpc606_5 gpc7073 (
      {stage1_59[256], stage1_59[257], stage1_59[258], stage1_59[259], stage1_59[260], stage1_59[261]},
      {stage1_61[162], stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167]},
      {stage2_63[27],stage2_62[32],stage2_61[51],stage2_60[72],stage2_59[112]}
   );
   gpc606_5 gpc7074 (
      {stage1_59[262], stage1_59[263], stage1_59[264], stage1_59[265], stage1_59[266], stage1_59[267]},
      {stage1_61[168], stage1_61[169], stage1_61[170], stage1_61[171], stage1_61[172], stage1_61[173]},
      {stage2_63[28],stage2_62[33],stage2_61[52],stage2_60[73],stage2_59[113]}
   );
   gpc1406_5 gpc7075 (
      {stage1_60[34], stage1_60[35], stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3]},
      {stage1_63[0]},
      {stage2_64[0],stage2_63[29],stage2_62[34],stage2_61[53],stage2_60[74]}
   );
   gpc606_5 gpc7076 (
      {stage1_60[40], stage1_60[41], stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45]},
      {stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9]},
      {stage2_64[1],stage2_63[30],stage2_62[35],stage2_61[54],stage2_60[75]}
   );
   gpc606_5 gpc7077 (
      {stage1_60[46], stage1_60[47], stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51]},
      {stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15]},
      {stage2_64[2],stage2_63[31],stage2_62[36],stage2_61[55],stage2_60[76]}
   );
   gpc606_5 gpc7078 (
      {stage1_60[52], stage1_60[53], stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57]},
      {stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21]},
      {stage2_64[3],stage2_63[32],stage2_62[37],stage2_61[56],stage2_60[77]}
   );
   gpc606_5 gpc7079 (
      {stage1_60[58], stage1_60[59], stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63]},
      {stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27]},
      {stage2_64[4],stage2_63[33],stage2_62[38],stage2_61[57],stage2_60[78]}
   );
   gpc606_5 gpc7080 (
      {stage1_60[64], stage1_60[65], stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69]},
      {stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33]},
      {stage2_64[5],stage2_63[34],stage2_62[39],stage2_61[58],stage2_60[79]}
   );
   gpc606_5 gpc7081 (
      {stage1_60[70], stage1_60[71], stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75]},
      {stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39]},
      {stage2_64[6],stage2_63[35],stage2_62[40],stage2_61[59],stage2_60[80]}
   );
   gpc606_5 gpc7082 (
      {stage1_60[76], stage1_60[77], stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81]},
      {stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage2_64[7],stage2_63[36],stage2_62[41],stage2_61[60],stage2_60[81]}
   );
   gpc606_5 gpc7083 (
      {stage1_60[82], stage1_60[83], stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87]},
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51]},
      {stage2_64[8],stage2_63[37],stage2_62[42],stage2_61[61],stage2_60[82]}
   );
   gpc606_5 gpc7084 (
      {stage1_60[88], stage1_60[89], stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93]},
      {stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57]},
      {stage2_64[9],stage2_63[38],stage2_62[43],stage2_61[62],stage2_60[83]}
   );
   gpc606_5 gpc7085 (
      {stage1_60[94], stage1_60[95], stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99]},
      {stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63]},
      {stage2_64[10],stage2_63[39],stage2_62[44],stage2_61[63],stage2_60[84]}
   );
   gpc606_5 gpc7086 (
      {stage1_60[100], stage1_60[101], stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105]},
      {stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69]},
      {stage2_64[11],stage2_63[40],stage2_62[45],stage2_61[64],stage2_60[85]}
   );
   gpc606_5 gpc7087 (
      {stage1_60[106], stage1_60[107], stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111]},
      {stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75]},
      {stage2_64[12],stage2_63[41],stage2_62[46],stage2_61[65],stage2_60[86]}
   );
   gpc606_5 gpc7088 (
      {stage1_60[112], stage1_60[113], stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117]},
      {stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79], stage1_62[80], stage1_62[81]},
      {stage2_64[13],stage2_63[42],stage2_62[47],stage2_61[66],stage2_60[87]}
   );
   gpc606_5 gpc7089 (
      {stage1_60[118], stage1_60[119], stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123]},
      {stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85], stage1_62[86], stage1_62[87]},
      {stage2_64[14],stage2_63[43],stage2_62[48],stage2_61[67],stage2_60[88]}
   );
   gpc606_5 gpc7090 (
      {stage1_60[124], stage1_60[125], stage1_60[126], stage1_60[127], stage1_60[128], stage1_60[129]},
      {stage1_62[88], stage1_62[89], stage1_62[90], stage1_62[91], stage1_62[92], stage1_62[93]},
      {stage2_64[15],stage2_63[44],stage2_62[49],stage2_61[68],stage2_60[89]}
   );
   gpc606_5 gpc7091 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[94], stage1_62[95], stage1_62[96], stage1_62[97], stage1_62[98], stage1_62[99]},
      {stage2_64[16],stage2_63[45],stage2_62[50],stage2_61[69],stage2_60[90]}
   );
   gpc606_5 gpc7092 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[100], stage1_62[101], stage1_62[102], stage1_62[103], stage1_62[104], stage1_62[105]},
      {stage2_64[17],stage2_63[46],stage2_62[51],stage2_61[70],stage2_60[91]}
   );
   gpc606_5 gpc7093 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[106], stage1_62[107], stage1_62[108], stage1_62[109], stage1_62[110], stage1_62[111]},
      {stage2_64[18],stage2_63[47],stage2_62[52],stage2_61[71],stage2_60[92]}
   );
   gpc606_5 gpc7094 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[112], stage1_62[113], stage1_62[114], stage1_62[115], stage1_62[116], stage1_62[117]},
      {stage2_64[19],stage2_63[48],stage2_62[53],stage2_61[72],stage2_60[93]}
   );
   gpc606_5 gpc7095 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[118], stage1_62[119], stage1_62[120], stage1_62[121], stage1_62[122], stage1_62[123]},
      {stage2_64[20],stage2_63[49],stage2_62[54],stage2_61[73],stage2_60[94]}
   );
   gpc615_5 gpc7096 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164]},
      {stage1_61[174]},
      {stage1_62[124], stage1_62[125], stage1_62[126], stage1_62[127], stage1_62[128], stage1_62[129]},
      {stage2_64[21],stage2_63[50],stage2_62[55],stage2_61[74],stage2_60[95]}
   );
   gpc615_5 gpc7097 (
      {stage1_60[165], stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169]},
      {stage1_61[175]},
      {stage1_62[130], stage1_62[131], stage1_62[132], stage1_62[133], stage1_62[134], stage1_62[135]},
      {stage2_64[22],stage2_63[51],stage2_62[56],stage2_61[75],stage2_60[96]}
   );
   gpc615_5 gpc7098 (
      {stage1_60[170], stage1_60[171], stage1_60[172], stage1_60[173], stage1_60[174]},
      {stage1_61[176]},
      {stage1_62[136], stage1_62[137], stage1_62[138], stage1_62[139], stage1_62[140], stage1_62[141]},
      {stage2_64[23],stage2_63[52],stage2_62[57],stage2_61[76],stage2_60[97]}
   );
   gpc615_5 gpc7099 (
      {stage1_60[175], stage1_60[176], stage1_60[177], stage1_60[178], stage1_60[179]},
      {stage1_61[177]},
      {stage1_62[142], stage1_62[143], stage1_62[144], stage1_62[145], stage1_62[146], stage1_62[147]},
      {stage2_64[24],stage2_63[53],stage2_62[58],stage2_61[77],stage2_60[98]}
   );
   gpc615_5 gpc7100 (
      {stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183], stage1_60[184]},
      {stage1_61[178]},
      {stage1_62[148], stage1_62[149], stage1_62[150], stage1_62[151], stage1_62[152], stage1_62[153]},
      {stage2_64[25],stage2_63[54],stage2_62[59],stage2_61[78],stage2_60[99]}
   );
   gpc615_5 gpc7101 (
      {stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188], stage1_60[189]},
      {stage1_61[179]},
      {stage1_62[154], stage1_62[155], stage1_62[156], stage1_62[157], stage1_62[158], stage1_62[159]},
      {stage2_64[26],stage2_63[55],stage2_62[60],stage2_61[79],stage2_60[100]}
   );
   gpc606_5 gpc7102 (
      {stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183], stage1_61[184], stage1_61[185]},
      {stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6]},
      {stage2_65[0],stage2_64[27],stage2_63[56],stage2_62[61],stage2_61[80]}
   );
   gpc606_5 gpc7103 (
      {stage1_61[186], stage1_61[187], stage1_61[188], stage1_61[189], stage1_61[190], stage1_61[191]},
      {stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12]},
      {stage2_65[1],stage2_64[28],stage2_63[57],stage2_62[62],stage2_61[81]}
   );
   gpc606_5 gpc7104 (
      {stage1_61[192], stage1_61[193], stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197]},
      {stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18]},
      {stage2_65[2],stage2_64[29],stage2_63[58],stage2_62[63],stage2_61[82]}
   );
   gpc1163_5 gpc7105 (
      {stage1_62[160], stage1_62[161], stage1_62[162]},
      {stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[3],stage2_64[30],stage2_63[59],stage2_62[64]}
   );
   gpc1163_5 gpc7106 (
      {stage1_62[163], stage1_62[164], stage1_62[165]},
      {stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29], stage1_63[30]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[4],stage2_64[31],stage2_63[60],stage2_62[65]}
   );
   gpc1163_5 gpc7107 (
      {stage1_62[166], stage1_62[167], stage1_62[168]},
      {stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35], stage1_63[36]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[5],stage2_64[32],stage2_63[61],stage2_62[66]}
   );
   gpc1163_5 gpc7108 (
      {stage1_62[169], stage1_62[170], stage1_62[171]},
      {stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41], stage1_63[42]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[6],stage2_64[33],stage2_63[62],stage2_62[67]}
   );
   gpc1163_5 gpc7109 (
      {stage1_62[172], stage1_62[173], stage1_62[174]},
      {stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47], stage1_63[48]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[7],stage2_64[34],stage2_63[63],stage2_62[68]}
   );
   gpc1163_5 gpc7110 (
      {stage1_62[175], stage1_62[176], stage1_62[177]},
      {stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53], stage1_63[54]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[8],stage2_64[35],stage2_63[64],stage2_62[69]}
   );
   gpc1163_5 gpc7111 (
      {stage1_62[178], stage1_62[179], stage1_62[180]},
      {stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59], stage1_63[60]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[9],stage2_64[36],stage2_63[65],stage2_62[70]}
   );
   gpc1163_5 gpc7112 (
      {stage1_62[181], stage1_62[182], stage1_62[183]},
      {stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65], stage1_63[66]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[10],stage2_64[37],stage2_63[66],stage2_62[71]}
   );
   gpc1163_5 gpc7113 (
      {stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71], stage1_63[72]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[11],stage2_64[38],stage2_63[67],stage2_62[72]}
   );
   gpc1163_5 gpc7114 (
      {stage1_62[187], stage1_62[188], stage1_62[189]},
      {stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77], stage1_63[78]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[12],stage2_64[39],stage2_63[68],stage2_62[73]}
   );
   gpc1163_5 gpc7115 (
      {stage1_62[190], stage1_62[191], stage1_62[192]},
      {stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83], stage1_63[84]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[13],stage2_64[40],stage2_63[69],stage2_62[74]}
   );
   gpc1163_5 gpc7116 (
      {stage1_62[193], stage1_62[194], stage1_62[195]},
      {stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89], stage1_63[90]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[14],stage2_64[41],stage2_63[70],stage2_62[75]}
   );
   gpc1163_5 gpc7117 (
      {stage1_62[196], stage1_62[197], stage1_62[198]},
      {stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95], stage1_63[96]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[15],stage2_64[42],stage2_63[71],stage2_62[76]}
   );
   gpc1163_5 gpc7118 (
      {stage1_62[199], stage1_62[200], stage1_62[201]},
      {stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101], stage1_63[102]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[16],stage2_64[43],stage2_63[72],stage2_62[77]}
   );
   gpc1163_5 gpc7119 (
      {stage1_62[202], stage1_62[203], stage1_62[204]},
      {stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107], stage1_63[108]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[17],stage2_64[44],stage2_63[73],stage2_62[78]}
   );
   gpc1163_5 gpc7120 (
      {stage1_62[205], stage1_62[206], stage1_62[207]},
      {stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113], stage1_63[114]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[18],stage2_64[45],stage2_63[74],stage2_62[79]}
   );
   gpc1163_5 gpc7121 (
      {stage1_62[208], stage1_62[209], stage1_62[210]},
      {stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119], stage1_63[120]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[19],stage2_64[46],stage2_63[75],stage2_62[80]}
   );
   gpc1163_5 gpc7122 (
      {stage1_62[211], stage1_62[212], stage1_62[213]},
      {stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125], stage1_63[126]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[20],stage2_64[47],stage2_63[76],stage2_62[81]}
   );
   gpc1163_5 gpc7123 (
      {stage1_62[214], stage1_62[215], stage1_62[216]},
      {stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131], stage1_63[132]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[21],stage2_64[48],stage2_63[77],stage2_62[82]}
   );
   gpc1163_5 gpc7124 (
      {stage1_62[217], stage1_62[218], stage1_62[219]},
      {stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137], stage1_63[138]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[22],stage2_64[49],stage2_63[78],stage2_62[83]}
   );
   gpc1163_5 gpc7125 (
      {stage1_62[220], stage1_62[221], stage1_62[222]},
      {stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143], stage1_63[144]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[23],stage2_64[50],stage2_63[79],stage2_62[84]}
   );
   gpc1163_5 gpc7126 (
      {stage1_62[223], stage1_62[224], stage1_62[225]},
      {stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149], stage1_63[150]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[24],stage2_64[51],stage2_63[80],stage2_62[85]}
   );
   gpc1163_5 gpc7127 (
      {stage1_62[226], stage1_62[227], stage1_62[228]},
      {stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155], stage1_63[156]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[25],stage2_64[52],stage2_63[81],stage2_62[86]}
   );
   gpc1163_5 gpc7128 (
      {stage1_62[229], stage1_62[230], stage1_62[231]},
      {stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161], stage1_63[162]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[26],stage2_64[53],stage2_63[82],stage2_62[87]}
   );
   gpc1163_5 gpc7129 (
      {stage1_62[232], stage1_62[233], stage1_62[234]},
      {stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167], stage1_63[168]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[27],stage2_64[54],stage2_63[83],stage2_62[88]}
   );
   gpc1163_5 gpc7130 (
      {stage1_62[235], stage1_62[236], stage1_62[237]},
      {stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173], stage1_63[174]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[28],stage2_64[55],stage2_63[84],stage2_62[89]}
   );
   gpc1163_5 gpc7131 (
      {stage1_62[238], stage1_62[239], stage1_62[240]},
      {stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179], stage1_63[180]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[29],stage2_64[56],stage2_63[85],stage2_62[90]}
   );
   gpc1163_5 gpc7132 (
      {stage1_62[241], stage1_62[242], stage1_62[243]},
      {stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185], stage1_63[186]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[30],stage2_64[57],stage2_63[86],stage2_62[91]}
   );
   gpc1163_5 gpc7133 (
      {stage1_62[244], stage1_62[245], stage1_62[246]},
      {stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191], stage1_63[192]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[31],stage2_64[58],stage2_63[87],stage2_62[92]}
   );
   gpc1163_5 gpc7134 (
      {stage1_62[247], stage1_62[248], stage1_62[249]},
      {stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197], stage1_63[198]},
      {stage1_64[29]},
      {stage1_65[29]},
      {stage2_66[29],stage2_65[32],stage2_64[59],stage2_63[88],stage2_62[93]}
   );
   gpc1163_5 gpc7135 (
      {stage1_62[250], stage1_62[251], stage1_62[252]},
      {stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203], stage1_63[204]},
      {stage1_64[30]},
      {stage1_65[30]},
      {stage2_66[30],stage2_65[33],stage2_64[60],stage2_63[89],stage2_62[94]}
   );
   gpc1163_5 gpc7136 (
      {stage1_62[253], stage1_62[254], stage1_62[255]},
      {stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209], stage1_63[210]},
      {stage1_64[31]},
      {stage1_65[31]},
      {stage2_66[31],stage2_65[34],stage2_64[61],stage2_63[90],stage2_62[95]}
   );
   gpc1163_5 gpc7137 (
      {stage1_62[256], stage1_62[257], stage1_62[258]},
      {stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215], stage1_63[216]},
      {stage1_64[32]},
      {stage1_65[32]},
      {stage2_66[32],stage2_65[35],stage2_64[62],stage2_63[91],stage2_62[96]}
   );
   gpc1163_5 gpc7138 (
      {stage1_62[259], stage1_62[260], stage1_62[261]},
      {stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221], stage1_63[222]},
      {stage1_64[33]},
      {stage1_65[33]},
      {stage2_66[33],stage2_65[36],stage2_64[63],stage2_63[92],stage2_62[97]}
   );
   gpc1163_5 gpc7139 (
      {stage1_62[262], stage1_62[263], stage1_62[264]},
      {stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227], stage1_63[228]},
      {stage1_64[34]},
      {stage1_65[34]},
      {stage2_66[34],stage2_65[37],stage2_64[64],stage2_63[93],stage2_62[98]}
   );
   gpc1163_5 gpc7140 (
      {stage1_62[265], stage1_62[266], stage1_62[267]},
      {stage1_63[229], stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[35]},
      {stage1_65[35]},
      {stage2_66[35],stage2_65[38],stage2_64[65],stage2_63[94],stage2_62[99]}
   );
   gpc1163_5 gpc7141 (
      {stage1_62[268], stage1_62[269], stage1_62[270]},
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239], stage1_63[240]},
      {stage1_64[36]},
      {stage1_65[36]},
      {stage2_66[36],stage2_65[39],stage2_64[66],stage2_63[95],stage2_62[100]}
   );
   gpc1163_5 gpc7142 (
      {stage1_62[271], stage1_62[272], stage1_62[273]},
      {stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_64[37]},
      {stage1_65[37]},
      {stage2_66[37],stage2_65[40],stage2_64[67],stage2_63[96],stage2_62[101]}
   );
   gpc1163_5 gpc7143 (
      {stage1_62[274], stage1_62[275], stage1_62[276]},
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252]},
      {stage1_64[38]},
      {stage1_65[38]},
      {stage2_66[38],stage2_65[41],stage2_64[68],stage2_63[97],stage2_62[102]}
   );
   gpc1163_5 gpc7144 (
      {stage1_62[277], stage1_62[278], stage1_62[279]},
      {stage1_63[253], stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258]},
      {stage1_64[39]},
      {stage1_65[39]},
      {stage2_66[39],stage2_65[42],stage2_64[69],stage2_63[98],stage2_62[103]}
   );
   gpc1163_5 gpc7145 (
      {stage1_62[280], stage1_62[281], stage1_62[282]},
      {stage1_63[259], stage1_63[260], stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264]},
      {stage1_64[40]},
      {stage1_65[40]},
      {stage2_66[40],stage2_65[43],stage2_64[70],stage2_63[99],stage2_62[104]}
   );
   gpc1163_5 gpc7146 (
      {stage1_62[283], stage1_62[284], stage1_62[285]},
      {stage1_63[265], stage1_63[266], stage1_63[267], stage1_63[268], stage1_63[269], stage1_63[270]},
      {stage1_64[41]},
      {stage1_65[41]},
      {stage2_66[41],stage2_65[44],stage2_64[71],stage2_63[100],stage2_62[105]}
   );
   gpc1163_5 gpc7147 (
      {stage1_62[286], stage1_62[287], stage1_62[288]},
      {stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274], stage1_63[275], stage1_63[276]},
      {stage1_64[42]},
      {stage1_65[42]},
      {stage2_66[42],stage2_65[45],stage2_64[72],stage2_63[101],stage2_62[106]}
   );
   gpc1163_5 gpc7148 (
      {stage1_62[289], stage1_62[290], stage1_62[291]},
      {stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281], stage1_63[282]},
      {stage1_64[43]},
      {stage1_65[43]},
      {stage2_66[43],stage2_65[46],stage2_64[73],stage2_63[102],stage2_62[107]}
   );
   gpc1163_5 gpc7149 (
      {stage1_62[292], stage1_62[293], stage1_62[294]},
      {stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_64[44]},
      {stage1_65[44]},
      {stage2_66[44],stage2_65[47],stage2_64[74],stage2_63[103],stage2_62[108]}
   );
   gpc1163_5 gpc7150 (
      {stage1_62[295], stage1_62[296], stage1_62[297]},
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294]},
      {stage1_64[45]},
      {stage1_65[45]},
      {stage2_66[45],stage2_65[48],stage2_64[75],stage2_63[104],stage2_62[109]}
   );
   gpc606_5 gpc7151 (
      {stage1_62[298], stage1_62[299], stage1_62[300], stage1_62[301], stage1_62[302], stage1_62[303]},
      {stage1_64[46], stage1_64[47], stage1_64[48], stage1_64[49], stage1_64[50], stage1_64[51]},
      {stage2_66[46],stage2_65[49],stage2_64[76],stage2_63[105],stage2_62[110]}
   );
   gpc606_5 gpc7152 (
      {stage1_62[304], stage1_62[305], stage1_62[306], stage1_62[307], stage1_62[308], stage1_62[309]},
      {stage1_64[52], stage1_64[53], stage1_64[54], stage1_64[55], stage1_64[56], stage1_64[57]},
      {stage2_66[47],stage2_65[50],stage2_64[77],stage2_63[106],stage2_62[111]}
   );
   gpc606_5 gpc7153 (
      {stage1_62[310], stage1_62[311], stage1_62[312], stage1_62[313], stage1_62[314], stage1_62[315]},
      {stage1_64[58], stage1_64[59], stage1_64[60], stage1_64[61], stage1_64[62], stage1_64[63]},
      {stage2_66[48],stage2_65[51],stage2_64[78],stage2_63[107],stage2_62[112]}
   );
   gpc606_5 gpc7154 (
      {stage1_62[316], stage1_62[317], stage1_62[318], stage1_62[319], stage1_62[320], stage1_62[321]},
      {stage1_64[64], stage1_64[65], stage1_64[66], stage1_64[67], stage1_64[68], stage1_64[69]},
      {stage2_66[49],stage2_65[52],stage2_64[79],stage2_63[108],stage2_62[113]}
   );
   gpc606_5 gpc7155 (
      {stage1_62[322], stage1_62[323], stage1_62[324], stage1_62[325], stage1_62[326], stage1_62[327]},
      {stage1_64[70], stage1_64[71], stage1_64[72], stage1_64[73], stage1_64[74], stage1_64[75]},
      {stage2_66[50],stage2_65[53],stage2_64[80],stage2_63[109],stage2_62[114]}
   );
   gpc606_5 gpc7156 (
      {stage1_62[328], stage1_62[329], stage1_62[330], stage1_62[331], stage1_62[332], stage1_62[333]},
      {stage1_64[76], stage1_64[77], stage1_64[78], stage1_64[79], stage1_64[80], stage1_64[81]},
      {stage2_66[51],stage2_65[54],stage2_64[81],stage2_63[110],stage2_62[115]}
   );
   gpc606_5 gpc7157 (
      {stage1_62[334], stage1_62[335], stage1_62[336], stage1_62[337], stage1_62[338], stage1_62[339]},
      {stage1_64[82], stage1_64[83], stage1_64[84], stage1_64[85], stage1_64[86], stage1_64[87]},
      {stage2_66[52],stage2_65[55],stage2_64[82],stage2_63[111],stage2_62[116]}
   );
   gpc606_5 gpc7158 (
      {stage1_62[340], stage1_62[341], stage1_62[342], stage1_62[343], stage1_62[344], stage1_62[345]},
      {stage1_64[88], stage1_64[89], stage1_64[90], stage1_64[91], stage1_64[92], stage1_64[93]},
      {stage2_66[53],stage2_65[56],stage2_64[83],stage2_63[112],stage2_62[117]}
   );
   gpc1_1 gpc7159 (
      {stage1_0[112]},
      {stage2_0[27]}
   );
   gpc1_1 gpc7160 (
      {stage1_0[113]},
      {stage2_0[28]}
   );
   gpc1_1 gpc7161 (
      {stage1_0[114]},
      {stage2_0[29]}
   );
   gpc1_1 gpc7162 (
      {stage1_0[115]},
      {stage2_0[30]}
   );
   gpc1_1 gpc7163 (
      {stage1_0[116]},
      {stage2_0[31]}
   );
   gpc1_1 gpc7164 (
      {stage1_0[117]},
      {stage2_0[32]}
   );
   gpc1_1 gpc7165 (
      {stage1_0[118]},
      {stage2_0[33]}
   );
   gpc1_1 gpc7166 (
      {stage1_2[208]},
      {stage2_2[60]}
   );
   gpc1_1 gpc7167 (
      {stage1_2[209]},
      {stage2_2[61]}
   );
   gpc1_1 gpc7168 (
      {stage1_2[210]},
      {stage2_2[62]}
   );
   gpc1_1 gpc7169 (
      {stage1_2[211]},
      {stage2_2[63]}
   );
   gpc1_1 gpc7170 (
      {stage1_2[212]},
      {stage2_2[64]}
   );
   gpc1_1 gpc7171 (
      {stage1_2[213]},
      {stage2_2[65]}
   );
   gpc1_1 gpc7172 (
      {stage1_2[214]},
      {stage2_2[66]}
   );
   gpc1_1 gpc7173 (
      {stage1_2[215]},
      {stage2_2[67]}
   );
   gpc1_1 gpc7174 (
      {stage1_2[216]},
      {stage2_2[68]}
   );
   gpc1_1 gpc7175 (
      {stage1_2[217]},
      {stage2_2[69]}
   );
   gpc1_1 gpc7176 (
      {stage1_2[218]},
      {stage2_2[70]}
   );
   gpc1_1 gpc7177 (
      {stage1_2[219]},
      {stage2_2[71]}
   );
   gpc1_1 gpc7178 (
      {stage1_2[220]},
      {stage2_2[72]}
   );
   gpc1_1 gpc7179 (
      {stage1_3[139]},
      {stage2_3[71]}
   );
   gpc1_1 gpc7180 (
      {stage1_3[140]},
      {stage2_3[72]}
   );
   gpc1_1 gpc7181 (
      {stage1_3[141]},
      {stage2_3[73]}
   );
   gpc1_1 gpc7182 (
      {stage1_3[142]},
      {stage2_3[74]}
   );
   gpc1_1 gpc7183 (
      {stage1_3[143]},
      {stage2_3[75]}
   );
   gpc1_1 gpc7184 (
      {stage1_3[144]},
      {stage2_3[76]}
   );
   gpc1_1 gpc7185 (
      {stage1_3[145]},
      {stage2_3[77]}
   );
   gpc1_1 gpc7186 (
      {stage1_3[146]},
      {stage2_3[78]}
   );
   gpc1_1 gpc7187 (
      {stage1_3[147]},
      {stage2_3[79]}
   );
   gpc1_1 gpc7188 (
      {stage1_3[148]},
      {stage2_3[80]}
   );
   gpc1_1 gpc7189 (
      {stage1_3[149]},
      {stage2_3[81]}
   );
   gpc1_1 gpc7190 (
      {stage1_3[150]},
      {stage2_3[82]}
   );
   gpc1_1 gpc7191 (
      {stage1_3[151]},
      {stage2_3[83]}
   );
   gpc1_1 gpc7192 (
      {stage1_3[152]},
      {stage2_3[84]}
   );
   gpc1_1 gpc7193 (
      {stage1_3[153]},
      {stage2_3[85]}
   );
   gpc1_1 gpc7194 (
      {stage1_3[154]},
      {stage2_3[86]}
   );
   gpc1_1 gpc7195 (
      {stage1_3[155]},
      {stage2_3[87]}
   );
   gpc1_1 gpc7196 (
      {stage1_3[156]},
      {stage2_3[88]}
   );
   gpc1_1 gpc7197 (
      {stage1_3[157]},
      {stage2_3[89]}
   );
   gpc1_1 gpc7198 (
      {stage1_3[158]},
      {stage2_3[90]}
   );
   gpc1_1 gpc7199 (
      {stage1_3[159]},
      {stage2_3[91]}
   );
   gpc1_1 gpc7200 (
      {stage1_3[160]},
      {stage2_3[92]}
   );
   gpc1_1 gpc7201 (
      {stage1_3[161]},
      {stage2_3[93]}
   );
   gpc1_1 gpc7202 (
      {stage1_3[162]},
      {stage2_3[94]}
   );
   gpc1_1 gpc7203 (
      {stage1_3[163]},
      {stage2_3[95]}
   );
   gpc1_1 gpc7204 (
      {stage1_3[164]},
      {stage2_3[96]}
   );
   gpc1_1 gpc7205 (
      {stage1_3[165]},
      {stage2_3[97]}
   );
   gpc1_1 gpc7206 (
      {stage1_3[166]},
      {stage2_3[98]}
   );
   gpc1_1 gpc7207 (
      {stage1_3[167]},
      {stage2_3[99]}
   );
   gpc1_1 gpc7208 (
      {stage1_3[168]},
      {stage2_3[100]}
   );
   gpc1_1 gpc7209 (
      {stage1_3[169]},
      {stage2_3[101]}
   );
   gpc1_1 gpc7210 (
      {stage1_3[170]},
      {stage2_3[102]}
   );
   gpc1_1 gpc7211 (
      {stage1_3[171]},
      {stage2_3[103]}
   );
   gpc1_1 gpc7212 (
      {stage1_3[172]},
      {stage2_3[104]}
   );
   gpc1_1 gpc7213 (
      {stage1_3[173]},
      {stage2_3[105]}
   );
   gpc1_1 gpc7214 (
      {stage1_3[174]},
      {stage2_3[106]}
   );
   gpc1_1 gpc7215 (
      {stage1_3[175]},
      {stage2_3[107]}
   );
   gpc1_1 gpc7216 (
      {stage1_3[176]},
      {stage2_3[108]}
   );
   gpc1_1 gpc7217 (
      {stage1_3[177]},
      {stage2_3[109]}
   );
   gpc1_1 gpc7218 (
      {stage1_3[178]},
      {stage2_3[110]}
   );
   gpc1_1 gpc7219 (
      {stage1_3[179]},
      {stage2_3[111]}
   );
   gpc1_1 gpc7220 (
      {stage1_3[180]},
      {stage2_3[112]}
   );
   gpc1_1 gpc7221 (
      {stage1_3[181]},
      {stage2_3[113]}
   );
   gpc1_1 gpc7222 (
      {stage1_3[182]},
      {stage2_3[114]}
   );
   gpc1_1 gpc7223 (
      {stage1_3[183]},
      {stage2_3[115]}
   );
   gpc1_1 gpc7224 (
      {stage1_3[184]},
      {stage2_3[116]}
   );
   gpc1_1 gpc7225 (
      {stage1_3[185]},
      {stage2_3[117]}
   );
   gpc1_1 gpc7226 (
      {stage1_3[186]},
      {stage2_3[118]}
   );
   gpc1_1 gpc7227 (
      {stage1_3[187]},
      {stage2_3[119]}
   );
   gpc1_1 gpc7228 (
      {stage1_3[188]},
      {stage2_3[120]}
   );
   gpc1_1 gpc7229 (
      {stage1_3[189]},
      {stage2_3[121]}
   );
   gpc1_1 gpc7230 (
      {stage1_3[190]},
      {stage2_3[122]}
   );
   gpc1_1 gpc7231 (
      {stage1_3[191]},
      {stage2_3[123]}
   );
   gpc1_1 gpc7232 (
      {stage1_3[192]},
      {stage2_3[124]}
   );
   gpc1_1 gpc7233 (
      {stage1_3[193]},
      {stage2_3[125]}
   );
   gpc1_1 gpc7234 (
      {stage1_3[194]},
      {stage2_3[126]}
   );
   gpc1_1 gpc7235 (
      {stage1_3[195]},
      {stage2_3[127]}
   );
   gpc1_1 gpc7236 (
      {stage1_3[196]},
      {stage2_3[128]}
   );
   gpc1_1 gpc7237 (
      {stage1_3[197]},
      {stage2_3[129]}
   );
   gpc1_1 gpc7238 (
      {stage1_3[198]},
      {stage2_3[130]}
   );
   gpc1_1 gpc7239 (
      {stage1_3[199]},
      {stage2_3[131]}
   );
   gpc1_1 gpc7240 (
      {stage1_3[200]},
      {stage2_3[132]}
   );
   gpc1_1 gpc7241 (
      {stage1_3[201]},
      {stage2_3[133]}
   );
   gpc1_1 gpc7242 (
      {stage1_3[202]},
      {stage2_3[134]}
   );
   gpc1_1 gpc7243 (
      {stage1_3[203]},
      {stage2_3[135]}
   );
   gpc1_1 gpc7244 (
      {stage1_3[204]},
      {stage2_3[136]}
   );
   gpc1_1 gpc7245 (
      {stage1_3[205]},
      {stage2_3[137]}
   );
   gpc1_1 gpc7246 (
      {stage1_3[206]},
      {stage2_3[138]}
   );
   gpc1_1 gpc7247 (
      {stage1_3[207]},
      {stage2_3[139]}
   );
   gpc1_1 gpc7248 (
      {stage1_3[208]},
      {stage2_3[140]}
   );
   gpc1_1 gpc7249 (
      {stage1_3[209]},
      {stage2_3[141]}
   );
   gpc1_1 gpc7250 (
      {stage1_3[210]},
      {stage2_3[142]}
   );
   gpc1_1 gpc7251 (
      {stage1_3[211]},
      {stage2_3[143]}
   );
   gpc1_1 gpc7252 (
      {stage1_3[212]},
      {stage2_3[144]}
   );
   gpc1_1 gpc7253 (
      {stage1_3[213]},
      {stage2_3[145]}
   );
   gpc1_1 gpc7254 (
      {stage1_3[214]},
      {stage2_3[146]}
   );
   gpc1_1 gpc7255 (
      {stage1_3[215]},
      {stage2_3[147]}
   );
   gpc1_1 gpc7256 (
      {stage1_3[216]},
      {stage2_3[148]}
   );
   gpc1_1 gpc7257 (
      {stage1_3[217]},
      {stage2_3[149]}
   );
   gpc1_1 gpc7258 (
      {stage1_3[218]},
      {stage2_3[150]}
   );
   gpc1_1 gpc7259 (
      {stage1_3[219]},
      {stage2_3[151]}
   );
   gpc1_1 gpc7260 (
      {stage1_3[220]},
      {stage2_3[152]}
   );
   gpc1_1 gpc7261 (
      {stage1_3[221]},
      {stage2_3[153]}
   );
   gpc1_1 gpc7262 (
      {stage1_3[222]},
      {stage2_3[154]}
   );
   gpc1_1 gpc7263 (
      {stage1_3[223]},
      {stage2_3[155]}
   );
   gpc1_1 gpc7264 (
      {stage1_3[224]},
      {stage2_3[156]}
   );
   gpc1_1 gpc7265 (
      {stage1_3[225]},
      {stage2_3[157]}
   );
   gpc1_1 gpc7266 (
      {stage1_3[226]},
      {stage2_3[158]}
   );
   gpc1_1 gpc7267 (
      {stage1_3[227]},
      {stage2_3[159]}
   );
   gpc1_1 gpc7268 (
      {stage1_3[228]},
      {stage2_3[160]}
   );
   gpc1_1 gpc7269 (
      {stage1_3[229]},
      {stage2_3[161]}
   );
   gpc1_1 gpc7270 (
      {stage1_3[230]},
      {stage2_3[162]}
   );
   gpc1_1 gpc7271 (
      {stage1_3[231]},
      {stage2_3[163]}
   );
   gpc1_1 gpc7272 (
      {stage1_3[232]},
      {stage2_3[164]}
   );
   gpc1_1 gpc7273 (
      {stage1_3[233]},
      {stage2_3[165]}
   );
   gpc1_1 gpc7274 (
      {stage1_3[234]},
      {stage2_3[166]}
   );
   gpc1_1 gpc7275 (
      {stage1_3[235]},
      {stage2_3[167]}
   );
   gpc1_1 gpc7276 (
      {stage1_3[236]},
      {stage2_3[168]}
   );
   gpc1_1 gpc7277 (
      {stage1_3[237]},
      {stage2_3[169]}
   );
   gpc1_1 gpc7278 (
      {stage1_3[238]},
      {stage2_3[170]}
   );
   gpc1_1 gpc7279 (
      {stage1_3[239]},
      {stage2_3[171]}
   );
   gpc1_1 gpc7280 (
      {stage1_3[240]},
      {stage2_3[172]}
   );
   gpc1_1 gpc7281 (
      {stage1_3[241]},
      {stage2_3[173]}
   );
   gpc1_1 gpc7282 (
      {stage1_3[242]},
      {stage2_3[174]}
   );
   gpc1_1 gpc7283 (
      {stage1_3[243]},
      {stage2_3[175]}
   );
   gpc1_1 gpc7284 (
      {stage1_3[244]},
      {stage2_3[176]}
   );
   gpc1_1 gpc7285 (
      {stage1_3[245]},
      {stage2_3[177]}
   );
   gpc1_1 gpc7286 (
      {stage1_3[246]},
      {stage2_3[178]}
   );
   gpc1_1 gpc7287 (
      {stage1_3[247]},
      {stage2_3[179]}
   );
   gpc1_1 gpc7288 (
      {stage1_3[248]},
      {stage2_3[180]}
   );
   gpc1_1 gpc7289 (
      {stage1_3[249]},
      {stage2_3[181]}
   );
   gpc1_1 gpc7290 (
      {stage1_3[250]},
      {stage2_3[182]}
   );
   gpc1_1 gpc7291 (
      {stage1_3[251]},
      {stage2_3[183]}
   );
   gpc1_1 gpc7292 (
      {stage1_3[252]},
      {stage2_3[184]}
   );
   gpc1_1 gpc7293 (
      {stage1_3[253]},
      {stage2_3[185]}
   );
   gpc1_1 gpc7294 (
      {stage1_3[254]},
      {stage2_3[186]}
   );
   gpc1_1 gpc7295 (
      {stage1_3[255]},
      {stage2_3[187]}
   );
   gpc1_1 gpc7296 (
      {stage1_3[256]},
      {stage2_3[188]}
   );
   gpc1_1 gpc7297 (
      {stage1_3[257]},
      {stage2_3[189]}
   );
   gpc1_1 gpc7298 (
      {stage1_3[258]},
      {stage2_3[190]}
   );
   gpc1_1 gpc7299 (
      {stage1_3[259]},
      {stage2_3[191]}
   );
   gpc1_1 gpc7300 (
      {stage1_3[260]},
      {stage2_3[192]}
   );
   gpc1_1 gpc7301 (
      {stage1_3[261]},
      {stage2_3[193]}
   );
   gpc1_1 gpc7302 (
      {stage1_3[262]},
      {stage2_3[194]}
   );
   gpc1_1 gpc7303 (
      {stage1_3[263]},
      {stage2_3[195]}
   );
   gpc1_1 gpc7304 (
      {stage1_3[264]},
      {stage2_3[196]}
   );
   gpc1_1 gpc7305 (
      {stage1_3[265]},
      {stage2_3[197]}
   );
   gpc1_1 gpc7306 (
      {stage1_3[266]},
      {stage2_3[198]}
   );
   gpc1_1 gpc7307 (
      {stage1_3[267]},
      {stage2_3[199]}
   );
   gpc1_1 gpc7308 (
      {stage1_3[268]},
      {stage2_3[200]}
   );
   gpc1_1 gpc7309 (
      {stage1_3[269]},
      {stage2_3[201]}
   );
   gpc1_1 gpc7310 (
      {stage1_3[270]},
      {stage2_3[202]}
   );
   gpc1_1 gpc7311 (
      {stage1_3[271]},
      {stage2_3[203]}
   );
   gpc1_1 gpc7312 (
      {stage1_3[272]},
      {stage2_3[204]}
   );
   gpc1_1 gpc7313 (
      {stage1_3[273]},
      {stage2_3[205]}
   );
   gpc1_1 gpc7314 (
      {stage1_3[274]},
      {stage2_3[206]}
   );
   gpc1_1 gpc7315 (
      {stage1_3[275]},
      {stage2_3[207]}
   );
   gpc1_1 gpc7316 (
      {stage1_3[276]},
      {stage2_3[208]}
   );
   gpc1_1 gpc7317 (
      {stage1_3[277]},
      {stage2_3[209]}
   );
   gpc1_1 gpc7318 (
      {stage1_3[278]},
      {stage2_3[210]}
   );
   gpc1_1 gpc7319 (
      {stage1_3[279]},
      {stage2_3[211]}
   );
   gpc1_1 gpc7320 (
      {stage1_3[280]},
      {stage2_3[212]}
   );
   gpc1_1 gpc7321 (
      {stage1_3[281]},
      {stage2_3[213]}
   );
   gpc1_1 gpc7322 (
      {stage1_3[282]},
      {stage2_3[214]}
   );
   gpc1_1 gpc7323 (
      {stage1_3[283]},
      {stage2_3[215]}
   );
   gpc1_1 gpc7324 (
      {stage1_3[284]},
      {stage2_3[216]}
   );
   gpc1_1 gpc7325 (
      {stage1_3[285]},
      {stage2_3[217]}
   );
   gpc1_1 gpc7326 (
      {stage1_3[286]},
      {stage2_3[218]}
   );
   gpc1_1 gpc7327 (
      {stage1_3[287]},
      {stage2_3[219]}
   );
   gpc1_1 gpc7328 (
      {stage1_3[288]},
      {stage2_3[220]}
   );
   gpc1_1 gpc7329 (
      {stage1_3[289]},
      {stage2_3[221]}
   );
   gpc1_1 gpc7330 (
      {stage1_3[290]},
      {stage2_3[222]}
   );
   gpc1_1 gpc7331 (
      {stage1_3[291]},
      {stage2_3[223]}
   );
   gpc1_1 gpc7332 (
      {stage1_3[292]},
      {stage2_3[224]}
   );
   gpc1_1 gpc7333 (
      {stage1_3[293]},
      {stage2_3[225]}
   );
   gpc1_1 gpc7334 (
      {stage1_3[294]},
      {stage2_3[226]}
   );
   gpc1_1 gpc7335 (
      {stage1_3[295]},
      {stage2_3[227]}
   );
   gpc1_1 gpc7336 (
      {stage1_3[296]},
      {stage2_3[228]}
   );
   gpc1_1 gpc7337 (
      {stage1_3[297]},
      {stage2_3[229]}
   );
   gpc1_1 gpc7338 (
      {stage1_3[298]},
      {stage2_3[230]}
   );
   gpc1_1 gpc7339 (
      {stage1_3[299]},
      {stage2_3[231]}
   );
   gpc1_1 gpc7340 (
      {stage1_3[300]},
      {stage2_3[232]}
   );
   gpc1_1 gpc7341 (
      {stage1_3[301]},
      {stage2_3[233]}
   );
   gpc1_1 gpc7342 (
      {stage1_3[302]},
      {stage2_3[234]}
   );
   gpc1_1 gpc7343 (
      {stage1_3[303]},
      {stage2_3[235]}
   );
   gpc1_1 gpc7344 (
      {stage1_3[304]},
      {stage2_3[236]}
   );
   gpc1_1 gpc7345 (
      {stage1_3[305]},
      {stage2_3[237]}
   );
   gpc1_1 gpc7346 (
      {stage1_3[306]},
      {stage2_3[238]}
   );
   gpc1_1 gpc7347 (
      {stage1_3[307]},
      {stage2_3[239]}
   );
   gpc1_1 gpc7348 (
      {stage1_3[308]},
      {stage2_3[240]}
   );
   gpc1_1 gpc7349 (
      {stage1_3[309]},
      {stage2_3[241]}
   );
   gpc1_1 gpc7350 (
      {stage1_3[310]},
      {stage2_3[242]}
   );
   gpc1_1 gpc7351 (
      {stage1_3[311]},
      {stage2_3[243]}
   );
   gpc1_1 gpc7352 (
      {stage1_3[312]},
      {stage2_3[244]}
   );
   gpc1_1 gpc7353 (
      {stage1_3[313]},
      {stage2_3[245]}
   );
   gpc1_1 gpc7354 (
      {stage1_3[314]},
      {stage2_3[246]}
   );
   gpc1_1 gpc7355 (
      {stage1_3[315]},
      {stage2_3[247]}
   );
   gpc1_1 gpc7356 (
      {stage1_3[316]},
      {stage2_3[248]}
   );
   gpc1_1 gpc7357 (
      {stage1_3[317]},
      {stage2_3[249]}
   );
   gpc1_1 gpc7358 (
      {stage1_3[318]},
      {stage2_3[250]}
   );
   gpc1_1 gpc7359 (
      {stage1_3[319]},
      {stage2_3[251]}
   );
   gpc1_1 gpc7360 (
      {stage1_3[320]},
      {stage2_3[252]}
   );
   gpc1_1 gpc7361 (
      {stage1_3[321]},
      {stage2_3[253]}
   );
   gpc1_1 gpc7362 (
      {stage1_4[247]},
      {stage2_4[89]}
   );
   gpc1_1 gpc7363 (
      {stage1_4[248]},
      {stage2_4[90]}
   );
   gpc1_1 gpc7364 (
      {stage1_4[249]},
      {stage2_4[91]}
   );
   gpc1_1 gpc7365 (
      {stage1_4[250]},
      {stage2_4[92]}
   );
   gpc1_1 gpc7366 (
      {stage1_5[188]},
      {stage2_5[83]}
   );
   gpc1_1 gpc7367 (
      {stage1_5[189]},
      {stage2_5[84]}
   );
   gpc1_1 gpc7368 (
      {stage1_5[190]},
      {stage2_5[85]}
   );
   gpc1_1 gpc7369 (
      {stage1_5[191]},
      {stage2_5[86]}
   );
   gpc1_1 gpc7370 (
      {stage1_5[192]},
      {stage2_5[87]}
   );
   gpc1_1 gpc7371 (
      {stage1_5[193]},
      {stage2_5[88]}
   );
   gpc1_1 gpc7372 (
      {stage1_5[194]},
      {stage2_5[89]}
   );
   gpc1_1 gpc7373 (
      {stage1_5[195]},
      {stage2_5[90]}
   );
   gpc1_1 gpc7374 (
      {stage1_5[196]},
      {stage2_5[91]}
   );
   gpc1_1 gpc7375 (
      {stage1_5[197]},
      {stage2_5[92]}
   );
   gpc1_1 gpc7376 (
      {stage1_5[198]},
      {stage2_5[93]}
   );
   gpc1_1 gpc7377 (
      {stage1_5[199]},
      {stage2_5[94]}
   );
   gpc1_1 gpc7378 (
      {stage1_5[200]},
      {stage2_5[95]}
   );
   gpc1_1 gpc7379 (
      {stage1_5[201]},
      {stage2_5[96]}
   );
   gpc1_1 gpc7380 (
      {stage1_5[202]},
      {stage2_5[97]}
   );
   gpc1_1 gpc7381 (
      {stage1_5[203]},
      {stage2_5[98]}
   );
   gpc1_1 gpc7382 (
      {stage1_5[204]},
      {stage2_5[99]}
   );
   gpc1_1 gpc7383 (
      {stage1_5[205]},
      {stage2_5[100]}
   );
   gpc1_1 gpc7384 (
      {stage1_5[206]},
      {stage2_5[101]}
   );
   gpc1_1 gpc7385 (
      {stage1_5[207]},
      {stage2_5[102]}
   );
   gpc1_1 gpc7386 (
      {stage1_5[208]},
      {stage2_5[103]}
   );
   gpc1_1 gpc7387 (
      {stage1_5[209]},
      {stage2_5[104]}
   );
   gpc1_1 gpc7388 (
      {stage1_5[210]},
      {stage2_5[105]}
   );
   gpc1_1 gpc7389 (
      {stage1_5[211]},
      {stage2_5[106]}
   );
   gpc1_1 gpc7390 (
      {stage1_5[212]},
      {stage2_5[107]}
   );
   gpc1_1 gpc7391 (
      {stage1_5[213]},
      {stage2_5[108]}
   );
   gpc1_1 gpc7392 (
      {stage1_5[214]},
      {stage2_5[109]}
   );
   gpc1_1 gpc7393 (
      {stage1_5[215]},
      {stage2_5[110]}
   );
   gpc1_1 gpc7394 (
      {stage1_5[216]},
      {stage2_5[111]}
   );
   gpc1_1 gpc7395 (
      {stage1_6[135]},
      {stage2_6[76]}
   );
   gpc1_1 gpc7396 (
      {stage1_6[136]},
      {stage2_6[77]}
   );
   gpc1_1 gpc7397 (
      {stage1_6[137]},
      {stage2_6[78]}
   );
   gpc1_1 gpc7398 (
      {stage1_6[138]},
      {stage2_6[79]}
   );
   gpc1_1 gpc7399 (
      {stage1_6[139]},
      {stage2_6[80]}
   );
   gpc1_1 gpc7400 (
      {stage1_6[140]},
      {stage2_6[81]}
   );
   gpc1_1 gpc7401 (
      {stage1_6[141]},
      {stage2_6[82]}
   );
   gpc1_1 gpc7402 (
      {stage1_6[142]},
      {stage2_6[83]}
   );
   gpc1_1 gpc7403 (
      {stage1_6[143]},
      {stage2_6[84]}
   );
   gpc1_1 gpc7404 (
      {stage1_6[144]},
      {stage2_6[85]}
   );
   gpc1_1 gpc7405 (
      {stage1_6[145]},
      {stage2_6[86]}
   );
   gpc1_1 gpc7406 (
      {stage1_6[146]},
      {stage2_6[87]}
   );
   gpc1_1 gpc7407 (
      {stage1_6[147]},
      {stage2_6[88]}
   );
   gpc1_1 gpc7408 (
      {stage1_6[148]},
      {stage2_6[89]}
   );
   gpc1_1 gpc7409 (
      {stage1_6[149]},
      {stage2_6[90]}
   );
   gpc1_1 gpc7410 (
      {stage1_6[150]},
      {stage2_6[91]}
   );
   gpc1_1 gpc7411 (
      {stage1_6[151]},
      {stage2_6[92]}
   );
   gpc1_1 gpc7412 (
      {stage1_6[152]},
      {stage2_6[93]}
   );
   gpc1_1 gpc7413 (
      {stage1_6[153]},
      {stage2_6[94]}
   );
   gpc1_1 gpc7414 (
      {stage1_6[154]},
      {stage2_6[95]}
   );
   gpc1_1 gpc7415 (
      {stage1_6[155]},
      {stage2_6[96]}
   );
   gpc1_1 gpc7416 (
      {stage1_6[156]},
      {stage2_6[97]}
   );
   gpc1_1 gpc7417 (
      {stage1_6[157]},
      {stage2_6[98]}
   );
   gpc1_1 gpc7418 (
      {stage1_6[158]},
      {stage2_6[99]}
   );
   gpc1_1 gpc7419 (
      {stage1_6[159]},
      {stage2_6[100]}
   );
   gpc1_1 gpc7420 (
      {stage1_6[160]},
      {stage2_6[101]}
   );
   gpc1_1 gpc7421 (
      {stage1_6[161]},
      {stage2_6[102]}
   );
   gpc1_1 gpc7422 (
      {stage1_6[162]},
      {stage2_6[103]}
   );
   gpc1_1 gpc7423 (
      {stage1_6[163]},
      {stage2_6[104]}
   );
   gpc1_1 gpc7424 (
      {stage1_6[164]},
      {stage2_6[105]}
   );
   gpc1_1 gpc7425 (
      {stage1_6[165]},
      {stage2_6[106]}
   );
   gpc1_1 gpc7426 (
      {stage1_6[166]},
      {stage2_6[107]}
   );
   gpc1_1 gpc7427 (
      {stage1_6[167]},
      {stage2_6[108]}
   );
   gpc1_1 gpc7428 (
      {stage1_6[168]},
      {stage2_6[109]}
   );
   gpc1_1 gpc7429 (
      {stage1_6[169]},
      {stage2_6[110]}
   );
   gpc1_1 gpc7430 (
      {stage1_6[170]},
      {stage2_6[111]}
   );
   gpc1_1 gpc7431 (
      {stage1_6[171]},
      {stage2_6[112]}
   );
   gpc1_1 gpc7432 (
      {stage1_6[172]},
      {stage2_6[113]}
   );
   gpc1_1 gpc7433 (
      {stage1_6[173]},
      {stage2_6[114]}
   );
   gpc1_1 gpc7434 (
      {stage1_6[174]},
      {stage2_6[115]}
   );
   gpc1_1 gpc7435 (
      {stage1_6[175]},
      {stage2_6[116]}
   );
   gpc1_1 gpc7436 (
      {stage1_6[176]},
      {stage2_6[117]}
   );
   gpc1_1 gpc7437 (
      {stage1_6[177]},
      {stage2_6[118]}
   );
   gpc1_1 gpc7438 (
      {stage1_6[178]},
      {stage2_6[119]}
   );
   gpc1_1 gpc7439 (
      {stage1_6[179]},
      {stage2_6[120]}
   );
   gpc1_1 gpc7440 (
      {stage1_8[168]},
      {stage2_8[102]}
   );
   gpc1_1 gpc7441 (
      {stage1_8[169]},
      {stage2_8[103]}
   );
   gpc1_1 gpc7442 (
      {stage1_8[170]},
      {stage2_8[104]}
   );
   gpc1_1 gpc7443 (
      {stage1_8[171]},
      {stage2_8[105]}
   );
   gpc1_1 gpc7444 (
      {stage1_8[172]},
      {stage2_8[106]}
   );
   gpc1_1 gpc7445 (
      {stage1_8[173]},
      {stage2_8[107]}
   );
   gpc1_1 gpc7446 (
      {stage1_8[174]},
      {stage2_8[108]}
   );
   gpc1_1 gpc7447 (
      {stage1_8[175]},
      {stage2_8[109]}
   );
   gpc1_1 gpc7448 (
      {stage1_8[176]},
      {stage2_8[110]}
   );
   gpc1_1 gpc7449 (
      {stage1_8[177]},
      {stage2_8[111]}
   );
   gpc1_1 gpc7450 (
      {stage1_8[178]},
      {stage2_8[112]}
   );
   gpc1_1 gpc7451 (
      {stage1_8[179]},
      {stage2_8[113]}
   );
   gpc1_1 gpc7452 (
      {stage1_8[180]},
      {stage2_8[114]}
   );
   gpc1_1 gpc7453 (
      {stage1_8[181]},
      {stage2_8[115]}
   );
   gpc1_1 gpc7454 (
      {stage1_8[182]},
      {stage2_8[116]}
   );
   gpc1_1 gpc7455 (
      {stage1_8[183]},
      {stage2_8[117]}
   );
   gpc1_1 gpc7456 (
      {stage1_8[184]},
      {stage2_8[118]}
   );
   gpc1_1 gpc7457 (
      {stage1_8[185]},
      {stage2_8[119]}
   );
   gpc1_1 gpc7458 (
      {stage1_8[186]},
      {stage2_8[120]}
   );
   gpc1_1 gpc7459 (
      {stage1_8[187]},
      {stage2_8[121]}
   );
   gpc1_1 gpc7460 (
      {stage1_8[188]},
      {stage2_8[122]}
   );
   gpc1_1 gpc7461 (
      {stage1_8[189]},
      {stage2_8[123]}
   );
   gpc1_1 gpc7462 (
      {stage1_8[190]},
      {stage2_8[124]}
   );
   gpc1_1 gpc7463 (
      {stage1_8[191]},
      {stage2_8[125]}
   );
   gpc1_1 gpc7464 (
      {stage1_8[192]},
      {stage2_8[126]}
   );
   gpc1_1 gpc7465 (
      {stage1_8[193]},
      {stage2_8[127]}
   );
   gpc1_1 gpc7466 (
      {stage1_8[194]},
      {stage2_8[128]}
   );
   gpc1_1 gpc7467 (
      {stage1_8[195]},
      {stage2_8[129]}
   );
   gpc1_1 gpc7468 (
      {stage1_8[196]},
      {stage2_8[130]}
   );
   gpc1_1 gpc7469 (
      {stage1_8[197]},
      {stage2_8[131]}
   );
   gpc1_1 gpc7470 (
      {stage1_8[198]},
      {stage2_8[132]}
   );
   gpc1_1 gpc7471 (
      {stage1_8[199]},
      {stage2_8[133]}
   );
   gpc1_1 gpc7472 (
      {stage1_8[200]},
      {stage2_8[134]}
   );
   gpc1_1 gpc7473 (
      {stage1_8[201]},
      {stage2_8[135]}
   );
   gpc1_1 gpc7474 (
      {stage1_8[202]},
      {stage2_8[136]}
   );
   gpc1_1 gpc7475 (
      {stage1_8[203]},
      {stage2_8[137]}
   );
   gpc1_1 gpc7476 (
      {stage1_8[204]},
      {stage2_8[138]}
   );
   gpc1_1 gpc7477 (
      {stage1_8[205]},
      {stage2_8[139]}
   );
   gpc1_1 gpc7478 (
      {stage1_8[206]},
      {stage2_8[140]}
   );
   gpc1_1 gpc7479 (
      {stage1_8[207]},
      {stage2_8[141]}
   );
   gpc1_1 gpc7480 (
      {stage1_8[208]},
      {stage2_8[142]}
   );
   gpc1_1 gpc7481 (
      {stage1_8[209]},
      {stage2_8[143]}
   );
   gpc1_1 gpc7482 (
      {stage1_8[210]},
      {stage2_8[144]}
   );
   gpc1_1 gpc7483 (
      {stage1_8[211]},
      {stage2_8[145]}
   );
   gpc1_1 gpc7484 (
      {stage1_8[212]},
      {stage2_8[146]}
   );
   gpc1_1 gpc7485 (
      {stage1_8[213]},
      {stage2_8[147]}
   );
   gpc1_1 gpc7486 (
      {stage1_8[214]},
      {stage2_8[148]}
   );
   gpc1_1 gpc7487 (
      {stage1_8[215]},
      {stage2_8[149]}
   );
   gpc1_1 gpc7488 (
      {stage1_8[216]},
      {stage2_8[150]}
   );
   gpc1_1 gpc7489 (
      {stage1_8[217]},
      {stage2_8[151]}
   );
   gpc1_1 gpc7490 (
      {stage1_8[218]},
      {stage2_8[152]}
   );
   gpc1_1 gpc7491 (
      {stage1_8[219]},
      {stage2_8[153]}
   );
   gpc1_1 gpc7492 (
      {stage1_8[220]},
      {stage2_8[154]}
   );
   gpc1_1 gpc7493 (
      {stage1_8[221]},
      {stage2_8[155]}
   );
   gpc1_1 gpc7494 (
      {stage1_8[222]},
      {stage2_8[156]}
   );
   gpc1_1 gpc7495 (
      {stage1_8[223]},
      {stage2_8[157]}
   );
   gpc1_1 gpc7496 (
      {stage1_8[224]},
      {stage2_8[158]}
   );
   gpc1_1 gpc7497 (
      {stage1_8[225]},
      {stage2_8[159]}
   );
   gpc1_1 gpc7498 (
      {stage1_8[226]},
      {stage2_8[160]}
   );
   gpc1_1 gpc7499 (
      {stage1_8[227]},
      {stage2_8[161]}
   );
   gpc1_1 gpc7500 (
      {stage1_8[228]},
      {stage2_8[162]}
   );
   gpc1_1 gpc7501 (
      {stage1_8[229]},
      {stage2_8[163]}
   );
   gpc1_1 gpc7502 (
      {stage1_8[230]},
      {stage2_8[164]}
   );
   gpc1_1 gpc7503 (
      {stage1_8[231]},
      {stage2_8[165]}
   );
   gpc1_1 gpc7504 (
      {stage1_8[232]},
      {stage2_8[166]}
   );
   gpc1_1 gpc7505 (
      {stage1_8[233]},
      {stage2_8[167]}
   );
   gpc1_1 gpc7506 (
      {stage1_8[234]},
      {stage2_8[168]}
   );
   gpc1_1 gpc7507 (
      {stage1_8[235]},
      {stage2_8[169]}
   );
   gpc1_1 gpc7508 (
      {stage1_8[236]},
      {stage2_8[170]}
   );
   gpc1_1 gpc7509 (
      {stage1_8[237]},
      {stage2_8[171]}
   );
   gpc1_1 gpc7510 (
      {stage1_8[238]},
      {stage2_8[172]}
   );
   gpc1_1 gpc7511 (
      {stage1_9[360]},
      {stage2_9[102]}
   );
   gpc1_1 gpc7512 (
      {stage1_9[361]},
      {stage2_9[103]}
   );
   gpc1_1 gpc7513 (
      {stage1_9[362]},
      {stage2_9[104]}
   );
   gpc1_1 gpc7514 (
      {stage1_10[101]},
      {stage2_10[82]}
   );
   gpc1_1 gpc7515 (
      {stage1_10[102]},
      {stage2_10[83]}
   );
   gpc1_1 gpc7516 (
      {stage1_10[103]},
      {stage2_10[84]}
   );
   gpc1_1 gpc7517 (
      {stage1_10[104]},
      {stage2_10[85]}
   );
   gpc1_1 gpc7518 (
      {stage1_10[105]},
      {stage2_10[86]}
   );
   gpc1_1 gpc7519 (
      {stage1_10[106]},
      {stage2_10[87]}
   );
   gpc1_1 gpc7520 (
      {stage1_10[107]},
      {stage2_10[88]}
   );
   gpc1_1 gpc7521 (
      {stage1_10[108]},
      {stage2_10[89]}
   );
   gpc1_1 gpc7522 (
      {stage1_10[109]},
      {stage2_10[90]}
   );
   gpc1_1 gpc7523 (
      {stage1_10[110]},
      {stage2_10[91]}
   );
   gpc1_1 gpc7524 (
      {stage1_10[111]},
      {stage2_10[92]}
   );
   gpc1_1 gpc7525 (
      {stage1_10[112]},
      {stage2_10[93]}
   );
   gpc1_1 gpc7526 (
      {stage1_10[113]},
      {stage2_10[94]}
   );
   gpc1_1 gpc7527 (
      {stage1_10[114]},
      {stage2_10[95]}
   );
   gpc1_1 gpc7528 (
      {stage1_10[115]},
      {stage2_10[96]}
   );
   gpc1_1 gpc7529 (
      {stage1_10[116]},
      {stage2_10[97]}
   );
   gpc1_1 gpc7530 (
      {stage1_10[117]},
      {stage2_10[98]}
   );
   gpc1_1 gpc7531 (
      {stage1_10[118]},
      {stage2_10[99]}
   );
   gpc1_1 gpc7532 (
      {stage1_10[119]},
      {stage2_10[100]}
   );
   gpc1_1 gpc7533 (
      {stage1_10[120]},
      {stage2_10[101]}
   );
   gpc1_1 gpc7534 (
      {stage1_10[121]},
      {stage2_10[102]}
   );
   gpc1_1 gpc7535 (
      {stage1_10[122]},
      {stage2_10[103]}
   );
   gpc1_1 gpc7536 (
      {stage1_10[123]},
      {stage2_10[104]}
   );
   gpc1_1 gpc7537 (
      {stage1_10[124]},
      {stage2_10[105]}
   );
   gpc1_1 gpc7538 (
      {stage1_10[125]},
      {stage2_10[106]}
   );
   gpc1_1 gpc7539 (
      {stage1_10[126]},
      {stage2_10[107]}
   );
   gpc1_1 gpc7540 (
      {stage1_10[127]},
      {stage2_10[108]}
   );
   gpc1_1 gpc7541 (
      {stage1_10[128]},
      {stage2_10[109]}
   );
   gpc1_1 gpc7542 (
      {stage1_10[129]},
      {stage2_10[110]}
   );
   gpc1_1 gpc7543 (
      {stage1_10[130]},
      {stage2_10[111]}
   );
   gpc1_1 gpc7544 (
      {stage1_10[131]},
      {stage2_10[112]}
   );
   gpc1_1 gpc7545 (
      {stage1_10[132]},
      {stage2_10[113]}
   );
   gpc1_1 gpc7546 (
      {stage1_10[133]},
      {stage2_10[114]}
   );
   gpc1_1 gpc7547 (
      {stage1_10[134]},
      {stage2_10[115]}
   );
   gpc1_1 gpc7548 (
      {stage1_10[135]},
      {stage2_10[116]}
   );
   gpc1_1 gpc7549 (
      {stage1_10[136]},
      {stage2_10[117]}
   );
   gpc1_1 gpc7550 (
      {stage1_10[137]},
      {stage2_10[118]}
   );
   gpc1_1 gpc7551 (
      {stage1_10[138]},
      {stage2_10[119]}
   );
   gpc1_1 gpc7552 (
      {stage1_10[139]},
      {stage2_10[120]}
   );
   gpc1_1 gpc7553 (
      {stage1_10[140]},
      {stage2_10[121]}
   );
   gpc1_1 gpc7554 (
      {stage1_10[141]},
      {stage2_10[122]}
   );
   gpc1_1 gpc7555 (
      {stage1_10[142]},
      {stage2_10[123]}
   );
   gpc1_1 gpc7556 (
      {stage1_10[143]},
      {stage2_10[124]}
   );
   gpc1_1 gpc7557 (
      {stage1_10[144]},
      {stage2_10[125]}
   );
   gpc1_1 gpc7558 (
      {stage1_10[145]},
      {stage2_10[126]}
   );
   gpc1_1 gpc7559 (
      {stage1_10[146]},
      {stage2_10[127]}
   );
   gpc1_1 gpc7560 (
      {stage1_10[147]},
      {stage2_10[128]}
   );
   gpc1_1 gpc7561 (
      {stage1_10[148]},
      {stage2_10[129]}
   );
   gpc1_1 gpc7562 (
      {stage1_10[149]},
      {stage2_10[130]}
   );
   gpc1_1 gpc7563 (
      {stage1_10[150]},
      {stage2_10[131]}
   );
   gpc1_1 gpc7564 (
      {stage1_10[151]},
      {stage2_10[132]}
   );
   gpc1_1 gpc7565 (
      {stage1_10[152]},
      {stage2_10[133]}
   );
   gpc1_1 gpc7566 (
      {stage1_11[307]},
      {stage2_11[125]}
   );
   gpc1_1 gpc7567 (
      {stage1_11[308]},
      {stage2_11[126]}
   );
   gpc1_1 gpc7568 (
      {stage1_11[309]},
      {stage2_11[127]}
   );
   gpc1_1 gpc7569 (
      {stage1_11[310]},
      {stage2_11[128]}
   );
   gpc1_1 gpc7570 (
      {stage1_11[311]},
      {stage2_11[129]}
   );
   gpc1_1 gpc7571 (
      {stage1_11[312]},
      {stage2_11[130]}
   );
   gpc1_1 gpc7572 (
      {stage1_11[313]},
      {stage2_11[131]}
   );
   gpc1_1 gpc7573 (
      {stage1_11[314]},
      {stage2_11[132]}
   );
   gpc1_1 gpc7574 (
      {stage1_11[315]},
      {stage2_11[133]}
   );
   gpc1_1 gpc7575 (
      {stage1_11[316]},
      {stage2_11[134]}
   );
   gpc1_1 gpc7576 (
      {stage1_11[317]},
      {stage2_11[135]}
   );
   gpc1_1 gpc7577 (
      {stage1_12[177]},
      {stage2_12[86]}
   );
   gpc1_1 gpc7578 (
      {stage1_12[178]},
      {stage2_12[87]}
   );
   gpc1_1 gpc7579 (
      {stage1_12[179]},
      {stage2_12[88]}
   );
   gpc1_1 gpc7580 (
      {stage1_12[180]},
      {stage2_12[89]}
   );
   gpc1_1 gpc7581 (
      {stage1_12[181]},
      {stage2_12[90]}
   );
   gpc1_1 gpc7582 (
      {stage1_12[182]},
      {stage2_12[91]}
   );
   gpc1_1 gpc7583 (
      {stage1_12[183]},
      {stage2_12[92]}
   );
   gpc1_1 gpc7584 (
      {stage1_12[184]},
      {stage2_12[93]}
   );
   gpc1_1 gpc7585 (
      {stage1_12[185]},
      {stage2_12[94]}
   );
   gpc1_1 gpc7586 (
      {stage1_12[186]},
      {stage2_12[95]}
   );
   gpc1_1 gpc7587 (
      {stage1_12[187]},
      {stage2_12[96]}
   );
   gpc1_1 gpc7588 (
      {stage1_12[188]},
      {stage2_12[97]}
   );
   gpc1_1 gpc7589 (
      {stage1_12[189]},
      {stage2_12[98]}
   );
   gpc1_1 gpc7590 (
      {stage1_12[190]},
      {stage2_12[99]}
   );
   gpc1_1 gpc7591 (
      {stage1_12[191]},
      {stage2_12[100]}
   );
   gpc1_1 gpc7592 (
      {stage1_12[192]},
      {stage2_12[101]}
   );
   gpc1_1 gpc7593 (
      {stage1_12[193]},
      {stage2_12[102]}
   );
   gpc1_1 gpc7594 (
      {stage1_12[194]},
      {stage2_12[103]}
   );
   gpc1_1 gpc7595 (
      {stage1_12[195]},
      {stage2_12[104]}
   );
   gpc1_1 gpc7596 (
      {stage1_12[196]},
      {stage2_12[105]}
   );
   gpc1_1 gpc7597 (
      {stage1_12[197]},
      {stage2_12[106]}
   );
   gpc1_1 gpc7598 (
      {stage1_12[198]},
      {stage2_12[107]}
   );
   gpc1_1 gpc7599 (
      {stage1_12[199]},
      {stage2_12[108]}
   );
   gpc1_1 gpc7600 (
      {stage1_12[200]},
      {stage2_12[109]}
   );
   gpc1_1 gpc7601 (
      {stage1_12[201]},
      {stage2_12[110]}
   );
   gpc1_1 gpc7602 (
      {stage1_12[202]},
      {stage2_12[111]}
   );
   gpc1_1 gpc7603 (
      {stage1_12[203]},
      {stage2_12[112]}
   );
   gpc1_1 gpc7604 (
      {stage1_12[204]},
      {stage2_12[113]}
   );
   gpc1_1 gpc7605 (
      {stage1_12[205]},
      {stage2_12[114]}
   );
   gpc1_1 gpc7606 (
      {stage1_12[206]},
      {stage2_12[115]}
   );
   gpc1_1 gpc7607 (
      {stage1_12[207]},
      {stage2_12[116]}
   );
   gpc1_1 gpc7608 (
      {stage1_12[208]},
      {stage2_12[117]}
   );
   gpc1_1 gpc7609 (
      {stage1_12[209]},
      {stage2_12[118]}
   );
   gpc1_1 gpc7610 (
      {stage1_12[210]},
      {stage2_12[119]}
   );
   gpc1_1 gpc7611 (
      {stage1_12[211]},
      {stage2_12[120]}
   );
   gpc1_1 gpc7612 (
      {stage1_12[212]},
      {stage2_12[121]}
   );
   gpc1_1 gpc7613 (
      {stage1_12[213]},
      {stage2_12[122]}
   );
   gpc1_1 gpc7614 (
      {stage1_12[214]},
      {stage2_12[123]}
   );
   gpc1_1 gpc7615 (
      {stage1_12[215]},
      {stage2_12[124]}
   );
   gpc1_1 gpc7616 (
      {stage1_12[216]},
      {stage2_12[125]}
   );
   gpc1_1 gpc7617 (
      {stage1_12[217]},
      {stage2_12[126]}
   );
   gpc1_1 gpc7618 (
      {stage1_12[218]},
      {stage2_12[127]}
   );
   gpc1_1 gpc7619 (
      {stage1_13[183]},
      {stage2_13[70]}
   );
   gpc1_1 gpc7620 (
      {stage1_13[184]},
      {stage2_13[71]}
   );
   gpc1_1 gpc7621 (
      {stage1_14[246]},
      {stage2_14[105]}
   );
   gpc1_1 gpc7622 (
      {stage1_14[247]},
      {stage2_14[106]}
   );
   gpc1_1 gpc7623 (
      {stage1_14[248]},
      {stage2_14[107]}
   );
   gpc1_1 gpc7624 (
      {stage1_14[249]},
      {stage2_14[108]}
   );
   gpc1_1 gpc7625 (
      {stage1_14[250]},
      {stage2_14[109]}
   );
   gpc1_1 gpc7626 (
      {stage1_14[251]},
      {stage2_14[110]}
   );
   gpc1_1 gpc7627 (
      {stage1_14[252]},
      {stage2_14[111]}
   );
   gpc1_1 gpc7628 (
      {stage1_14[253]},
      {stage2_14[112]}
   );
   gpc1_1 gpc7629 (
      {stage1_14[254]},
      {stage2_14[113]}
   );
   gpc1_1 gpc7630 (
      {stage1_14[255]},
      {stage2_14[114]}
   );
   gpc1_1 gpc7631 (
      {stage1_15[255]},
      {stage2_15[112]}
   );
   gpc1_1 gpc7632 (
      {stage1_15[256]},
      {stage2_15[113]}
   );
   gpc1_1 gpc7633 (
      {stage1_15[257]},
      {stage2_15[114]}
   );
   gpc1_1 gpc7634 (
      {stage1_16[182]},
      {stage2_16[68]}
   );
   gpc1_1 gpc7635 (
      {stage1_16[183]},
      {stage2_16[69]}
   );
   gpc1_1 gpc7636 (
      {stage1_16[184]},
      {stage2_16[70]}
   );
   gpc1_1 gpc7637 (
      {stage1_16[185]},
      {stage2_16[71]}
   );
   gpc1_1 gpc7638 (
      {stage1_16[186]},
      {stage2_16[72]}
   );
   gpc1_1 gpc7639 (
      {stage1_16[187]},
      {stage2_16[73]}
   );
   gpc1_1 gpc7640 (
      {stage1_16[188]},
      {stage2_16[74]}
   );
   gpc1_1 gpc7641 (
      {stage1_16[189]},
      {stage2_16[75]}
   );
   gpc1_1 gpc7642 (
      {stage1_16[190]},
      {stage2_16[76]}
   );
   gpc1_1 gpc7643 (
      {stage1_16[191]},
      {stage2_16[77]}
   );
   gpc1_1 gpc7644 (
      {stage1_16[192]},
      {stage2_16[78]}
   );
   gpc1_1 gpc7645 (
      {stage1_16[193]},
      {stage2_16[79]}
   );
   gpc1_1 gpc7646 (
      {stage1_16[194]},
      {stage2_16[80]}
   );
   gpc1_1 gpc7647 (
      {stage1_16[195]},
      {stage2_16[81]}
   );
   gpc1_1 gpc7648 (
      {stage1_16[196]},
      {stage2_16[82]}
   );
   gpc1_1 gpc7649 (
      {stage1_16[197]},
      {stage2_16[83]}
   );
   gpc1_1 gpc7650 (
      {stage1_16[198]},
      {stage2_16[84]}
   );
   gpc1_1 gpc7651 (
      {stage1_16[199]},
      {stage2_16[85]}
   );
   gpc1_1 gpc7652 (
      {stage1_16[200]},
      {stage2_16[86]}
   );
   gpc1_1 gpc7653 (
      {stage1_16[201]},
      {stage2_16[87]}
   );
   gpc1_1 gpc7654 (
      {stage1_16[202]},
      {stage2_16[88]}
   );
   gpc1_1 gpc7655 (
      {stage1_16[203]},
      {stage2_16[89]}
   );
   gpc1_1 gpc7656 (
      {stage1_16[204]},
      {stage2_16[90]}
   );
   gpc1_1 gpc7657 (
      {stage1_16[205]},
      {stage2_16[91]}
   );
   gpc1_1 gpc7658 (
      {stage1_16[206]},
      {stage2_16[92]}
   );
   gpc1_1 gpc7659 (
      {stage1_16[207]},
      {stage2_16[93]}
   );
   gpc1_1 gpc7660 (
      {stage1_16[208]},
      {stage2_16[94]}
   );
   gpc1_1 gpc7661 (
      {stage1_16[209]},
      {stage2_16[95]}
   );
   gpc1_1 gpc7662 (
      {stage1_16[210]},
      {stage2_16[96]}
   );
   gpc1_1 gpc7663 (
      {stage1_16[211]},
      {stage2_16[97]}
   );
   gpc1_1 gpc7664 (
      {stage1_16[212]},
      {stage2_16[98]}
   );
   gpc1_1 gpc7665 (
      {stage1_16[213]},
      {stage2_16[99]}
   );
   gpc1_1 gpc7666 (
      {stage1_16[214]},
      {stage2_16[100]}
   );
   gpc1_1 gpc7667 (
      {stage1_16[215]},
      {stage2_16[101]}
   );
   gpc1_1 gpc7668 (
      {stage1_16[216]},
      {stage2_16[102]}
   );
   gpc1_1 gpc7669 (
      {stage1_16[217]},
      {stage2_16[103]}
   );
   gpc1_1 gpc7670 (
      {stage1_16[218]},
      {stage2_16[104]}
   );
   gpc1_1 gpc7671 (
      {stage1_16[219]},
      {stage2_16[105]}
   );
   gpc1_1 gpc7672 (
      {stage1_16[220]},
      {stage2_16[106]}
   );
   gpc1_1 gpc7673 (
      {stage1_16[221]},
      {stage2_16[107]}
   );
   gpc1_1 gpc7674 (
      {stage1_16[222]},
      {stage2_16[108]}
   );
   gpc1_1 gpc7675 (
      {stage1_16[223]},
      {stage2_16[109]}
   );
   gpc1_1 gpc7676 (
      {stage1_18[204]},
      {stage2_18[124]}
   );
   gpc1_1 gpc7677 (
      {stage1_18[205]},
      {stage2_18[125]}
   );
   gpc1_1 gpc7678 (
      {stage1_18[206]},
      {stage2_18[126]}
   );
   gpc1_1 gpc7679 (
      {stage1_18[207]},
      {stage2_18[127]}
   );
   gpc1_1 gpc7680 (
      {stage1_18[208]},
      {stage2_18[128]}
   );
   gpc1_1 gpc7681 (
      {stage1_18[209]},
      {stage2_18[129]}
   );
   gpc1_1 gpc7682 (
      {stage1_18[210]},
      {stage2_18[130]}
   );
   gpc1_1 gpc7683 (
      {stage1_18[211]},
      {stage2_18[131]}
   );
   gpc1_1 gpc7684 (
      {stage1_18[212]},
      {stage2_18[132]}
   );
   gpc1_1 gpc7685 (
      {stage1_18[213]},
      {stage2_18[133]}
   );
   gpc1_1 gpc7686 (
      {stage1_18[214]},
      {stage2_18[134]}
   );
   gpc1_1 gpc7687 (
      {stage1_18[215]},
      {stage2_18[135]}
   );
   gpc1_1 gpc7688 (
      {stage1_18[216]},
      {stage2_18[136]}
   );
   gpc1_1 gpc7689 (
      {stage1_18[217]},
      {stage2_18[137]}
   );
   gpc1_1 gpc7690 (
      {stage1_18[218]},
      {stage2_18[138]}
   );
   gpc1_1 gpc7691 (
      {stage1_18[219]},
      {stage2_18[139]}
   );
   gpc1_1 gpc7692 (
      {stage1_18[220]},
      {stage2_18[140]}
   );
   gpc1_1 gpc7693 (
      {stage1_18[221]},
      {stage2_18[141]}
   );
   gpc1_1 gpc7694 (
      {stage1_18[222]},
      {stage2_18[142]}
   );
   gpc1_1 gpc7695 (
      {stage1_18[223]},
      {stage2_18[143]}
   );
   gpc1_1 gpc7696 (
      {stage1_18[224]},
      {stage2_18[144]}
   );
   gpc1_1 gpc7697 (
      {stage1_18[225]},
      {stage2_18[145]}
   );
   gpc1_1 gpc7698 (
      {stage1_18[226]},
      {stage2_18[146]}
   );
   gpc1_1 gpc7699 (
      {stage1_18[227]},
      {stage2_18[147]}
   );
   gpc1_1 gpc7700 (
      {stage1_18[228]},
      {stage2_18[148]}
   );
   gpc1_1 gpc7701 (
      {stage1_18[229]},
      {stage2_18[149]}
   );
   gpc1_1 gpc7702 (
      {stage1_18[230]},
      {stage2_18[150]}
   );
   gpc1_1 gpc7703 (
      {stage1_18[231]},
      {stage2_18[151]}
   );
   gpc1_1 gpc7704 (
      {stage1_18[232]},
      {stage2_18[152]}
   );
   gpc1_1 gpc7705 (
      {stage1_18[233]},
      {stage2_18[153]}
   );
   gpc1_1 gpc7706 (
      {stage1_18[234]},
      {stage2_18[154]}
   );
   gpc1_1 gpc7707 (
      {stage1_18[235]},
      {stage2_18[155]}
   );
   gpc1_1 gpc7708 (
      {stage1_18[236]},
      {stage2_18[156]}
   );
   gpc1_1 gpc7709 (
      {stage1_18[237]},
      {stage2_18[157]}
   );
   gpc1_1 gpc7710 (
      {stage1_18[238]},
      {stage2_18[158]}
   );
   gpc1_1 gpc7711 (
      {stage1_18[239]},
      {stage2_18[159]}
   );
   gpc1_1 gpc7712 (
      {stage1_18[240]},
      {stage2_18[160]}
   );
   gpc1_1 gpc7713 (
      {stage1_18[241]},
      {stage2_18[161]}
   );
   gpc1_1 gpc7714 (
      {stage1_19[201]},
      {stage2_19[76]}
   );
   gpc1_1 gpc7715 (
      {stage1_19[202]},
      {stage2_19[77]}
   );
   gpc1_1 gpc7716 (
      {stage1_19[203]},
      {stage2_19[78]}
   );
   gpc1_1 gpc7717 (
      {stage1_19[204]},
      {stage2_19[79]}
   );
   gpc1_1 gpc7718 (
      {stage1_19[205]},
      {stage2_19[80]}
   );
   gpc1_1 gpc7719 (
      {stage1_19[206]},
      {stage2_19[81]}
   );
   gpc1_1 gpc7720 (
      {stage1_19[207]},
      {stage2_19[82]}
   );
   gpc1_1 gpc7721 (
      {stage1_19[208]},
      {stage2_19[83]}
   );
   gpc1_1 gpc7722 (
      {stage1_19[209]},
      {stage2_19[84]}
   );
   gpc1_1 gpc7723 (
      {stage1_19[210]},
      {stage2_19[85]}
   );
   gpc1_1 gpc7724 (
      {stage1_19[211]},
      {stage2_19[86]}
   );
   gpc1_1 gpc7725 (
      {stage1_19[212]},
      {stage2_19[87]}
   );
   gpc1_1 gpc7726 (
      {stage1_19[213]},
      {stage2_19[88]}
   );
   gpc1_1 gpc7727 (
      {stage1_19[214]},
      {stage2_19[89]}
   );
   gpc1_1 gpc7728 (
      {stage1_19[215]},
      {stage2_19[90]}
   );
   gpc1_1 gpc7729 (
      {stage1_19[216]},
      {stage2_19[91]}
   );
   gpc1_1 gpc7730 (
      {stage1_19[217]},
      {stage2_19[92]}
   );
   gpc1_1 gpc7731 (
      {stage1_19[218]},
      {stage2_19[93]}
   );
   gpc1_1 gpc7732 (
      {stage1_20[227]},
      {stage2_20[71]}
   );
   gpc1_1 gpc7733 (
      {stage1_20[228]},
      {stage2_20[72]}
   );
   gpc1_1 gpc7734 (
      {stage1_20[229]},
      {stage2_20[73]}
   );
   gpc1_1 gpc7735 (
      {stage1_20[230]},
      {stage2_20[74]}
   );
   gpc1_1 gpc7736 (
      {stage1_20[231]},
      {stage2_20[75]}
   );
   gpc1_1 gpc7737 (
      {stage1_20[232]},
      {stage2_20[76]}
   );
   gpc1_1 gpc7738 (
      {stage1_20[233]},
      {stage2_20[77]}
   );
   gpc1_1 gpc7739 (
      {stage1_20[234]},
      {stage2_20[78]}
   );
   gpc1_1 gpc7740 (
      {stage1_20[235]},
      {stage2_20[79]}
   );
   gpc1_1 gpc7741 (
      {stage1_20[236]},
      {stage2_20[80]}
   );
   gpc1_1 gpc7742 (
      {stage1_20[237]},
      {stage2_20[81]}
   );
   gpc1_1 gpc7743 (
      {stage1_20[238]},
      {stage2_20[82]}
   );
   gpc1_1 gpc7744 (
      {stage1_20[239]},
      {stage2_20[83]}
   );
   gpc1_1 gpc7745 (
      {stage1_20[240]},
      {stage2_20[84]}
   );
   gpc1_1 gpc7746 (
      {stage1_20[241]},
      {stage2_20[85]}
   );
   gpc1_1 gpc7747 (
      {stage1_20[242]},
      {stage2_20[86]}
   );
   gpc1_1 gpc7748 (
      {stage1_20[243]},
      {stage2_20[87]}
   );
   gpc1_1 gpc7749 (
      {stage1_21[186]},
      {stage2_21[93]}
   );
   gpc1_1 gpc7750 (
      {stage1_21[187]},
      {stage2_21[94]}
   );
   gpc1_1 gpc7751 (
      {stage1_21[188]},
      {stage2_21[95]}
   );
   gpc1_1 gpc7752 (
      {stage1_21[189]},
      {stage2_21[96]}
   );
   gpc1_1 gpc7753 (
      {stage1_21[190]},
      {stage2_21[97]}
   );
   gpc1_1 gpc7754 (
      {stage1_21[191]},
      {stage2_21[98]}
   );
   gpc1_1 gpc7755 (
      {stage1_21[192]},
      {stage2_21[99]}
   );
   gpc1_1 gpc7756 (
      {stage1_21[193]},
      {stage2_21[100]}
   );
   gpc1_1 gpc7757 (
      {stage1_21[194]},
      {stage2_21[101]}
   );
   gpc1_1 gpc7758 (
      {stage1_21[195]},
      {stage2_21[102]}
   );
   gpc1_1 gpc7759 (
      {stage1_21[196]},
      {stage2_21[103]}
   );
   gpc1_1 gpc7760 (
      {stage1_21[197]},
      {stage2_21[104]}
   );
   gpc1_1 gpc7761 (
      {stage1_21[198]},
      {stage2_21[105]}
   );
   gpc1_1 gpc7762 (
      {stage1_21[199]},
      {stage2_21[106]}
   );
   gpc1_1 gpc7763 (
      {stage1_21[200]},
      {stage2_21[107]}
   );
   gpc1_1 gpc7764 (
      {stage1_21[201]},
      {stage2_21[108]}
   );
   gpc1_1 gpc7765 (
      {stage1_21[202]},
      {stage2_21[109]}
   );
   gpc1_1 gpc7766 (
      {stage1_21[203]},
      {stage2_21[110]}
   );
   gpc1_1 gpc7767 (
      {stage1_21[204]},
      {stage2_21[111]}
   );
   gpc1_1 gpc7768 (
      {stage1_22[194]},
      {stage2_22[103]}
   );
   gpc1_1 gpc7769 (
      {stage1_22[195]},
      {stage2_22[104]}
   );
   gpc1_1 gpc7770 (
      {stage1_22[196]},
      {stage2_22[105]}
   );
   gpc1_1 gpc7771 (
      {stage1_22[197]},
      {stage2_22[106]}
   );
   gpc1_1 gpc7772 (
      {stage1_22[198]},
      {stage2_22[107]}
   );
   gpc1_1 gpc7773 (
      {stage1_22[199]},
      {stage2_22[108]}
   );
   gpc1_1 gpc7774 (
      {stage1_22[200]},
      {stage2_22[109]}
   );
   gpc1_1 gpc7775 (
      {stage1_23[290]},
      {stage2_23[89]}
   );
   gpc1_1 gpc7776 (
      {stage1_23[291]},
      {stage2_23[90]}
   );
   gpc1_1 gpc7777 (
      {stage1_23[292]},
      {stage2_23[91]}
   );
   gpc1_1 gpc7778 (
      {stage1_23[293]},
      {stage2_23[92]}
   );
   gpc1_1 gpc7779 (
      {stage1_23[294]},
      {stage2_23[93]}
   );
   gpc1_1 gpc7780 (
      {stage1_23[295]},
      {stage2_23[94]}
   );
   gpc1_1 gpc7781 (
      {stage1_23[296]},
      {stage2_23[95]}
   );
   gpc1_1 gpc7782 (
      {stage1_23[297]},
      {stage2_23[96]}
   );
   gpc1_1 gpc7783 (
      {stage1_23[298]},
      {stage2_23[97]}
   );
   gpc1_1 gpc7784 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc7785 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc7786 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc7787 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc7788 (
      {stage1_25[184]},
      {stage2_25[96]}
   );
   gpc1_1 gpc7789 (
      {stage1_25[185]},
      {stage2_25[97]}
   );
   gpc1_1 gpc7790 (
      {stage1_25[186]},
      {stage2_25[98]}
   );
   gpc1_1 gpc7791 (
      {stage1_25[187]},
      {stage2_25[99]}
   );
   gpc1_1 gpc7792 (
      {stage1_25[188]},
      {stage2_25[100]}
   );
   gpc1_1 gpc7793 (
      {stage1_25[189]},
      {stage2_25[101]}
   );
   gpc1_1 gpc7794 (
      {stage1_25[190]},
      {stage2_25[102]}
   );
   gpc1_1 gpc7795 (
      {stage1_25[191]},
      {stage2_25[103]}
   );
   gpc1_1 gpc7796 (
      {stage1_25[192]},
      {stage2_25[104]}
   );
   gpc1_1 gpc7797 (
      {stage1_25[193]},
      {stage2_25[105]}
   );
   gpc1_1 gpc7798 (
      {stage1_25[194]},
      {stage2_25[106]}
   );
   gpc1_1 gpc7799 (
      {stage1_25[195]},
      {stage2_25[107]}
   );
   gpc1_1 gpc7800 (
      {stage1_25[196]},
      {stage2_25[108]}
   );
   gpc1_1 gpc7801 (
      {stage1_25[197]},
      {stage2_25[109]}
   );
   gpc1_1 gpc7802 (
      {stage1_25[198]},
      {stage2_25[110]}
   );
   gpc1_1 gpc7803 (
      {stage1_25[199]},
      {stage2_25[111]}
   );
   gpc1_1 gpc7804 (
      {stage1_25[200]},
      {stage2_25[112]}
   );
   gpc1_1 gpc7805 (
      {stage1_25[201]},
      {stage2_25[113]}
   );
   gpc1_1 gpc7806 (
      {stage1_25[202]},
      {stage2_25[114]}
   );
   gpc1_1 gpc7807 (
      {stage1_25[203]},
      {stage2_25[115]}
   );
   gpc1_1 gpc7808 (
      {stage1_25[204]},
      {stage2_25[116]}
   );
   gpc1_1 gpc7809 (
      {stage1_25[205]},
      {stage2_25[117]}
   );
   gpc1_1 gpc7810 (
      {stage1_25[206]},
      {stage2_25[118]}
   );
   gpc1_1 gpc7811 (
      {stage1_25[207]},
      {stage2_25[119]}
   );
   gpc1_1 gpc7812 (
      {stage1_25[208]},
      {stage2_25[120]}
   );
   gpc1_1 gpc7813 (
      {stage1_25[209]},
      {stage2_25[121]}
   );
   gpc1_1 gpc7814 (
      {stage1_25[210]},
      {stage2_25[122]}
   );
   gpc1_1 gpc7815 (
      {stage1_26[154]},
      {stage2_26[96]}
   );
   gpc1_1 gpc7816 (
      {stage1_26[155]},
      {stage2_26[97]}
   );
   gpc1_1 gpc7817 (
      {stage1_26[156]},
      {stage2_26[98]}
   );
   gpc1_1 gpc7818 (
      {stage1_26[157]},
      {stage2_26[99]}
   );
   gpc1_1 gpc7819 (
      {stage1_26[158]},
      {stage2_26[100]}
   );
   gpc1_1 gpc7820 (
      {stage1_26[159]},
      {stage2_26[101]}
   );
   gpc1_1 gpc7821 (
      {stage1_26[160]},
      {stage2_26[102]}
   );
   gpc1_1 gpc7822 (
      {stage1_26[161]},
      {stage2_26[103]}
   );
   gpc1_1 gpc7823 (
      {stage1_26[162]},
      {stage2_26[104]}
   );
   gpc1_1 gpc7824 (
      {stage1_26[163]},
      {stage2_26[105]}
   );
   gpc1_1 gpc7825 (
      {stage1_26[164]},
      {stage2_26[106]}
   );
   gpc1_1 gpc7826 (
      {stage1_26[165]},
      {stage2_26[107]}
   );
   gpc1_1 gpc7827 (
      {stage1_26[166]},
      {stage2_26[108]}
   );
   gpc1_1 gpc7828 (
      {stage1_26[167]},
      {stage2_26[109]}
   );
   gpc1_1 gpc7829 (
      {stage1_26[168]},
      {stage2_26[110]}
   );
   gpc1_1 gpc7830 (
      {stage1_26[169]},
      {stage2_26[111]}
   );
   gpc1_1 gpc7831 (
      {stage1_26[170]},
      {stage2_26[112]}
   );
   gpc1_1 gpc7832 (
      {stage1_26[171]},
      {stage2_26[113]}
   );
   gpc1_1 gpc7833 (
      {stage1_26[172]},
      {stage2_26[114]}
   );
   gpc1_1 gpc7834 (
      {stage1_26[173]},
      {stage2_26[115]}
   );
   gpc1_1 gpc7835 (
      {stage1_26[174]},
      {stage2_26[116]}
   );
   gpc1_1 gpc7836 (
      {stage1_26[175]},
      {stage2_26[117]}
   );
   gpc1_1 gpc7837 (
      {stage1_26[176]},
      {stage2_26[118]}
   );
   gpc1_1 gpc7838 (
      {stage1_26[177]},
      {stage2_26[119]}
   );
   gpc1_1 gpc7839 (
      {stage1_26[178]},
      {stage2_26[120]}
   );
   gpc1_1 gpc7840 (
      {stage1_26[179]},
      {stage2_26[121]}
   );
   gpc1_1 gpc7841 (
      {stage1_26[180]},
      {stage2_26[122]}
   );
   gpc1_1 gpc7842 (
      {stage1_26[181]},
      {stage2_26[123]}
   );
   gpc1_1 gpc7843 (
      {stage1_26[182]},
      {stage2_26[124]}
   );
   gpc1_1 gpc7844 (
      {stage1_26[183]},
      {stage2_26[125]}
   );
   gpc1_1 gpc7845 (
      {stage1_26[184]},
      {stage2_26[126]}
   );
   gpc1_1 gpc7846 (
      {stage1_26[185]},
      {stage2_26[127]}
   );
   gpc1_1 gpc7847 (
      {stage1_26[186]},
      {stage2_26[128]}
   );
   gpc1_1 gpc7848 (
      {stage1_26[187]},
      {stage2_26[129]}
   );
   gpc1_1 gpc7849 (
      {stage1_26[188]},
      {stage2_26[130]}
   );
   gpc1_1 gpc7850 (
      {stage1_27[211]},
      {stage2_27[85]}
   );
   gpc1_1 gpc7851 (
      {stage1_28[240]},
      {stage2_28[71]}
   );
   gpc1_1 gpc7852 (
      {stage1_28[241]},
      {stage2_28[72]}
   );
   gpc1_1 gpc7853 (
      {stage1_28[242]},
      {stage2_28[73]}
   );
   gpc1_1 gpc7854 (
      {stage1_28[243]},
      {stage2_28[74]}
   );
   gpc1_1 gpc7855 (
      {stage1_28[244]},
      {stage2_28[75]}
   );
   gpc1_1 gpc7856 (
      {stage1_28[245]},
      {stage2_28[76]}
   );
   gpc1_1 gpc7857 (
      {stage1_28[246]},
      {stage2_28[77]}
   );
   gpc1_1 gpc7858 (
      {stage1_28[247]},
      {stage2_28[78]}
   );
   gpc1_1 gpc7859 (
      {stage1_28[248]},
      {stage2_28[79]}
   );
   gpc1_1 gpc7860 (
      {stage1_29[186]},
      {stage2_29[77]}
   );
   gpc1_1 gpc7861 (
      {stage1_29[187]},
      {stage2_29[78]}
   );
   gpc1_1 gpc7862 (
      {stage1_29[188]},
      {stage2_29[79]}
   );
   gpc1_1 gpc7863 (
      {stage1_29[189]},
      {stage2_29[80]}
   );
   gpc1_1 gpc7864 (
      {stage1_29[190]},
      {stage2_29[81]}
   );
   gpc1_1 gpc7865 (
      {stage1_29[191]},
      {stage2_29[82]}
   );
   gpc1_1 gpc7866 (
      {stage1_29[192]},
      {stage2_29[83]}
   );
   gpc1_1 gpc7867 (
      {stage1_29[193]},
      {stage2_29[84]}
   );
   gpc1_1 gpc7868 (
      {stage1_29[194]},
      {stage2_29[85]}
   );
   gpc1_1 gpc7869 (
      {stage1_29[195]},
      {stage2_29[86]}
   );
   gpc1_1 gpc7870 (
      {stage1_29[196]},
      {stage2_29[87]}
   );
   gpc1_1 gpc7871 (
      {stage1_29[197]},
      {stage2_29[88]}
   );
   gpc1_1 gpc7872 (
      {stage1_29[198]},
      {stage2_29[89]}
   );
   gpc1_1 gpc7873 (
      {stage1_29[199]},
      {stage2_29[90]}
   );
   gpc1_1 gpc7874 (
      {stage1_29[200]},
      {stage2_29[91]}
   );
   gpc1_1 gpc7875 (
      {stage1_29[201]},
      {stage2_29[92]}
   );
   gpc1_1 gpc7876 (
      {stage1_29[202]},
      {stage2_29[93]}
   );
   gpc1_1 gpc7877 (
      {stage1_29[203]},
      {stage2_29[94]}
   );
   gpc1_1 gpc7878 (
      {stage1_29[204]},
      {stage2_29[95]}
   );
   gpc1_1 gpc7879 (
      {stage1_29[205]},
      {stage2_29[96]}
   );
   gpc1_1 gpc7880 (
      {stage1_29[206]},
      {stage2_29[97]}
   );
   gpc1_1 gpc7881 (
      {stage1_29[207]},
      {stage2_29[98]}
   );
   gpc1_1 gpc7882 (
      {stage1_29[208]},
      {stage2_29[99]}
   );
   gpc1_1 gpc7883 (
      {stage1_29[209]},
      {stage2_29[100]}
   );
   gpc1_1 gpc7884 (
      {stage1_29[210]},
      {stage2_29[101]}
   );
   gpc1_1 gpc7885 (
      {stage1_29[211]},
      {stage2_29[102]}
   );
   gpc1_1 gpc7886 (
      {stage1_29[212]},
      {stage2_29[103]}
   );
   gpc1_1 gpc7887 (
      {stage1_29[213]},
      {stage2_29[104]}
   );
   gpc1_1 gpc7888 (
      {stage1_29[214]},
      {stage2_29[105]}
   );
   gpc1_1 gpc7889 (
      {stage1_29[215]},
      {stage2_29[106]}
   );
   gpc1_1 gpc7890 (
      {stage1_29[216]},
      {stage2_29[107]}
   );
   gpc1_1 gpc7891 (
      {stage1_29[217]},
      {stage2_29[108]}
   );
   gpc1_1 gpc7892 (
      {stage1_29[218]},
      {stage2_29[109]}
   );
   gpc1_1 gpc7893 (
      {stage1_29[219]},
      {stage2_29[110]}
   );
   gpc1_1 gpc7894 (
      {stage1_29[220]},
      {stage2_29[111]}
   );
   gpc1_1 gpc7895 (
      {stage1_30[232]},
      {stage2_30[99]}
   );
   gpc1_1 gpc7896 (
      {stage1_31[180]},
      {stage2_31[96]}
   );
   gpc1_1 gpc7897 (
      {stage1_31[181]},
      {stage2_31[97]}
   );
   gpc1_1 gpc7898 (
      {stage1_31[182]},
      {stage2_31[98]}
   );
   gpc1_1 gpc7899 (
      {stage1_31[183]},
      {stage2_31[99]}
   );
   gpc1_1 gpc7900 (
      {stage1_31[184]},
      {stage2_31[100]}
   );
   gpc1_1 gpc7901 (
      {stage1_31[185]},
      {stage2_31[101]}
   );
   gpc1_1 gpc7902 (
      {stage1_31[186]},
      {stage2_31[102]}
   );
   gpc1_1 gpc7903 (
      {stage1_31[187]},
      {stage2_31[103]}
   );
   gpc1_1 gpc7904 (
      {stage1_31[188]},
      {stage2_31[104]}
   );
   gpc1_1 gpc7905 (
      {stage1_31[189]},
      {stage2_31[105]}
   );
   gpc1_1 gpc7906 (
      {stage1_31[190]},
      {stage2_31[106]}
   );
   gpc1_1 gpc7907 (
      {stage1_31[191]},
      {stage2_31[107]}
   );
   gpc1_1 gpc7908 (
      {stage1_31[192]},
      {stage2_31[108]}
   );
   gpc1_1 gpc7909 (
      {stage1_31[193]},
      {stage2_31[109]}
   );
   gpc1_1 gpc7910 (
      {stage1_31[194]},
      {stage2_31[110]}
   );
   gpc1_1 gpc7911 (
      {stage1_31[195]},
      {stage2_31[111]}
   );
   gpc1_1 gpc7912 (
      {stage1_31[196]},
      {stage2_31[112]}
   );
   gpc1_1 gpc7913 (
      {stage1_31[197]},
      {stage2_31[113]}
   );
   gpc1_1 gpc7914 (
      {stage1_31[198]},
      {stage2_31[114]}
   );
   gpc1_1 gpc7915 (
      {stage1_31[199]},
      {stage2_31[115]}
   );
   gpc1_1 gpc7916 (
      {stage1_31[200]},
      {stage2_31[116]}
   );
   gpc1_1 gpc7917 (
      {stage1_31[201]},
      {stage2_31[117]}
   );
   gpc1_1 gpc7918 (
      {stage1_31[202]},
      {stage2_31[118]}
   );
   gpc1_1 gpc7919 (
      {stage1_31[203]},
      {stage2_31[119]}
   );
   gpc1_1 gpc7920 (
      {stage1_31[204]},
      {stage2_31[120]}
   );
   gpc1_1 gpc7921 (
      {stage1_31[205]},
      {stage2_31[121]}
   );
   gpc1_1 gpc7922 (
      {stage1_31[206]},
      {stage2_31[122]}
   );
   gpc1_1 gpc7923 (
      {stage1_31[207]},
      {stage2_31[123]}
   );
   gpc1_1 gpc7924 (
      {stage1_31[208]},
      {stage2_31[124]}
   );
   gpc1_1 gpc7925 (
      {stage1_31[209]},
      {stage2_31[125]}
   );
   gpc1_1 gpc7926 (
      {stage1_31[210]},
      {stage2_31[126]}
   );
   gpc1_1 gpc7927 (
      {stage1_31[211]},
      {stage2_31[127]}
   );
   gpc1_1 gpc7928 (
      {stage1_32[404]},
      {stage2_32[107]}
   );
   gpc1_1 gpc7929 (
      {stage1_32[405]},
      {stage2_32[108]}
   );
   gpc1_1 gpc7930 (
      {stage1_32[406]},
      {stage2_32[109]}
   );
   gpc1_1 gpc7931 (
      {stage1_32[407]},
      {stage2_32[110]}
   );
   gpc1_1 gpc7932 (
      {stage1_32[408]},
      {stage2_32[111]}
   );
   gpc1_1 gpc7933 (
      {stage1_32[409]},
      {stage2_32[112]}
   );
   gpc1_1 gpc7934 (
      {stage1_32[410]},
      {stage2_32[113]}
   );
   gpc1_1 gpc7935 (
      {stage1_32[411]},
      {stage2_32[114]}
   );
   gpc1_1 gpc7936 (
      {stage1_32[412]},
      {stage2_32[115]}
   );
   gpc1_1 gpc7937 (
      {stage1_32[413]},
      {stage2_32[116]}
   );
   gpc1_1 gpc7938 (
      {stage1_32[414]},
      {stage2_32[117]}
   );
   gpc1_1 gpc7939 (
      {stage1_34[242]},
      {stage2_34[102]}
   );
   gpc1_1 gpc7940 (
      {stage1_34[243]},
      {stage2_34[103]}
   );
   gpc1_1 gpc7941 (
      {stage1_34[244]},
      {stage2_34[104]}
   );
   gpc1_1 gpc7942 (
      {stage1_34[245]},
      {stage2_34[105]}
   );
   gpc1_1 gpc7943 (
      {stage1_34[246]},
      {stage2_34[106]}
   );
   gpc1_1 gpc7944 (
      {stage1_34[247]},
      {stage2_34[107]}
   );
   gpc1_1 gpc7945 (
      {stage1_34[248]},
      {stage2_34[108]}
   );
   gpc1_1 gpc7946 (
      {stage1_34[249]},
      {stage2_34[109]}
   );
   gpc1_1 gpc7947 (
      {stage1_34[250]},
      {stage2_34[110]}
   );
   gpc1_1 gpc7948 (
      {stage1_34[251]},
      {stage2_34[111]}
   );
   gpc1_1 gpc7949 (
      {stage1_34[252]},
      {stage2_34[112]}
   );
   gpc1_1 gpc7950 (
      {stage1_34[253]},
      {stage2_34[113]}
   );
   gpc1_1 gpc7951 (
      {stage1_34[254]},
      {stage2_34[114]}
   );
   gpc1_1 gpc7952 (
      {stage1_34[255]},
      {stage2_34[115]}
   );
   gpc1_1 gpc7953 (
      {stage1_34[256]},
      {stage2_34[116]}
   );
   gpc1_1 gpc7954 (
      {stage1_34[257]},
      {stage2_34[117]}
   );
   gpc1_1 gpc7955 (
      {stage1_34[258]},
      {stage2_34[118]}
   );
   gpc1_1 gpc7956 (
      {stage1_34[259]},
      {stage2_34[119]}
   );
   gpc1_1 gpc7957 (
      {stage1_34[260]},
      {stage2_34[120]}
   );
   gpc1_1 gpc7958 (
      {stage1_34[261]},
      {stage2_34[121]}
   );
   gpc1_1 gpc7959 (
      {stage1_34[262]},
      {stage2_34[122]}
   );
   gpc1_1 gpc7960 (
      {stage1_34[263]},
      {stage2_34[123]}
   );
   gpc1_1 gpc7961 (
      {stage1_34[264]},
      {stage2_34[124]}
   );
   gpc1_1 gpc7962 (
      {stage1_34[265]},
      {stage2_34[125]}
   );
   gpc1_1 gpc7963 (
      {stage1_34[266]},
      {stage2_34[126]}
   );
   gpc1_1 gpc7964 (
      {stage1_34[267]},
      {stage2_34[127]}
   );
   gpc1_1 gpc7965 (
      {stage1_35[173]},
      {stage2_35[100]}
   );
   gpc1_1 gpc7966 (
      {stage1_35[174]},
      {stage2_35[101]}
   );
   gpc1_1 gpc7967 (
      {stage1_35[175]},
      {stage2_35[102]}
   );
   gpc1_1 gpc7968 (
      {stage1_35[176]},
      {stage2_35[103]}
   );
   gpc1_1 gpc7969 (
      {stage1_35[177]},
      {stage2_35[104]}
   );
   gpc1_1 gpc7970 (
      {stage1_35[178]},
      {stage2_35[105]}
   );
   gpc1_1 gpc7971 (
      {stage1_35[179]},
      {stage2_35[106]}
   );
   gpc1_1 gpc7972 (
      {stage1_35[180]},
      {stage2_35[107]}
   );
   gpc1_1 gpc7973 (
      {stage1_35[181]},
      {stage2_35[108]}
   );
   gpc1_1 gpc7974 (
      {stage1_35[182]},
      {stage2_35[109]}
   );
   gpc1_1 gpc7975 (
      {stage1_35[183]},
      {stage2_35[110]}
   );
   gpc1_1 gpc7976 (
      {stage1_35[184]},
      {stage2_35[111]}
   );
   gpc1_1 gpc7977 (
      {stage1_35[185]},
      {stage2_35[112]}
   );
   gpc1_1 gpc7978 (
      {stage1_35[186]},
      {stage2_35[113]}
   );
   gpc1_1 gpc7979 (
      {stage1_35[187]},
      {stage2_35[114]}
   );
   gpc1_1 gpc7980 (
      {stage1_35[188]},
      {stage2_35[115]}
   );
   gpc1_1 gpc7981 (
      {stage1_35[189]},
      {stage2_35[116]}
   );
   gpc1_1 gpc7982 (
      {stage1_35[190]},
      {stage2_35[117]}
   );
   gpc1_1 gpc7983 (
      {stage1_37[297]},
      {stage2_37[108]}
   );
   gpc1_1 gpc7984 (
      {stage1_37[298]},
      {stage2_37[109]}
   );
   gpc1_1 gpc7985 (
      {stage1_37[299]},
      {stage2_37[110]}
   );
   gpc1_1 gpc7986 (
      {stage1_37[300]},
      {stage2_37[111]}
   );
   gpc1_1 gpc7987 (
      {stage1_37[301]},
      {stage2_37[112]}
   );
   gpc1_1 gpc7988 (
      {stage1_37[302]},
      {stage2_37[113]}
   );
   gpc1_1 gpc7989 (
      {stage1_39[194]},
      {stage2_39[105]}
   );
   gpc1_1 gpc7990 (
      {stage1_39[195]},
      {stage2_39[106]}
   );
   gpc1_1 gpc7991 (
      {stage1_39[196]},
      {stage2_39[107]}
   );
   gpc1_1 gpc7992 (
      {stage1_40[203]},
      {stage2_40[113]}
   );
   gpc1_1 gpc7993 (
      {stage1_40[204]},
      {stage2_40[114]}
   );
   gpc1_1 gpc7994 (
      {stage1_40[205]},
      {stage2_40[115]}
   );
   gpc1_1 gpc7995 (
      {stage1_40[206]},
      {stage2_40[116]}
   );
   gpc1_1 gpc7996 (
      {stage1_40[207]},
      {stage2_40[117]}
   );
   gpc1_1 gpc7997 (
      {stage1_40[208]},
      {stage2_40[118]}
   );
   gpc1_1 gpc7998 (
      {stage1_40[209]},
      {stage2_40[119]}
   );
   gpc1_1 gpc7999 (
      {stage1_40[210]},
      {stage2_40[120]}
   );
   gpc1_1 gpc8000 (
      {stage1_40[211]},
      {stage2_40[121]}
   );
   gpc1_1 gpc8001 (
      {stage1_40[212]},
      {stage2_40[122]}
   );
   gpc1_1 gpc8002 (
      {stage1_40[213]},
      {stage2_40[123]}
   );
   gpc1_1 gpc8003 (
      {stage1_40[214]},
      {stage2_40[124]}
   );
   gpc1_1 gpc8004 (
      {stage1_40[215]},
      {stage2_40[125]}
   );
   gpc1_1 gpc8005 (
      {stage1_40[216]},
      {stage2_40[126]}
   );
   gpc1_1 gpc8006 (
      {stage1_40[217]},
      {stage2_40[127]}
   );
   gpc1_1 gpc8007 (
      {stage1_40[218]},
      {stage2_40[128]}
   );
   gpc1_1 gpc8008 (
      {stage1_40[219]},
      {stage2_40[129]}
   );
   gpc1_1 gpc8009 (
      {stage1_40[220]},
      {stage2_40[130]}
   );
   gpc1_1 gpc8010 (
      {stage1_40[221]},
      {stage2_40[131]}
   );
   gpc1_1 gpc8011 (
      {stage1_40[222]},
      {stage2_40[132]}
   );
   gpc1_1 gpc8012 (
      {stage1_40[223]},
      {stage2_40[133]}
   );
   gpc1_1 gpc8013 (
      {stage1_40[224]},
      {stage2_40[134]}
   );
   gpc1_1 gpc8014 (
      {stage1_40[225]},
      {stage2_40[135]}
   );
   gpc1_1 gpc8015 (
      {stage1_40[226]},
      {stage2_40[136]}
   );
   gpc1_1 gpc8016 (
      {stage1_40[227]},
      {stage2_40[137]}
   );
   gpc1_1 gpc8017 (
      {stage1_40[228]},
      {stage2_40[138]}
   );
   gpc1_1 gpc8018 (
      {stage1_40[229]},
      {stage2_40[139]}
   );
   gpc1_1 gpc8019 (
      {stage1_41[252]},
      {stage2_41[98]}
   );
   gpc1_1 gpc8020 (
      {stage1_41[253]},
      {stage2_41[99]}
   );
   gpc1_1 gpc8021 (
      {stage1_41[254]},
      {stage2_41[100]}
   );
   gpc1_1 gpc8022 (
      {stage1_41[255]},
      {stage2_41[101]}
   );
   gpc1_1 gpc8023 (
      {stage1_41[256]},
      {stage2_41[102]}
   );
   gpc1_1 gpc8024 (
      {stage1_41[257]},
      {stage2_41[103]}
   );
   gpc1_1 gpc8025 (
      {stage1_41[258]},
      {stage2_41[104]}
   );
   gpc1_1 gpc8026 (
      {stage1_41[259]},
      {stage2_41[105]}
   );
   gpc1_1 gpc8027 (
      {stage1_41[260]},
      {stage2_41[106]}
   );
   gpc1_1 gpc8028 (
      {stage1_41[261]},
      {stage2_41[107]}
   );
   gpc1_1 gpc8029 (
      {stage1_41[262]},
      {stage2_41[108]}
   );
   gpc1_1 gpc8030 (
      {stage1_41[263]},
      {stage2_41[109]}
   );
   gpc1_1 gpc8031 (
      {stage1_41[264]},
      {stage2_41[110]}
   );
   gpc1_1 gpc8032 (
      {stage1_41[265]},
      {stage2_41[111]}
   );
   gpc1_1 gpc8033 (
      {stage1_41[266]},
      {stage2_41[112]}
   );
   gpc1_1 gpc8034 (
      {stage1_41[267]},
      {stage2_41[113]}
   );
   gpc1_1 gpc8035 (
      {stage1_41[268]},
      {stage2_41[114]}
   );
   gpc1_1 gpc8036 (
      {stage1_41[269]},
      {stage2_41[115]}
   );
   gpc1_1 gpc8037 (
      {stage1_41[270]},
      {stage2_41[116]}
   );
   gpc1_1 gpc8038 (
      {stage1_41[271]},
      {stage2_41[117]}
   );
   gpc1_1 gpc8039 (
      {stage1_41[272]},
      {stage2_41[118]}
   );
   gpc1_1 gpc8040 (
      {stage1_41[273]},
      {stage2_41[119]}
   );
   gpc1_1 gpc8041 (
      {stage1_41[274]},
      {stage2_41[120]}
   );
   gpc1_1 gpc8042 (
      {stage1_41[275]},
      {stage2_41[121]}
   );
   gpc1_1 gpc8043 (
      {stage1_41[276]},
      {stage2_41[122]}
   );
   gpc1_1 gpc8044 (
      {stage1_42[228]},
      {stage2_42[81]}
   );
   gpc1_1 gpc8045 (
      {stage1_43[218]},
      {stage2_43[85]}
   );
   gpc1_1 gpc8046 (
      {stage1_43[219]},
      {stage2_43[86]}
   );
   gpc1_1 gpc8047 (
      {stage1_43[220]},
      {stage2_43[87]}
   );
   gpc1_1 gpc8048 (
      {stage1_43[221]},
      {stage2_43[88]}
   );
   gpc1_1 gpc8049 (
      {stage1_43[222]},
      {stage2_43[89]}
   );
   gpc1_1 gpc8050 (
      {stage1_43[223]},
      {stage2_43[90]}
   );
   gpc1_1 gpc8051 (
      {stage1_43[224]},
      {stage2_43[91]}
   );
   gpc1_1 gpc8052 (
      {stage1_43[225]},
      {stage2_43[92]}
   );
   gpc1_1 gpc8053 (
      {stage1_43[226]},
      {stage2_43[93]}
   );
   gpc1_1 gpc8054 (
      {stage1_43[227]},
      {stage2_43[94]}
   );
   gpc1_1 gpc8055 (
      {stage1_43[228]},
      {stage2_43[95]}
   );
   gpc1_1 gpc8056 (
      {stage1_43[229]},
      {stage2_43[96]}
   );
   gpc1_1 gpc8057 (
      {stage1_43[230]},
      {stage2_43[97]}
   );
   gpc1_1 gpc8058 (
      {stage1_43[231]},
      {stage2_43[98]}
   );
   gpc1_1 gpc8059 (
      {stage1_43[232]},
      {stage2_43[99]}
   );
   gpc1_1 gpc8060 (
      {stage1_43[233]},
      {stage2_43[100]}
   );
   gpc1_1 gpc8061 (
      {stage1_43[234]},
      {stage2_43[101]}
   );
   gpc1_1 gpc8062 (
      {stage1_43[235]},
      {stage2_43[102]}
   );
   gpc1_1 gpc8063 (
      {stage1_43[236]},
      {stage2_43[103]}
   );
   gpc1_1 gpc8064 (
      {stage1_43[237]},
      {stage2_43[104]}
   );
   gpc1_1 gpc8065 (
      {stage1_43[238]},
      {stage2_43[105]}
   );
   gpc1_1 gpc8066 (
      {stage1_43[239]},
      {stage2_43[106]}
   );
   gpc1_1 gpc8067 (
      {stage1_43[240]},
      {stage2_43[107]}
   );
   gpc1_1 gpc8068 (
      {stage1_43[241]},
      {stage2_43[108]}
   );
   gpc1_1 gpc8069 (
      {stage1_43[242]},
      {stage2_43[109]}
   );
   gpc1_1 gpc8070 (
      {stage1_43[243]},
      {stage2_43[110]}
   );
   gpc1_1 gpc8071 (
      {stage1_44[244]},
      {stage2_44[113]}
   );
   gpc1_1 gpc8072 (
      {stage1_44[245]},
      {stage2_44[114]}
   );
   gpc1_1 gpc8073 (
      {stage1_44[246]},
      {stage2_44[115]}
   );
   gpc1_1 gpc8074 (
      {stage1_44[247]},
      {stage2_44[116]}
   );
   gpc1_1 gpc8075 (
      {stage1_44[248]},
      {stage2_44[117]}
   );
   gpc1_1 gpc8076 (
      {stage1_44[249]},
      {stage2_44[118]}
   );
   gpc1_1 gpc8077 (
      {stage1_44[250]},
      {stage2_44[119]}
   );
   gpc1_1 gpc8078 (
      {stage1_44[251]},
      {stage2_44[120]}
   );
   gpc1_1 gpc8079 (
      {stage1_44[252]},
      {stage2_44[121]}
   );
   gpc1_1 gpc8080 (
      {stage1_44[253]},
      {stage2_44[122]}
   );
   gpc1_1 gpc8081 (
      {stage1_44[254]},
      {stage2_44[123]}
   );
   gpc1_1 gpc8082 (
      {stage1_44[255]},
      {stage2_44[124]}
   );
   gpc1_1 gpc8083 (
      {stage1_44[256]},
      {stage2_44[125]}
   );
   gpc1_1 gpc8084 (
      {stage1_44[257]},
      {stage2_44[126]}
   );
   gpc1_1 gpc8085 (
      {stage1_44[258]},
      {stage2_44[127]}
   );
   gpc1_1 gpc8086 (
      {stage1_44[259]},
      {stage2_44[128]}
   );
   gpc1_1 gpc8087 (
      {stage1_44[260]},
      {stage2_44[129]}
   );
   gpc1_1 gpc8088 (
      {stage1_44[261]},
      {stage2_44[130]}
   );
   gpc1_1 gpc8089 (
      {stage1_44[262]},
      {stage2_44[131]}
   );
   gpc1_1 gpc8090 (
      {stage1_44[263]},
      {stage2_44[132]}
   );
   gpc1_1 gpc8091 (
      {stage1_44[264]},
      {stage2_44[133]}
   );
   gpc1_1 gpc8092 (
      {stage1_44[265]},
      {stage2_44[134]}
   );
   gpc1_1 gpc8093 (
      {stage1_44[266]},
      {stage2_44[135]}
   );
   gpc1_1 gpc8094 (
      {stage1_44[267]},
      {stage2_44[136]}
   );
   gpc1_1 gpc8095 (
      {stage1_44[268]},
      {stage2_44[137]}
   );
   gpc1_1 gpc8096 (
      {stage1_45[157]},
      {stage2_45[100]}
   );
   gpc1_1 gpc8097 (
      {stage1_45[158]},
      {stage2_45[101]}
   );
   gpc1_1 gpc8098 (
      {stage1_45[159]},
      {stage2_45[102]}
   );
   gpc1_1 gpc8099 (
      {stage1_45[160]},
      {stage2_45[103]}
   );
   gpc1_1 gpc8100 (
      {stage1_45[161]},
      {stage2_45[104]}
   );
   gpc1_1 gpc8101 (
      {stage1_45[162]},
      {stage2_45[105]}
   );
   gpc1_1 gpc8102 (
      {stage1_45[163]},
      {stage2_45[106]}
   );
   gpc1_1 gpc8103 (
      {stage1_45[164]},
      {stage2_45[107]}
   );
   gpc1_1 gpc8104 (
      {stage1_45[165]},
      {stage2_45[108]}
   );
   gpc1_1 gpc8105 (
      {stage1_45[166]},
      {stage2_45[109]}
   );
   gpc1_1 gpc8106 (
      {stage1_45[167]},
      {stage2_45[110]}
   );
   gpc1_1 gpc8107 (
      {stage1_45[168]},
      {stage2_45[111]}
   );
   gpc1_1 gpc8108 (
      {stage1_45[169]},
      {stage2_45[112]}
   );
   gpc1_1 gpc8109 (
      {stage1_45[170]},
      {stage2_45[113]}
   );
   gpc1_1 gpc8110 (
      {stage1_45[171]},
      {stage2_45[114]}
   );
   gpc1_1 gpc8111 (
      {stage1_45[172]},
      {stage2_45[115]}
   );
   gpc1_1 gpc8112 (
      {stage1_45[173]},
      {stage2_45[116]}
   );
   gpc1_1 gpc8113 (
      {stage1_45[174]},
      {stage2_45[117]}
   );
   gpc1_1 gpc8114 (
      {stage1_45[175]},
      {stage2_45[118]}
   );
   gpc1_1 gpc8115 (
      {stage1_45[176]},
      {stage2_45[119]}
   );
   gpc1_1 gpc8116 (
      {stage1_45[177]},
      {stage2_45[120]}
   );
   gpc1_1 gpc8117 (
      {stage1_45[178]},
      {stage2_45[121]}
   );
   gpc1_1 gpc8118 (
      {stage1_45[179]},
      {stage2_45[122]}
   );
   gpc1_1 gpc8119 (
      {stage1_45[180]},
      {stage2_45[123]}
   );
   gpc1_1 gpc8120 (
      {stage1_45[181]},
      {stage2_45[124]}
   );
   gpc1_1 gpc8121 (
      {stage1_45[182]},
      {stage2_45[125]}
   );
   gpc1_1 gpc8122 (
      {stage1_45[183]},
      {stage2_45[126]}
   );
   gpc1_1 gpc8123 (
      {stage1_45[184]},
      {stage2_45[127]}
   );
   gpc1_1 gpc8124 (
      {stage1_45[185]},
      {stage2_45[128]}
   );
   gpc1_1 gpc8125 (
      {stage1_45[186]},
      {stage2_45[129]}
   );
   gpc1_1 gpc8126 (
      {stage1_45[187]},
      {stage2_45[130]}
   );
   gpc1_1 gpc8127 (
      {stage1_45[188]},
      {stage2_45[131]}
   );
   gpc1_1 gpc8128 (
      {stage1_46[285]},
      {stage2_46[78]}
   );
   gpc1_1 gpc8129 (
      {stage1_46[286]},
      {stage2_46[79]}
   );
   gpc1_1 gpc8130 (
      {stage1_46[287]},
      {stage2_46[80]}
   );
   gpc1_1 gpc8131 (
      {stage1_46[288]},
      {stage2_46[81]}
   );
   gpc1_1 gpc8132 (
      {stage1_46[289]},
      {stage2_46[82]}
   );
   gpc1_1 gpc8133 (
      {stage1_46[290]},
      {stage2_46[83]}
   );
   gpc1_1 gpc8134 (
      {stage1_46[291]},
      {stage2_46[84]}
   );
   gpc1_1 gpc8135 (
      {stage1_46[292]},
      {stage2_46[85]}
   );
   gpc1_1 gpc8136 (
      {stage1_46[293]},
      {stage2_46[86]}
   );
   gpc1_1 gpc8137 (
      {stage1_46[294]},
      {stage2_46[87]}
   );
   gpc1_1 gpc8138 (
      {stage1_46[295]},
      {stage2_46[88]}
   );
   gpc1_1 gpc8139 (
      {stage1_46[296]},
      {stage2_46[89]}
   );
   gpc1_1 gpc8140 (
      {stage1_46[297]},
      {stage2_46[90]}
   );
   gpc1_1 gpc8141 (
      {stage1_46[298]},
      {stage2_46[91]}
   );
   gpc1_1 gpc8142 (
      {stage1_46[299]},
      {stage2_46[92]}
   );
   gpc1_1 gpc8143 (
      {stage1_47[270]},
      {stage2_47[100]}
   );
   gpc1_1 gpc8144 (
      {stage1_47[271]},
      {stage2_47[101]}
   );
   gpc1_1 gpc8145 (
      {stage1_47[272]},
      {stage2_47[102]}
   );
   gpc1_1 gpc8146 (
      {stage1_47[273]},
      {stage2_47[103]}
   );
   gpc1_1 gpc8147 (
      {stage1_47[274]},
      {stage2_47[104]}
   );
   gpc1_1 gpc8148 (
      {stage1_47[275]},
      {stage2_47[105]}
   );
   gpc1_1 gpc8149 (
      {stage1_47[276]},
      {stage2_47[106]}
   );
   gpc1_1 gpc8150 (
      {stage1_47[277]},
      {stage2_47[107]}
   );
   gpc1_1 gpc8151 (
      {stage1_48[166]},
      {stage2_48[109]}
   );
   gpc1_1 gpc8152 (
      {stage1_48[167]},
      {stage2_48[110]}
   );
   gpc1_1 gpc8153 (
      {stage1_48[168]},
      {stage2_48[111]}
   );
   gpc1_1 gpc8154 (
      {stage1_48[169]},
      {stage2_48[112]}
   );
   gpc1_1 gpc8155 (
      {stage1_48[170]},
      {stage2_48[113]}
   );
   gpc1_1 gpc8156 (
      {stage1_48[171]},
      {stage2_48[114]}
   );
   gpc1_1 gpc8157 (
      {stage1_48[172]},
      {stage2_48[115]}
   );
   gpc1_1 gpc8158 (
      {stage1_48[173]},
      {stage2_48[116]}
   );
   gpc1_1 gpc8159 (
      {stage1_48[174]},
      {stage2_48[117]}
   );
   gpc1_1 gpc8160 (
      {stage1_48[175]},
      {stage2_48[118]}
   );
   gpc1_1 gpc8161 (
      {stage1_48[176]},
      {stage2_48[119]}
   );
   gpc1_1 gpc8162 (
      {stage1_48[177]},
      {stage2_48[120]}
   );
   gpc1_1 gpc8163 (
      {stage1_48[178]},
      {stage2_48[121]}
   );
   gpc1_1 gpc8164 (
      {stage1_48[179]},
      {stage2_48[122]}
   );
   gpc1_1 gpc8165 (
      {stage1_48[180]},
      {stage2_48[123]}
   );
   gpc1_1 gpc8166 (
      {stage1_48[181]},
      {stage2_48[124]}
   );
   gpc1_1 gpc8167 (
      {stage1_48[182]},
      {stage2_48[125]}
   );
   gpc1_1 gpc8168 (
      {stage1_48[183]},
      {stage2_48[126]}
   );
   gpc1_1 gpc8169 (
      {stage1_48[184]},
      {stage2_48[127]}
   );
   gpc1_1 gpc8170 (
      {stage1_48[185]},
      {stage2_48[128]}
   );
   gpc1_1 gpc8171 (
      {stage1_48[186]},
      {stage2_48[129]}
   );
   gpc1_1 gpc8172 (
      {stage1_48[187]},
      {stage2_48[130]}
   );
   gpc1_1 gpc8173 (
      {stage1_48[188]},
      {stage2_48[131]}
   );
   gpc1_1 gpc8174 (
      {stage1_48[189]},
      {stage2_48[132]}
   );
   gpc1_1 gpc8175 (
      {stage1_48[190]},
      {stage2_48[133]}
   );
   gpc1_1 gpc8176 (
      {stage1_48[191]},
      {stage2_48[134]}
   );
   gpc1_1 gpc8177 (
      {stage1_48[192]},
      {stage2_48[135]}
   );
   gpc1_1 gpc8178 (
      {stage1_48[193]},
      {stage2_48[136]}
   );
   gpc1_1 gpc8179 (
      {stage1_48[194]},
      {stage2_48[137]}
   );
   gpc1_1 gpc8180 (
      {stage1_48[195]},
      {stage2_48[138]}
   );
   gpc1_1 gpc8181 (
      {stage1_48[196]},
      {stage2_48[139]}
   );
   gpc1_1 gpc8182 (
      {stage1_48[197]},
      {stage2_48[140]}
   );
   gpc1_1 gpc8183 (
      {stage1_48[198]},
      {stage2_48[141]}
   );
   gpc1_1 gpc8184 (
      {stage1_48[199]},
      {stage2_48[142]}
   );
   gpc1_1 gpc8185 (
      {stage1_48[200]},
      {stage2_48[143]}
   );
   gpc1_1 gpc8186 (
      {stage1_48[201]},
      {stage2_48[144]}
   );
   gpc1_1 gpc8187 (
      {stage1_48[202]},
      {stage2_48[145]}
   );
   gpc1_1 gpc8188 (
      {stage1_48[203]},
      {stage2_48[146]}
   );
   gpc1_1 gpc8189 (
      {stage1_48[204]},
      {stage2_48[147]}
   );
   gpc1_1 gpc8190 (
      {stage1_48[205]},
      {stage2_48[148]}
   );
   gpc1_1 gpc8191 (
      {stage1_48[206]},
      {stage2_48[149]}
   );
   gpc1_1 gpc8192 (
      {stage1_48[207]},
      {stage2_48[150]}
   );
   gpc1_1 gpc8193 (
      {stage1_48[208]},
      {stage2_48[151]}
   );
   gpc1_1 gpc8194 (
      {stage1_48[209]},
      {stage2_48[152]}
   );
   gpc1_1 gpc8195 (
      {stage1_48[210]},
      {stage2_48[153]}
   );
   gpc1_1 gpc8196 (
      {stage1_49[203]},
      {stage2_49[77]}
   );
   gpc1_1 gpc8197 (
      {stage1_49[204]},
      {stage2_49[78]}
   );
   gpc1_1 gpc8198 (
      {stage1_49[205]},
      {stage2_49[79]}
   );
   gpc1_1 gpc8199 (
      {stage1_49[206]},
      {stage2_49[80]}
   );
   gpc1_1 gpc8200 (
      {stage1_49[207]},
      {stage2_49[81]}
   );
   gpc1_1 gpc8201 (
      {stage1_49[208]},
      {stage2_49[82]}
   );
   gpc1_1 gpc8202 (
      {stage1_49[209]},
      {stage2_49[83]}
   );
   gpc1_1 gpc8203 (
      {stage1_49[210]},
      {stage2_49[84]}
   );
   gpc1_1 gpc8204 (
      {stage1_49[211]},
      {stage2_49[85]}
   );
   gpc1_1 gpc8205 (
      {stage1_49[212]},
      {stage2_49[86]}
   );
   gpc1_1 gpc8206 (
      {stage1_49[213]},
      {stage2_49[87]}
   );
   gpc1_1 gpc8207 (
      {stage1_49[214]},
      {stage2_49[88]}
   );
   gpc1_1 gpc8208 (
      {stage1_49[215]},
      {stage2_49[89]}
   );
   gpc1_1 gpc8209 (
      {stage1_49[216]},
      {stage2_49[90]}
   );
   gpc1_1 gpc8210 (
      {stage1_49[217]},
      {stage2_49[91]}
   );
   gpc1_1 gpc8211 (
      {stage1_49[218]},
      {stage2_49[92]}
   );
   gpc1_1 gpc8212 (
      {stage1_49[219]},
      {stage2_49[93]}
   );
   gpc1_1 gpc8213 (
      {stage1_49[220]},
      {stage2_49[94]}
   );
   gpc1_1 gpc8214 (
      {stage1_49[221]},
      {stage2_49[95]}
   );
   gpc1_1 gpc8215 (
      {stage1_49[222]},
      {stage2_49[96]}
   );
   gpc1_1 gpc8216 (
      {stage1_49[223]},
      {stage2_49[97]}
   );
   gpc1_1 gpc8217 (
      {stage1_49[224]},
      {stage2_49[98]}
   );
   gpc1_1 gpc8218 (
      {stage1_49[225]},
      {stage2_49[99]}
   );
   gpc1_1 gpc8219 (
      {stage1_49[226]},
      {stage2_49[100]}
   );
   gpc1_1 gpc8220 (
      {stage1_49[227]},
      {stage2_49[101]}
   );
   gpc1_1 gpc8221 (
      {stage1_49[228]},
      {stage2_49[102]}
   );
   gpc1_1 gpc8222 (
      {stage1_49[229]},
      {stage2_49[103]}
   );
   gpc1_1 gpc8223 (
      {stage1_49[230]},
      {stage2_49[104]}
   );
   gpc1_1 gpc8224 (
      {stage1_49[231]},
      {stage2_49[105]}
   );
   gpc1_1 gpc8225 (
      {stage1_49[232]},
      {stage2_49[106]}
   );
   gpc1_1 gpc8226 (
      {stage1_49[233]},
      {stage2_49[107]}
   );
   gpc1_1 gpc8227 (
      {stage1_49[234]},
      {stage2_49[108]}
   );
   gpc1_1 gpc8228 (
      {stage1_49[235]},
      {stage2_49[109]}
   );
   gpc1_1 gpc8229 (
      {stage1_49[236]},
      {stage2_49[110]}
   );
   gpc1_1 gpc8230 (
      {stage1_49[237]},
      {stage2_49[111]}
   );
   gpc1_1 gpc8231 (
      {stage1_49[238]},
      {stage2_49[112]}
   );
   gpc1_1 gpc8232 (
      {stage1_49[239]},
      {stage2_49[113]}
   );
   gpc1_1 gpc8233 (
      {stage1_49[240]},
      {stage2_49[114]}
   );
   gpc1_1 gpc8234 (
      {stage1_49[241]},
      {stage2_49[115]}
   );
   gpc1_1 gpc8235 (
      {stage1_50[134]},
      {stage2_50[70]}
   );
   gpc1_1 gpc8236 (
      {stage1_50[135]},
      {stage2_50[71]}
   );
   gpc1_1 gpc8237 (
      {stage1_50[136]},
      {stage2_50[72]}
   );
   gpc1_1 gpc8238 (
      {stage1_50[137]},
      {stage2_50[73]}
   );
   gpc1_1 gpc8239 (
      {stage1_50[138]},
      {stage2_50[74]}
   );
   gpc1_1 gpc8240 (
      {stage1_50[139]},
      {stage2_50[75]}
   );
   gpc1_1 gpc8241 (
      {stage1_50[140]},
      {stage2_50[76]}
   );
   gpc1_1 gpc8242 (
      {stage1_50[141]},
      {stage2_50[77]}
   );
   gpc1_1 gpc8243 (
      {stage1_50[142]},
      {stage2_50[78]}
   );
   gpc1_1 gpc8244 (
      {stage1_50[143]},
      {stage2_50[79]}
   );
   gpc1_1 gpc8245 (
      {stage1_50[144]},
      {stage2_50[80]}
   );
   gpc1_1 gpc8246 (
      {stage1_50[145]},
      {stage2_50[81]}
   );
   gpc1_1 gpc8247 (
      {stage1_50[146]},
      {stage2_50[82]}
   );
   gpc1_1 gpc8248 (
      {stage1_50[147]},
      {stage2_50[83]}
   );
   gpc1_1 gpc8249 (
      {stage1_50[148]},
      {stage2_50[84]}
   );
   gpc1_1 gpc8250 (
      {stage1_50[149]},
      {stage2_50[85]}
   );
   gpc1_1 gpc8251 (
      {stage1_50[150]},
      {stage2_50[86]}
   );
   gpc1_1 gpc8252 (
      {stage1_50[151]},
      {stage2_50[87]}
   );
   gpc1_1 gpc8253 (
      {stage1_50[152]},
      {stage2_50[88]}
   );
   gpc1_1 gpc8254 (
      {stage1_50[153]},
      {stage2_50[89]}
   );
   gpc1_1 gpc8255 (
      {stage1_50[154]},
      {stage2_50[90]}
   );
   gpc1_1 gpc8256 (
      {stage1_50[155]},
      {stage2_50[91]}
   );
   gpc1_1 gpc8257 (
      {stage1_50[156]},
      {stage2_50[92]}
   );
   gpc1_1 gpc8258 (
      {stage1_50[157]},
      {stage2_50[93]}
   );
   gpc1_1 gpc8259 (
      {stage1_50[158]},
      {stage2_50[94]}
   );
   gpc1_1 gpc8260 (
      {stage1_50[159]},
      {stage2_50[95]}
   );
   gpc1_1 gpc8261 (
      {stage1_50[160]},
      {stage2_50[96]}
   );
   gpc1_1 gpc8262 (
      {stage1_50[161]},
      {stage2_50[97]}
   );
   gpc1_1 gpc8263 (
      {stage1_50[162]},
      {stage2_50[98]}
   );
   gpc1_1 gpc8264 (
      {stage1_50[163]},
      {stage2_50[99]}
   );
   gpc1_1 gpc8265 (
      {stage1_50[164]},
      {stage2_50[100]}
   );
   gpc1_1 gpc8266 (
      {stage1_50[165]},
      {stage2_50[101]}
   );
   gpc1_1 gpc8267 (
      {stage1_50[166]},
      {stage2_50[102]}
   );
   gpc1_1 gpc8268 (
      {stage1_50[167]},
      {stage2_50[103]}
   );
   gpc1_1 gpc8269 (
      {stage1_50[168]},
      {stage2_50[104]}
   );
   gpc1_1 gpc8270 (
      {stage1_50[169]},
      {stage2_50[105]}
   );
   gpc1_1 gpc8271 (
      {stage1_50[170]},
      {stage2_50[106]}
   );
   gpc1_1 gpc8272 (
      {stage1_50[171]},
      {stage2_50[107]}
   );
   gpc1_1 gpc8273 (
      {stage1_50[172]},
      {stage2_50[108]}
   );
   gpc1_1 gpc8274 (
      {stage1_50[173]},
      {stage2_50[109]}
   );
   gpc1_1 gpc8275 (
      {stage1_50[174]},
      {stage2_50[110]}
   );
   gpc1_1 gpc8276 (
      {stage1_50[175]},
      {stage2_50[111]}
   );
   gpc1_1 gpc8277 (
      {stage1_50[176]},
      {stage2_50[112]}
   );
   gpc1_1 gpc8278 (
      {stage1_50[177]},
      {stage2_50[113]}
   );
   gpc1_1 gpc8279 (
      {stage1_50[178]},
      {stage2_50[114]}
   );
   gpc1_1 gpc8280 (
      {stage1_50[179]},
      {stage2_50[115]}
   );
   gpc1_1 gpc8281 (
      {stage1_50[180]},
      {stage2_50[116]}
   );
   gpc1_1 gpc8282 (
      {stage1_50[181]},
      {stage2_50[117]}
   );
   gpc1_1 gpc8283 (
      {stage1_50[182]},
      {stage2_50[118]}
   );
   gpc1_1 gpc8284 (
      {stage1_50[183]},
      {stage2_50[119]}
   );
   gpc1_1 gpc8285 (
      {stage1_50[184]},
      {stage2_50[120]}
   );
   gpc1_1 gpc8286 (
      {stage1_50[185]},
      {stage2_50[121]}
   );
   gpc1_1 gpc8287 (
      {stage1_50[186]},
      {stage2_50[122]}
   );
   gpc1_1 gpc8288 (
      {stage1_50[187]},
      {stage2_50[123]}
   );
   gpc1_1 gpc8289 (
      {stage1_50[188]},
      {stage2_50[124]}
   );
   gpc1_1 gpc8290 (
      {stage1_50[189]},
      {stage2_50[125]}
   );
   gpc1_1 gpc8291 (
      {stage1_50[190]},
      {stage2_50[126]}
   );
   gpc1_1 gpc8292 (
      {stage1_50[191]},
      {stage2_50[127]}
   );
   gpc1_1 gpc8293 (
      {stage1_50[192]},
      {stage2_50[128]}
   );
   gpc1_1 gpc8294 (
      {stage1_50[193]},
      {stage2_50[129]}
   );
   gpc1_1 gpc8295 (
      {stage1_50[194]},
      {stage2_50[130]}
   );
   gpc1_1 gpc8296 (
      {stage1_50[195]},
      {stage2_50[131]}
   );
   gpc1_1 gpc8297 (
      {stage1_50[196]},
      {stage2_50[132]}
   );
   gpc1_1 gpc8298 (
      {stage1_50[197]},
      {stage2_50[133]}
   );
   gpc1_1 gpc8299 (
      {stage1_50[198]},
      {stage2_50[134]}
   );
   gpc1_1 gpc8300 (
      {stage1_50[199]},
      {stage2_50[135]}
   );
   gpc1_1 gpc8301 (
      {stage1_50[200]},
      {stage2_50[136]}
   );
   gpc1_1 gpc8302 (
      {stage1_50[201]},
      {stage2_50[137]}
   );
   gpc1_1 gpc8303 (
      {stage1_50[202]},
      {stage2_50[138]}
   );
   gpc1_1 gpc8304 (
      {stage1_50[203]},
      {stage2_50[139]}
   );
   gpc1_1 gpc8305 (
      {stage1_50[204]},
      {stage2_50[140]}
   );
   gpc1_1 gpc8306 (
      {stage1_50[205]},
      {stage2_50[141]}
   );
   gpc1_1 gpc8307 (
      {stage1_50[206]},
      {stage2_50[142]}
   );
   gpc1_1 gpc8308 (
      {stage1_50[207]},
      {stage2_50[143]}
   );
   gpc1_1 gpc8309 (
      {stage1_50[208]},
      {stage2_50[144]}
   );
   gpc1_1 gpc8310 (
      {stage1_50[209]},
      {stage2_50[145]}
   );
   gpc1_1 gpc8311 (
      {stage1_50[210]},
      {stage2_50[146]}
   );
   gpc1_1 gpc8312 (
      {stage1_50[211]},
      {stage2_50[147]}
   );
   gpc1_1 gpc8313 (
      {stage1_50[212]},
      {stage2_50[148]}
   );
   gpc1_1 gpc8314 (
      {stage1_50[213]},
      {stage2_50[149]}
   );
   gpc1_1 gpc8315 (
      {stage1_50[214]},
      {stage2_50[150]}
   );
   gpc1_1 gpc8316 (
      {stage1_50[215]},
      {stage2_50[151]}
   );
   gpc1_1 gpc8317 (
      {stage1_50[216]},
      {stage2_50[152]}
   );
   gpc1_1 gpc8318 (
      {stage1_51[224]},
      {stage2_51[85]}
   );
   gpc1_1 gpc8319 (
      {stage1_51[225]},
      {stage2_51[86]}
   );
   gpc1_1 gpc8320 (
      {stage1_51[226]},
      {stage2_51[87]}
   );
   gpc1_1 gpc8321 (
      {stage1_52[269]},
      {stage2_52[93]}
   );
   gpc1_1 gpc8322 (
      {stage1_52[270]},
      {stage2_52[94]}
   );
   gpc1_1 gpc8323 (
      {stage1_52[271]},
      {stage2_52[95]}
   );
   gpc1_1 gpc8324 (
      {stage1_52[272]},
      {stage2_52[96]}
   );
   gpc1_1 gpc8325 (
      {stage1_52[273]},
      {stage2_52[97]}
   );
   gpc1_1 gpc8326 (
      {stage1_52[274]},
      {stage2_52[98]}
   );
   gpc1_1 gpc8327 (
      {stage1_52[275]},
      {stage2_52[99]}
   );
   gpc1_1 gpc8328 (
      {stage1_52[276]},
      {stage2_52[100]}
   );
   gpc1_1 gpc8329 (
      {stage1_52[277]},
      {stage2_52[101]}
   );
   gpc1_1 gpc8330 (
      {stage1_52[278]},
      {stage2_52[102]}
   );
   gpc1_1 gpc8331 (
      {stage1_52[279]},
      {stage2_52[103]}
   );
   gpc1_1 gpc8332 (
      {stage1_52[280]},
      {stage2_52[104]}
   );
   gpc1_1 gpc8333 (
      {stage1_52[281]},
      {stage2_52[105]}
   );
   gpc1_1 gpc8334 (
      {stage1_52[282]},
      {stage2_52[106]}
   );
   gpc1_1 gpc8335 (
      {stage1_52[283]},
      {stage2_52[107]}
   );
   gpc1_1 gpc8336 (
      {stage1_52[284]},
      {stage2_52[108]}
   );
   gpc1_1 gpc8337 (
      {stage1_52[285]},
      {stage2_52[109]}
   );
   gpc1_1 gpc8338 (
      {stage1_52[286]},
      {stage2_52[110]}
   );
   gpc1_1 gpc8339 (
      {stage1_52[287]},
      {stage2_52[111]}
   );
   gpc1_1 gpc8340 (
      {stage1_52[288]},
      {stage2_52[112]}
   );
   gpc1_1 gpc8341 (
      {stage1_52[289]},
      {stage2_52[113]}
   );
   gpc1_1 gpc8342 (
      {stage1_52[290]},
      {stage2_52[114]}
   );
   gpc1_1 gpc8343 (
      {stage1_52[291]},
      {stage2_52[115]}
   );
   gpc1_1 gpc8344 (
      {stage1_52[292]},
      {stage2_52[116]}
   );
   gpc1_1 gpc8345 (
      {stage1_52[293]},
      {stage2_52[117]}
   );
   gpc1_1 gpc8346 (
      {stage1_52[294]},
      {stage2_52[118]}
   );
   gpc1_1 gpc8347 (
      {stage1_52[295]},
      {stage2_52[119]}
   );
   gpc1_1 gpc8348 (
      {stage1_52[296]},
      {stage2_52[120]}
   );
   gpc1_1 gpc8349 (
      {stage1_52[297]},
      {stage2_52[121]}
   );
   gpc1_1 gpc8350 (
      {stage1_52[298]},
      {stage2_52[122]}
   );
   gpc1_1 gpc8351 (
      {stage1_52[299]},
      {stage2_52[123]}
   );
   gpc1_1 gpc8352 (
      {stage1_52[300]},
      {stage2_52[124]}
   );
   gpc1_1 gpc8353 (
      {stage1_52[301]},
      {stage2_52[125]}
   );
   gpc1_1 gpc8354 (
      {stage1_52[302]},
      {stage2_52[126]}
   );
   gpc1_1 gpc8355 (
      {stage1_52[303]},
      {stage2_52[127]}
   );
   gpc1_1 gpc8356 (
      {stage1_53[173]},
      {stage2_53[83]}
   );
   gpc1_1 gpc8357 (
      {stage1_53[174]},
      {stage2_53[84]}
   );
   gpc1_1 gpc8358 (
      {stage1_53[175]},
      {stage2_53[85]}
   );
   gpc1_1 gpc8359 (
      {stage1_53[176]},
      {stage2_53[86]}
   );
   gpc1_1 gpc8360 (
      {stage1_53[177]},
      {stage2_53[87]}
   );
   gpc1_1 gpc8361 (
      {stage1_53[178]},
      {stage2_53[88]}
   );
   gpc1_1 gpc8362 (
      {stage1_53[179]},
      {stage2_53[89]}
   );
   gpc1_1 gpc8363 (
      {stage1_53[180]},
      {stage2_53[90]}
   );
   gpc1_1 gpc8364 (
      {stage1_53[181]},
      {stage2_53[91]}
   );
   gpc1_1 gpc8365 (
      {stage1_53[182]},
      {stage2_53[92]}
   );
   gpc1_1 gpc8366 (
      {stage1_53[183]},
      {stage2_53[93]}
   );
   gpc1_1 gpc8367 (
      {stage1_53[184]},
      {stage2_53[94]}
   );
   gpc1_1 gpc8368 (
      {stage1_53[185]},
      {stage2_53[95]}
   );
   gpc1_1 gpc8369 (
      {stage1_53[186]},
      {stage2_53[96]}
   );
   gpc1_1 gpc8370 (
      {stage1_54[216]},
      {stage2_54[77]}
   );
   gpc1_1 gpc8371 (
      {stage1_54[217]},
      {stage2_54[78]}
   );
   gpc1_1 gpc8372 (
      {stage1_54[218]},
      {stage2_54[79]}
   );
   gpc1_1 gpc8373 (
      {stage1_54[219]},
      {stage2_54[80]}
   );
   gpc1_1 gpc8374 (
      {stage1_54[220]},
      {stage2_54[81]}
   );
   gpc1_1 gpc8375 (
      {stage1_54[221]},
      {stage2_54[82]}
   );
   gpc1_1 gpc8376 (
      {stage1_54[222]},
      {stage2_54[83]}
   );
   gpc1_1 gpc8377 (
      {stage1_54[223]},
      {stage2_54[84]}
   );
   gpc1_1 gpc8378 (
      {stage1_54[224]},
      {stage2_54[85]}
   );
   gpc1_1 gpc8379 (
      {stage1_54[225]},
      {stage2_54[86]}
   );
   gpc1_1 gpc8380 (
      {stage1_54[226]},
      {stage2_54[87]}
   );
   gpc1_1 gpc8381 (
      {stage1_54[227]},
      {stage2_54[88]}
   );
   gpc1_1 gpc8382 (
      {stage1_54[228]},
      {stage2_54[89]}
   );
   gpc1_1 gpc8383 (
      {stage1_54[229]},
      {stage2_54[90]}
   );
   gpc1_1 gpc8384 (
      {stage1_54[230]},
      {stage2_54[91]}
   );
   gpc1_1 gpc8385 (
      {stage1_54[231]},
      {stage2_54[92]}
   );
   gpc1_1 gpc8386 (
      {stage1_54[232]},
      {stage2_54[93]}
   );
   gpc1_1 gpc8387 (
      {stage1_54[233]},
      {stage2_54[94]}
   );
   gpc1_1 gpc8388 (
      {stage1_54[234]},
      {stage2_54[95]}
   );
   gpc1_1 gpc8389 (
      {stage1_54[235]},
      {stage2_54[96]}
   );
   gpc1_1 gpc8390 (
      {stage1_54[236]},
      {stage2_54[97]}
   );
   gpc1_1 gpc8391 (
      {stage1_54[237]},
      {stage2_54[98]}
   );
   gpc1_1 gpc8392 (
      {stage1_54[238]},
      {stage2_54[99]}
   );
   gpc1_1 gpc8393 (
      {stage1_54[239]},
      {stage2_54[100]}
   );
   gpc1_1 gpc8394 (
      {stage1_54[240]},
      {stage2_54[101]}
   );
   gpc1_1 gpc8395 (
      {stage1_54[241]},
      {stage2_54[102]}
   );
   gpc1_1 gpc8396 (
      {stage1_54[242]},
      {stage2_54[103]}
   );
   gpc1_1 gpc8397 (
      {stage1_54[243]},
      {stage2_54[104]}
   );
   gpc1_1 gpc8398 (
      {stage1_54[244]},
      {stage2_54[105]}
   );
   gpc1_1 gpc8399 (
      {stage1_54[245]},
      {stage2_54[106]}
   );
   gpc1_1 gpc8400 (
      {stage1_54[246]},
      {stage2_54[107]}
   );
   gpc1_1 gpc8401 (
      {stage1_54[247]},
      {stage2_54[108]}
   );
   gpc1_1 gpc8402 (
      {stage1_54[248]},
      {stage2_54[109]}
   );
   gpc1_1 gpc8403 (
      {stage1_54[249]},
      {stage2_54[110]}
   );
   gpc1_1 gpc8404 (
      {stage1_54[250]},
      {stage2_54[111]}
   );
   gpc1_1 gpc8405 (
      {stage1_54[251]},
      {stage2_54[112]}
   );
   gpc1_1 gpc8406 (
      {stage1_54[252]},
      {stage2_54[113]}
   );
   gpc1_1 gpc8407 (
      {stage1_54[253]},
      {stage2_54[114]}
   );
   gpc1_1 gpc8408 (
      {stage1_54[254]},
      {stage2_54[115]}
   );
   gpc1_1 gpc8409 (
      {stage1_54[255]},
      {stage2_54[116]}
   );
   gpc1_1 gpc8410 (
      {stage1_54[256]},
      {stage2_54[117]}
   );
   gpc1_1 gpc8411 (
      {stage1_54[257]},
      {stage2_54[118]}
   );
   gpc1_1 gpc8412 (
      {stage1_54[258]},
      {stage2_54[119]}
   );
   gpc1_1 gpc8413 (
      {stage1_54[259]},
      {stage2_54[120]}
   );
   gpc1_1 gpc8414 (
      {stage1_54[260]},
      {stage2_54[121]}
   );
   gpc1_1 gpc8415 (
      {stage1_54[261]},
      {stage2_54[122]}
   );
   gpc1_1 gpc8416 (
      {stage1_54[262]},
      {stage2_54[123]}
   );
   gpc1_1 gpc8417 (
      {stage1_55[219]},
      {stage2_55[104]}
   );
   gpc1_1 gpc8418 (
      {stage1_55[220]},
      {stage2_55[105]}
   );
   gpc1_1 gpc8419 (
      {stage1_55[221]},
      {stage2_55[106]}
   );
   gpc1_1 gpc8420 (
      {stage1_55[222]},
      {stage2_55[107]}
   );
   gpc1_1 gpc8421 (
      {stage1_55[223]},
      {stage2_55[108]}
   );
   gpc1_1 gpc8422 (
      {stage1_55[224]},
      {stage2_55[109]}
   );
   gpc1_1 gpc8423 (
      {stage1_55[225]},
      {stage2_55[110]}
   );
   gpc1_1 gpc8424 (
      {stage1_56[225]},
      {stage2_56[100]}
   );
   gpc1_1 gpc8425 (
      {stage1_56[226]},
      {stage2_56[101]}
   );
   gpc1_1 gpc8426 (
      {stage1_56[227]},
      {stage2_56[102]}
   );
   gpc1_1 gpc8427 (
      {stage1_56[228]},
      {stage2_56[103]}
   );
   gpc1_1 gpc8428 (
      {stage1_56[229]},
      {stage2_56[104]}
   );
   gpc1_1 gpc8429 (
      {stage1_56[230]},
      {stage2_56[105]}
   );
   gpc1_1 gpc8430 (
      {stage1_56[231]},
      {stage2_56[106]}
   );
   gpc1_1 gpc8431 (
      {stage1_56[232]},
      {stage2_56[107]}
   );
   gpc1_1 gpc8432 (
      {stage1_56[233]},
      {stage2_56[108]}
   );
   gpc1_1 gpc8433 (
      {stage1_56[234]},
      {stage2_56[109]}
   );
   gpc1_1 gpc8434 (
      {stage1_56[235]},
      {stage2_56[110]}
   );
   gpc1_1 gpc8435 (
      {stage1_56[236]},
      {stage2_56[111]}
   );
   gpc1_1 gpc8436 (
      {stage1_56[237]},
      {stage2_56[112]}
   );
   gpc1_1 gpc8437 (
      {stage1_56[238]},
      {stage2_56[113]}
   );
   gpc1_1 gpc8438 (
      {stage1_56[239]},
      {stage2_56[114]}
   );
   gpc1_1 gpc8439 (
      {stage1_56[240]},
      {stage2_56[115]}
   );
   gpc1_1 gpc8440 (
      {stage1_56[241]},
      {stage2_56[116]}
   );
   gpc1_1 gpc8441 (
      {stage1_56[242]},
      {stage2_56[117]}
   );
   gpc1_1 gpc8442 (
      {stage1_56[243]},
      {stage2_56[118]}
   );
   gpc1_1 gpc8443 (
      {stage1_56[244]},
      {stage2_56[119]}
   );
   gpc1_1 gpc8444 (
      {stage1_56[245]},
      {stage2_56[120]}
   );
   gpc1_1 gpc8445 (
      {stage1_56[246]},
      {stage2_56[121]}
   );
   gpc1_1 gpc8446 (
      {stage1_56[247]},
      {stage2_56[122]}
   );
   gpc1_1 gpc8447 (
      {stage1_56[248]},
      {stage2_56[123]}
   );
   gpc1_1 gpc8448 (
      {stage1_56[249]},
      {stage2_56[124]}
   );
   gpc1_1 gpc8449 (
      {stage1_56[250]},
      {stage2_56[125]}
   );
   gpc1_1 gpc8450 (
      {stage1_56[251]},
      {stage2_56[126]}
   );
   gpc1_1 gpc8451 (
      {stage1_56[252]},
      {stage2_56[127]}
   );
   gpc1_1 gpc8452 (
      {stage1_56[253]},
      {stage2_56[128]}
   );
   gpc1_1 gpc8453 (
      {stage1_56[254]},
      {stage2_56[129]}
   );
   gpc1_1 gpc8454 (
      {stage1_56[255]},
      {stage2_56[130]}
   );
   gpc1_1 gpc8455 (
      {stage1_56[256]},
      {stage2_56[131]}
   );
   gpc1_1 gpc8456 (
      {stage1_59[268]},
      {stage2_59[114]}
   );
   gpc1_1 gpc8457 (
      {stage1_59[269]},
      {stage2_59[115]}
   );
   gpc1_1 gpc8458 (
      {stage1_59[270]},
      {stage2_59[116]}
   );
   gpc1_1 gpc8459 (
      {stage1_59[271]},
      {stage2_59[117]}
   );
   gpc1_1 gpc8460 (
      {stage1_59[272]},
      {stage2_59[118]}
   );
   gpc1_1 gpc8461 (
      {stage1_59[273]},
      {stage2_59[119]}
   );
   gpc1_1 gpc8462 (
      {stage1_59[274]},
      {stage2_59[120]}
   );
   gpc1_1 gpc8463 (
      {stage1_59[275]},
      {stage2_59[121]}
   );
   gpc1_1 gpc8464 (
      {stage1_59[276]},
      {stage2_59[122]}
   );
   gpc1_1 gpc8465 (
      {stage1_59[277]},
      {stage2_59[123]}
   );
   gpc1_1 gpc8466 (
      {stage1_59[278]},
      {stage2_59[124]}
   );
   gpc1_1 gpc8467 (
      {stage1_59[279]},
      {stage2_59[125]}
   );
   gpc1_1 gpc8468 (
      {stage1_59[280]},
      {stage2_59[126]}
   );
   gpc1_1 gpc8469 (
      {stage1_59[281]},
      {stage2_59[127]}
   );
   gpc1_1 gpc8470 (
      {stage1_59[282]},
      {stage2_59[128]}
   );
   gpc1_1 gpc8471 (
      {stage1_59[283]},
      {stage2_59[129]}
   );
   gpc1_1 gpc8472 (
      {stage1_59[284]},
      {stage2_59[130]}
   );
   gpc1_1 gpc8473 (
      {stage1_59[285]},
      {stage2_59[131]}
   );
   gpc1_1 gpc8474 (
      {stage1_59[286]},
      {stage2_59[132]}
   );
   gpc1_1 gpc8475 (
      {stage1_59[287]},
      {stage2_59[133]}
   );
   gpc1_1 gpc8476 (
      {stage1_59[288]},
      {stage2_59[134]}
   );
   gpc1_1 gpc8477 (
      {stage1_59[289]},
      {stage2_59[135]}
   );
   gpc1_1 gpc8478 (
      {stage1_59[290]},
      {stage2_59[136]}
   );
   gpc1_1 gpc8479 (
      {stage1_59[291]},
      {stage2_59[137]}
   );
   gpc1_1 gpc8480 (
      {stage1_59[292]},
      {stage2_59[138]}
   );
   gpc1_1 gpc8481 (
      {stage1_59[293]},
      {stage2_59[139]}
   );
   gpc1_1 gpc8482 (
      {stage1_60[190]},
      {stage2_60[101]}
   );
   gpc1_1 gpc8483 (
      {stage1_60[191]},
      {stage2_60[102]}
   );
   gpc1_1 gpc8484 (
      {stage1_60[192]},
      {stage2_60[103]}
   );
   gpc1_1 gpc8485 (
      {stage1_60[193]},
      {stage2_60[104]}
   );
   gpc1_1 gpc8486 (
      {stage1_60[194]},
      {stage2_60[105]}
   );
   gpc1_1 gpc8487 (
      {stage1_60[195]},
      {stage2_60[106]}
   );
   gpc1_1 gpc8488 (
      {stage1_60[196]},
      {stage2_60[107]}
   );
   gpc1_1 gpc8489 (
      {stage1_60[197]},
      {stage2_60[108]}
   );
   gpc1_1 gpc8490 (
      {stage1_60[198]},
      {stage2_60[109]}
   );
   gpc1_1 gpc8491 (
      {stage1_60[199]},
      {stage2_60[110]}
   );
   gpc1_1 gpc8492 (
      {stage1_61[198]},
      {stage2_61[83]}
   );
   gpc1_1 gpc8493 (
      {stage1_61[199]},
      {stage2_61[84]}
   );
   gpc1_1 gpc8494 (
      {stage1_61[200]},
      {stage2_61[85]}
   );
   gpc1_1 gpc8495 (
      {stage1_61[201]},
      {stage2_61[86]}
   );
   gpc1_1 gpc8496 (
      {stage1_61[202]},
      {stage2_61[87]}
   );
   gpc1_1 gpc8497 (
      {stage1_61[203]},
      {stage2_61[88]}
   );
   gpc1_1 gpc8498 (
      {stage1_61[204]},
      {stage2_61[89]}
   );
   gpc1_1 gpc8499 (
      {stage1_61[205]},
      {stage2_61[90]}
   );
   gpc1_1 gpc8500 (
      {stage1_61[206]},
      {stage2_61[91]}
   );
   gpc1_1 gpc8501 (
      {stage1_61[207]},
      {stage2_61[92]}
   );
   gpc1_1 gpc8502 (
      {stage1_61[208]},
      {stage2_61[93]}
   );
   gpc1_1 gpc8503 (
      {stage1_61[209]},
      {stage2_61[94]}
   );
   gpc1_1 gpc8504 (
      {stage1_61[210]},
      {stage2_61[95]}
   );
   gpc1_1 gpc8505 (
      {stage1_61[211]},
      {stage2_61[96]}
   );
   gpc1_1 gpc8506 (
      {stage1_61[212]},
      {stage2_61[97]}
   );
   gpc1_1 gpc8507 (
      {stage1_61[213]},
      {stage2_61[98]}
   );
   gpc1_1 gpc8508 (
      {stage1_61[214]},
      {stage2_61[99]}
   );
   gpc1_1 gpc8509 (
      {stage1_61[215]},
      {stage2_61[100]}
   );
   gpc1_1 gpc8510 (
      {stage1_61[216]},
      {stage2_61[101]}
   );
   gpc1_1 gpc8511 (
      {stage1_62[346]},
      {stage2_62[118]}
   );
   gpc1_1 gpc8512 (
      {stage1_62[347]},
      {stage2_62[119]}
   );
   gpc1_1 gpc8513 (
      {stage1_62[348]},
      {stage2_62[120]}
   );
   gpc1_1 gpc8514 (
      {stage1_62[349]},
      {stage2_62[121]}
   );
   gpc1_1 gpc8515 (
      {stage1_62[350]},
      {stage2_62[122]}
   );
   gpc1_1 gpc8516 (
      {stage1_62[351]},
      {stage2_62[123]}
   );
   gpc1_1 gpc8517 (
      {stage1_62[352]},
      {stage2_62[124]}
   );
   gpc1_1 gpc8518 (
      {stage1_62[353]},
      {stage2_62[125]}
   );
   gpc1_1 gpc8519 (
      {stage1_62[354]},
      {stage2_62[126]}
   );
   gpc1_1 gpc8520 (
      {stage1_62[355]},
      {stage2_62[127]}
   );
   gpc1_1 gpc8521 (
      {stage1_62[356]},
      {stage2_62[128]}
   );
   gpc1_1 gpc8522 (
      {stage1_62[357]},
      {stage2_62[129]}
   );
   gpc1_1 gpc8523 (
      {stage1_62[358]},
      {stage2_62[130]}
   );
   gpc1_1 gpc8524 (
      {stage1_62[359]},
      {stage2_62[131]}
   );
   gpc1_1 gpc8525 (
      {stage1_62[360]},
      {stage2_62[132]}
   );
   gpc1_1 gpc8526 (
      {stage1_62[361]},
      {stage2_62[133]}
   );
   gpc1_1 gpc8527 (
      {stage1_62[362]},
      {stage2_62[134]}
   );
   gpc1_1 gpc8528 (
      {stage1_62[363]},
      {stage2_62[135]}
   );
   gpc1_1 gpc8529 (
      {stage1_62[364]},
      {stage2_62[136]}
   );
   gpc1_1 gpc8530 (
      {stage1_62[365]},
      {stage2_62[137]}
   );
   gpc1_1 gpc8531 (
      {stage1_62[366]},
      {stage2_62[138]}
   );
   gpc1_1 gpc8532 (
      {stage1_62[367]},
      {stage2_62[139]}
   );
   gpc1_1 gpc8533 (
      {stage1_62[368]},
      {stage2_62[140]}
   );
   gpc1_1 gpc8534 (
      {stage1_62[369]},
      {stage2_62[141]}
   );
   gpc1_1 gpc8535 (
      {stage1_62[370]},
      {stage2_62[142]}
   );
   gpc1_1 gpc8536 (
      {stage1_62[371]},
      {stage2_62[143]}
   );
   gpc1_1 gpc8537 (
      {stage1_62[372]},
      {stage2_62[144]}
   );
   gpc1_1 gpc8538 (
      {stage1_64[94]},
      {stage2_64[84]}
   );
   gpc1_1 gpc8539 (
      {stage1_64[95]},
      {stage2_64[85]}
   );
   gpc1_1 gpc8540 (
      {stage1_64[96]},
      {stage2_64[86]}
   );
   gpc1_1 gpc8541 (
      {stage1_64[97]},
      {stage2_64[87]}
   );
   gpc1_1 gpc8542 (
      {stage1_64[98]},
      {stage2_64[88]}
   );
   gpc1_1 gpc8543 (
      {stage1_64[99]},
      {stage2_64[89]}
   );
   gpc1_1 gpc8544 (
      {stage1_64[100]},
      {stage2_64[90]}
   );
   gpc1_1 gpc8545 (
      {stage1_64[101]},
      {stage2_64[91]}
   );
   gpc1_1 gpc8546 (
      {stage1_64[102]},
      {stage2_64[92]}
   );
   gpc1_1 gpc8547 (
      {stage1_64[103]},
      {stage2_64[93]}
   );
   gpc1_1 gpc8548 (
      {stage1_64[104]},
      {stage2_64[94]}
   );
   gpc1_1 gpc8549 (
      {stage1_64[105]},
      {stage2_64[95]}
   );
   gpc1_1 gpc8550 (
      {stage1_64[106]},
      {stage2_64[96]}
   );
   gpc1_1 gpc8551 (
      {stage1_64[107]},
      {stage2_64[97]}
   );
   gpc1_1 gpc8552 (
      {stage1_64[108]},
      {stage2_64[98]}
   );
   gpc1_1 gpc8553 (
      {stage1_64[109]},
      {stage2_64[99]}
   );
   gpc1_1 gpc8554 (
      {stage1_64[110]},
      {stage2_64[100]}
   );
   gpc1_1 gpc8555 (
      {stage1_64[111]},
      {stage2_64[101]}
   );
   gpc1_1 gpc8556 (
      {stage1_65[46]},
      {stage2_65[57]}
   );
   gpc1_1 gpc8557 (
      {stage1_65[47]},
      {stage2_65[58]}
   );
   gpc1_1 gpc8558 (
      {stage1_65[48]},
      {stage2_65[59]}
   );
   gpc1_1 gpc8559 (
      {stage1_65[49]},
      {stage2_65[60]}
   );
   gpc1_1 gpc8560 (
      {stage1_65[50]},
      {stage2_65[61]}
   );
   gpc1_1 gpc8561 (
      {stage1_65[51]},
      {stage2_65[62]}
   );
   gpc1_1 gpc8562 (
      {stage1_65[52]},
      {stage2_65[63]}
   );
   gpc1_1 gpc8563 (
      {stage1_65[53]},
      {stage2_65[64]}
   );
   gpc1_1 gpc8564 (
      {stage1_65[54]},
      {stage2_65[65]}
   );
   gpc1_1 gpc8565 (
      {stage1_65[55]},
      {stage2_65[66]}
   );
   gpc1_1 gpc8566 (
      {stage1_65[56]},
      {stage2_65[67]}
   );
   gpc1163_5 gpc8567 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc8568 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc8569 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[6]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc8570 (
      {stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18]},
      {stage2_1[7]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc615_5 gpc8571 (
      {stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_1[8]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc615_5 gpc8572 (
      {stage2_0[24], stage2_0[25], stage2_0[26], stage2_0[27], stage2_0[28]},
      {stage2_1[9]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1343_5 gpc8573 (
      {stage2_1[10], stage2_1[11], stage2_1[12]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[1], stage2_3[2], stage2_3[3]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc1343_5 gpc8574 (
      {stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[1]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc8575 (
      {stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc8576 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage3_6[0],stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9]}
   );
   gpc606_5 gpc8577 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49], stage2_2[50]},
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage3_6[1],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc8578 (
      {stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54], stage2_2[55], stage2_2[56]},
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage3_6[2],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc606_5 gpc8579 (
      {stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60], stage2_2[61], stage2_2[62]},
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage3_6[3],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc8580 (
      {stage2_2[63], stage2_2[64], stage2_2[65], stage2_2[66], stage2_2[67], stage2_2[68]},
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage3_6[4],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc8581 (
      {stage2_2[69], stage2_2[70], stage2_2[71], stage2_2[72], 1'b0, 1'b0},
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage3_6[5],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc207_4 gpc8582 (
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_5[0], stage2_5[1]},
      {stage3_6[6],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc207_4 gpc8583 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26]},
      {stage2_5[2], stage2_5[3]},
      {stage3_6[7],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc207_4 gpc8584 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_5[4], stage2_5[5]},
      {stage3_6[8],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc207_4 gpc8585 (
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40]},
      {stage2_5[6], stage2_5[7]},
      {stage3_6[9],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc207_4 gpc8586 (
      {stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[8], stage2_5[9]},
      {stage3_6[10],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc207_4 gpc8587 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_5[10], stage2_5[11]},
      {stage3_6[11],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc207_4 gpc8588 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_5[12], stage2_5[13]},
      {stage3_6[12],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc207_4 gpc8589 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_5[14], stage2_5[15]},
      {stage3_6[13],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc207_4 gpc8590 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75]},
      {stage2_5[16], stage2_5[17]},
      {stage3_6[14],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc207_4 gpc8591 (
      {stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_5[18], stage2_5[19]},
      {stage3_6[15],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc207_4 gpc8592 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_5[20], stage2_5[21]},
      {stage3_6[16],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc207_4 gpc8593 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96]},
      {stage2_5[22], stage2_5[23]},
      {stage3_6[17],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc207_4 gpc8594 (
      {stage2_3[97], stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103]},
      {stage2_5[24], stage2_5[25]},
      {stage3_6[18],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc207_4 gpc8595 (
      {stage2_3[104], stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109], stage2_3[110]},
      {stage2_5[26], stage2_5[27]},
      {stage3_6[19],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc207_4 gpc8596 (
      {stage2_3[111], stage2_3[112], stage2_3[113], stage2_3[114], stage2_3[115], stage2_3[116], stage2_3[117]},
      {stage2_5[28], stage2_5[29]},
      {stage3_6[20],stage3_5[23],stage3_4[29],stage3_3[29]}
   );
   gpc207_4 gpc8597 (
      {stage2_3[118], stage2_3[119], stage2_3[120], stage2_3[121], stage2_3[122], stage2_3[123], stage2_3[124]},
      {stage2_5[30], stage2_5[31]},
      {stage3_6[21],stage3_5[24],stage3_4[30],stage3_3[30]}
   );
   gpc207_4 gpc8598 (
      {stage2_3[125], stage2_3[126], stage2_3[127], stage2_3[128], stage2_3[129], stage2_3[130], stage2_3[131]},
      {stage2_5[32], stage2_5[33]},
      {stage3_6[22],stage3_5[25],stage3_4[31],stage3_3[31]}
   );
   gpc207_4 gpc8599 (
      {stage2_3[132], stage2_3[133], stage2_3[134], stage2_3[135], stage2_3[136], stage2_3[137], stage2_3[138]},
      {stage2_5[34], stage2_5[35]},
      {stage3_6[23],stage3_5[26],stage3_4[32],stage3_3[32]}
   );
   gpc207_4 gpc8600 (
      {stage2_3[139], stage2_3[140], stage2_3[141], stage2_3[142], stage2_3[143], stage2_3[144], stage2_3[145]},
      {stage2_5[36], stage2_5[37]},
      {stage3_6[24],stage3_5[27],stage3_4[33],stage3_3[33]}
   );
   gpc207_4 gpc8601 (
      {stage2_3[146], stage2_3[147], stage2_3[148], stage2_3[149], stage2_3[150], stage2_3[151], stage2_3[152]},
      {stage2_5[38], stage2_5[39]},
      {stage3_6[25],stage3_5[28],stage3_4[34],stage3_3[34]}
   );
   gpc207_4 gpc8602 (
      {stage2_3[153], stage2_3[154], stage2_3[155], stage2_3[156], stage2_3[157], stage2_3[158], stage2_3[159]},
      {stage2_5[40], stage2_5[41]},
      {stage3_6[26],stage3_5[29],stage3_4[35],stage3_3[35]}
   );
   gpc207_4 gpc8603 (
      {stage2_3[160], stage2_3[161], stage2_3[162], stage2_3[163], stage2_3[164], stage2_3[165], stage2_3[166]},
      {stage2_5[42], stage2_5[43]},
      {stage3_6[27],stage3_5[30],stage3_4[36],stage3_3[36]}
   );
   gpc207_4 gpc8604 (
      {stage2_3[167], stage2_3[168], stage2_3[169], stage2_3[170], stage2_3[171], stage2_3[172], stage2_3[173]},
      {stage2_5[44], stage2_5[45]},
      {stage3_6[28],stage3_5[31],stage3_4[37],stage3_3[37]}
   );
   gpc207_4 gpc8605 (
      {stage2_3[174], stage2_3[175], stage2_3[176], stage2_3[177], stage2_3[178], stage2_3[179], stage2_3[180]},
      {stage2_5[46], stage2_5[47]},
      {stage3_6[29],stage3_5[32],stage3_4[38],stage3_3[38]}
   );
   gpc207_4 gpc8606 (
      {stage2_3[181], stage2_3[182], stage2_3[183], stage2_3[184], stage2_3[185], stage2_3[186], stage2_3[187]},
      {stage2_5[48], stage2_5[49]},
      {stage3_6[30],stage3_5[33],stage3_4[39],stage3_3[39]}
   );
   gpc207_4 gpc8607 (
      {stage2_3[188], stage2_3[189], stage2_3[190], stage2_3[191], stage2_3[192], stage2_3[193], stage2_3[194]},
      {stage2_5[50], stage2_5[51]},
      {stage3_6[31],stage3_5[34],stage3_4[40],stage3_3[40]}
   );
   gpc207_4 gpc8608 (
      {stage2_3[195], stage2_3[196], stage2_3[197], stage2_3[198], stage2_3[199], stage2_3[200], stage2_3[201]},
      {stage2_5[52], stage2_5[53]},
      {stage3_6[32],stage3_5[35],stage3_4[41],stage3_3[41]}
   );
   gpc207_4 gpc8609 (
      {stage2_3[202], stage2_3[203], stage2_3[204], stage2_3[205], stage2_3[206], stage2_3[207], stage2_3[208]},
      {stage2_5[54], stage2_5[55]},
      {stage3_6[33],stage3_5[36],stage3_4[42],stage3_3[42]}
   );
   gpc207_4 gpc8610 (
      {stage2_3[209], stage2_3[210], stage2_3[211], stage2_3[212], stage2_3[213], stage2_3[214], stage2_3[215]},
      {stage2_5[56], stage2_5[57]},
      {stage3_6[34],stage3_5[37],stage3_4[43],stage3_3[43]}
   );
   gpc615_5 gpc8611 (
      {stage2_3[216], stage2_3[217], stage2_3[218], stage2_3[219], stage2_3[220]},
      {stage2_4[38]},
      {stage2_5[58], stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63]},
      {stage3_7[0],stage3_6[35],stage3_5[38],stage3_4[44],stage3_3[44]}
   );
   gpc615_5 gpc8612 (
      {stage2_3[221], stage2_3[222], stage2_3[223], stage2_3[224], stage2_3[225]},
      {stage2_4[39]},
      {stage2_5[64], stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage3_7[1],stage3_6[36],stage3_5[39],stage3_4[45],stage3_3[45]}
   );
   gpc615_5 gpc8613 (
      {stage2_3[226], stage2_3[227], stage2_3[228], stage2_3[229], stage2_3[230]},
      {stage2_4[40]},
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75]},
      {stage3_7[2],stage3_6[37],stage3_5[40],stage3_4[46],stage3_3[46]}
   );
   gpc615_5 gpc8614 (
      {stage2_3[231], stage2_3[232], stage2_3[233], stage2_3[234], stage2_3[235]},
      {stage2_4[41]},
      {stage2_5[76], stage2_5[77], stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81]},
      {stage3_7[3],stage3_6[38],stage3_5[41],stage3_4[47],stage3_3[47]}
   );
   gpc615_5 gpc8615 (
      {stage2_3[236], stage2_3[237], stage2_3[238], stage2_3[239], stage2_3[240]},
      {stage2_4[42]},
      {stage2_5[82], stage2_5[83], stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87]},
      {stage3_7[4],stage3_6[39],stage3_5[42],stage3_4[48],stage3_3[48]}
   );
   gpc615_5 gpc8616 (
      {stage2_3[241], stage2_3[242], stage2_3[243], stage2_3[244], stage2_3[245]},
      {stage2_4[43]},
      {stage2_5[88], stage2_5[89], stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93]},
      {stage3_7[5],stage3_6[40],stage3_5[43],stage3_4[49],stage3_3[49]}
   );
   gpc615_5 gpc8617 (
      {stage2_3[246], stage2_3[247], stage2_3[248], stage2_3[249], stage2_3[250]},
      {stage2_4[44]},
      {stage2_5[94], stage2_5[95], stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99]},
      {stage3_7[6],stage3_6[41],stage3_5[44],stage3_4[50],stage3_3[50]}
   );
   gpc615_5 gpc8618 (
      {stage2_3[251], stage2_3[252], stage2_3[253], 1'b0, 1'b0},
      {stage2_4[45]},
      {stage2_5[100], stage2_5[101], stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105]},
      {stage3_7[7],stage3_6[42],stage3_5[45],stage3_4[51],stage3_3[51]}
   );
   gpc606_5 gpc8619 (
      {stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[43],stage3_5[46],stage3_4[52]}
   );
   gpc606_5 gpc8620 (
      {stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[44],stage3_5[47],stage3_4[53]}
   );
   gpc606_5 gpc8621 (
      {stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[45],stage3_5[48],stage3_4[54]}
   );
   gpc606_5 gpc8622 (
      {stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[46],stage3_5[49],stage3_4[55]}
   );
   gpc606_5 gpc8623 (
      {stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[47],stage3_5[50],stage3_4[56]}
   );
   gpc606_5 gpc8624 (
      {stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[48],stage3_5[51],stage3_4[57]}
   );
   gpc606_5 gpc8625 (
      {stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[14],stage3_6[49],stage3_5[52],stage3_4[58]}
   );
   gpc606_5 gpc8626 (
      {stage2_4[88], stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], 1'b0},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[15],stage3_6[50],stage3_5[53],stage3_4[59]}
   );
   gpc606_5 gpc8627 (
      {stage2_5[106], stage2_5[107], stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[16],stage3_6[51],stage3_5[54]}
   );
   gpc615_5 gpc8628 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[9],stage3_7[17],stage3_6[52]}
   );
   gpc615_5 gpc8629 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[7]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[10],stage3_7[18],stage3_6[53]}
   );
   gpc615_5 gpc8630 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[8]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[11],stage3_7[19],stage3_6[54]}
   );
   gpc615_5 gpc8631 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[9]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[4],stage3_8[12],stage3_7[20],stage3_6[55]}
   );
   gpc615_5 gpc8632 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[10]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[5],stage3_8[13],stage3_7[21],stage3_6[56]}
   );
   gpc615_5 gpc8633 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[11]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[6],stage3_8[14],stage3_7[22],stage3_6[57]}
   );
   gpc615_5 gpc8634 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[12]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[7],stage3_8[15],stage3_7[23],stage3_6[58]}
   );
   gpc615_5 gpc8635 (
      {stage2_6[83], stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87]},
      {stage2_7[13]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[8],stage3_8[16],stage3_7[24],stage3_6[59]}
   );
   gpc615_5 gpc8636 (
      {stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91], stage2_6[92]},
      {stage2_7[14]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[9],stage3_8[17],stage3_7[25],stage3_6[60]}
   );
   gpc615_5 gpc8637 (
      {stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_7[15]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[10],stage3_8[18],stage3_7[26],stage3_6[61]}
   );
   gpc615_5 gpc8638 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102]},
      {stage2_7[16]},
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage3_10[10],stage3_9[11],stage3_8[19],stage3_7[27],stage3_6[62]}
   );
   gpc615_5 gpc8639 (
      {stage2_6[103], stage2_6[104], stage2_6[105], stage2_6[106], stage2_6[107]},
      {stage2_7[17]},
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage3_10[11],stage3_9[12],stage3_8[20],stage3_7[28],stage3_6[63]}
   );
   gpc615_5 gpc8640 (
      {stage2_6[108], stage2_6[109], stage2_6[110], stage2_6[111], stage2_6[112]},
      {stage2_7[18]},
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage3_10[12],stage3_9[13],stage3_8[21],stage3_7[29],stage3_6[64]}
   );
   gpc615_5 gpc8641 (
      {stage2_6[113], stage2_6[114], stage2_6[115], stage2_6[116], stage2_6[117]},
      {stage2_7[19]},
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage3_10[13],stage3_9[14],stage3_8[22],stage3_7[30],stage3_6[65]}
   );
   gpc615_5 gpc8642 (
      {stage2_6[118], stage2_6[119], stage2_6[120], 1'b0, 1'b0},
      {stage2_7[20]},
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage3_10[14],stage3_9[15],stage3_8[23],stage3_7[31],stage3_6[66]}
   );
   gpc2116_5 gpc8643 (
      {stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[90]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[15],stage3_9[16],stage3_8[24],stage3_7[32]}
   );
   gpc2116_5 gpc8644 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[91]},
      {stage2_9[1]},
      {stage2_10[2], stage2_10[3]},
      {stage3_11[1],stage3_10[16],stage3_9[17],stage3_8[25],stage3_7[33]}
   );
   gpc2116_5 gpc8645 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[92]},
      {stage2_9[2]},
      {stage2_10[4], stage2_10[5]},
      {stage3_11[2],stage3_10[17],stage3_9[18],stage3_8[26],stage3_7[34]}
   );
   gpc2116_5 gpc8646 (
      {stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44]},
      {stage2_8[93]},
      {stage2_9[3]},
      {stage2_10[6], stage2_10[7]},
      {stage3_11[3],stage3_10[18],stage3_9[19],stage3_8[27],stage3_7[35]}
   );
   gpc2116_5 gpc8647 (
      {stage2_7[45], stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[94]},
      {stage2_9[4]},
      {stage2_10[8], stage2_10[9]},
      {stage3_11[4],stage3_10[19],stage3_9[20],stage3_8[28],stage3_7[36]}
   );
   gpc2116_5 gpc8648 (
      {stage2_7[51], stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[95]},
      {stage2_9[5]},
      {stage2_10[10], stage2_10[11]},
      {stage3_11[5],stage3_10[20],stage3_9[21],stage3_8[29],stage3_7[37]}
   );
   gpc2116_5 gpc8649 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62]},
      {stage2_8[96]},
      {stage2_9[6]},
      {stage2_10[12], stage2_10[13]},
      {stage3_11[6],stage3_10[21],stage3_9[22],stage3_8[30],stage3_7[38]}
   );
   gpc2116_5 gpc8650 (
      {stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[97]},
      {stage2_9[7]},
      {stage2_10[14], stage2_10[15]},
      {stage3_11[7],stage3_10[22],stage3_9[23],stage3_8[31],stage3_7[39]}
   );
   gpc2116_5 gpc8651 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73], stage2_7[74]},
      {stage2_8[98]},
      {stage2_9[8]},
      {stage2_10[16], stage2_10[17]},
      {stage3_11[8],stage3_10[23],stage3_9[24],stage3_8[32],stage3_7[40]}
   );
   gpc615_5 gpc8652 (
      {stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78], stage2_7[79]},
      {stage2_8[99]},
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage3_11[9],stage3_10[24],stage3_9[25],stage3_8[33],stage3_7[41]}
   );
   gpc615_5 gpc8653 (
      {stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83], stage2_7[84]},
      {stage2_8[100]},
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage3_11[10],stage3_10[25],stage3_9[26],stage3_8[34],stage3_7[42]}
   );
   gpc606_5 gpc8654 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[0],stage3_11[11],stage3_10[26],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc8655 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[1],stage3_11[12],stage3_10[27],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc8656 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[2],stage3_11[13],stage3_10[28],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc8657 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[3],stage3_11[14],stage3_10[29],stage3_9[30],stage3_8[38]}
   );
   gpc606_5 gpc8658 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[4],stage3_11[15],stage3_10[30],stage3_9[31],stage3_8[39]}
   );
   gpc606_5 gpc8659 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[5],stage3_11[16],stage3_10[31],stage3_9[32],stage3_8[40]}
   );
   gpc606_5 gpc8660 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[6],stage3_11[17],stage3_10[32],stage3_9[33],stage3_8[41]}
   );
   gpc606_5 gpc8661 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[7],stage3_11[18],stage3_10[33],stage3_9[34],stage3_8[42]}
   );
   gpc606_5 gpc8662 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[8],stage3_11[19],stage3_10[34],stage3_9[35],stage3_8[43]}
   );
   gpc606_5 gpc8663 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], stage2_8[160]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[9],stage3_11[20],stage3_10[35],stage3_9[36],stage3_8[44]}
   );
   gpc606_5 gpc8664 (
      {stage2_8[161], stage2_8[162], stage2_8[163], stage2_8[164], stage2_8[165], stage2_8[166]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[10],stage3_11[21],stage3_10[36],stage3_9[37],stage3_8[45]}
   );
   gpc606_5 gpc8665 (
      {stage2_8[167], stage2_8[168], stage2_8[169], stage2_8[170], stage2_8[171], stage2_8[172]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[11],stage3_11[22],stage3_10[37],stage3_9[38],stage3_8[46]}
   );
   gpc606_5 gpc8666 (
      {stage2_9[21], stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[12],stage3_11[23],stage3_10[38],stage3_9[39]}
   );
   gpc606_5 gpc8667 (
      {stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30], stage2_9[31], stage2_9[32]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[13],stage3_11[24],stage3_10[39],stage3_9[40]}
   );
   gpc606_5 gpc8668 (
      {stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37], stage2_9[38]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[14],stage3_11[25],stage3_10[40],stage3_9[41]}
   );
   gpc606_5 gpc8669 (
      {stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43], stage2_9[44]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[15],stage3_11[26],stage3_10[41],stage3_9[42]}
   );
   gpc606_5 gpc8670 (
      {stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49], stage2_9[50]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[16],stage3_11[27],stage3_10[42],stage3_9[43]}
   );
   gpc606_5 gpc8671 (
      {stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[17],stage3_11[28],stage3_10[43],stage3_9[44]}
   );
   gpc606_5 gpc8672 (
      {stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[18],stage3_11[29],stage3_10[44],stage3_9[45]}
   );
   gpc606_5 gpc8673 (
      {stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67], stage2_9[68]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[19],stage3_11[30],stage3_10[45],stage3_9[46]}
   );
   gpc606_5 gpc8674 (
      {stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[20],stage3_11[31],stage3_10[46],stage3_9[47]}
   );
   gpc606_5 gpc8675 (
      {stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[21],stage3_11[32],stage3_10[47],stage3_9[48]}
   );
   gpc606_5 gpc8676 (
      {stage2_9[81], stage2_9[82], stage2_9[83], stage2_9[84], stage2_9[85], stage2_9[86]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[22],stage3_11[33],stage3_10[48],stage3_9[49]}
   );
   gpc606_5 gpc8677 (
      {stage2_9[87], stage2_9[88], stage2_9[89], stage2_9[90], stage2_9[91], stage2_9[92]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[23],stage3_11[34],stage3_10[49],stage3_9[50]}
   );
   gpc606_5 gpc8678 (
      {stage2_9[93], stage2_9[94], stage2_9[95], stage2_9[96], stage2_9[97], stage2_9[98]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[24],stage3_11[35],stage3_10[50],stage3_9[51]}
   );
   gpc606_5 gpc8679 (
      {stage2_9[99], stage2_9[100], stage2_9[101], stage2_9[102], stage2_9[103], stage2_9[104]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[25],stage3_11[36],stage3_10[51],stage3_9[52]}
   );
   gpc215_4 gpc8680 (
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94]},
      {stage2_11[84]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[14],stage3_12[26],stage3_11[37],stage3_10[52]}
   );
   gpc215_4 gpc8681 (
      {stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99]},
      {stage2_11[85]},
      {stage2_12[2], stage2_12[3]},
      {stage3_13[15],stage3_12[27],stage3_11[38],stage3_10[53]}
   );
   gpc215_4 gpc8682 (
      {stage2_10[100], stage2_10[101], stage2_10[102], stage2_10[103], stage2_10[104]},
      {stage2_11[86]},
      {stage2_12[4], stage2_12[5]},
      {stage3_13[16],stage3_12[28],stage3_11[39],stage3_10[54]}
   );
   gpc615_5 gpc8683 (
      {stage2_10[105], stage2_10[106], stage2_10[107], stage2_10[108], stage2_10[109]},
      {stage2_11[87]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[0],stage3_13[17],stage3_12[29],stage3_11[40],stage3_10[55]}
   );
   gpc615_5 gpc8684 (
      {stage2_10[110], stage2_10[111], stage2_10[112], stage2_10[113], stage2_10[114]},
      {stage2_11[88]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[1],stage3_13[18],stage3_12[30],stage3_11[41],stage3_10[56]}
   );
   gpc615_5 gpc8685 (
      {stage2_10[115], stage2_10[116], stage2_10[117], stage2_10[118], stage2_10[119]},
      {stage2_11[89]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[2],stage3_13[19],stage3_12[31],stage3_11[42],stage3_10[57]}
   );
   gpc615_5 gpc8686 (
      {stage2_10[120], stage2_10[121], stage2_10[122], stage2_10[123], stage2_10[124]},
      {stage2_11[90]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[3],stage3_13[20],stage3_12[32],stage3_11[43],stage3_10[58]}
   );
   gpc606_5 gpc8687 (
      {stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[4],stage3_13[21],stage3_12[33],stage3_11[44]}
   );
   gpc606_5 gpc8688 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[5],stage3_13[22],stage3_12[34],stage3_11[45]}
   );
   gpc606_5 gpc8689 (
      {stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[6],stage3_13[23],stage3_12[35],stage3_11[46]}
   );
   gpc606_5 gpc8690 (
      {stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[7],stage3_13[24],stage3_12[36],stage3_11[47]}
   );
   gpc615_5 gpc8691 (
      {stage2_11[115], stage2_11[116], stage2_11[117], stage2_11[118], stage2_11[119]},
      {stage2_12[30]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[8],stage3_13[25],stage3_12[37],stage3_11[48]}
   );
   gpc615_5 gpc8692 (
      {stage2_11[120], stage2_11[121], stage2_11[122], stage2_11[123], stage2_11[124]},
      {stage2_12[31]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[9],stage3_13[26],stage3_12[38],stage3_11[49]}
   );
   gpc606_5 gpc8693 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[6],stage3_14[10],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc8694 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[7],stage3_14[11],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc8695 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[8],stage3_14[12],stage3_13[29],stage3_12[41]}
   );
   gpc606_5 gpc8696 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[9],stage3_14[13],stage3_13[30],stage3_12[42]}
   );
   gpc606_5 gpc8697 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[10],stage3_14[14],stage3_13[31],stage3_12[43]}
   );
   gpc606_5 gpc8698 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[11],stage3_14[15],stage3_13[32],stage3_12[44]}
   );
   gpc606_5 gpc8699 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[12],stage3_14[16],stage3_13[33],stage3_12[45]}
   );
   gpc606_5 gpc8700 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[13],stage3_14[17],stage3_13[34],stage3_12[46]}
   );
   gpc606_5 gpc8701 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[14],stage3_14[18],stage3_13[35],stage3_12[47]}
   );
   gpc606_5 gpc8702 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[15],stage3_14[19],stage3_13[36],stage3_12[48]}
   );
   gpc623_5 gpc8703 (
      {stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_13[36], stage2_13[37]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[16],stage3_14[20],stage3_13[37],stage3_12[49]}
   );
   gpc623_5 gpc8704 (
      {stage2_12[95], stage2_12[96], stage2_12[97]},
      {stage2_13[38], stage2_13[39]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[17],stage3_14[21],stage3_13[38],stage3_12[50]}
   );
   gpc615_5 gpc8705 (
      {stage2_13[40], stage2_13[41], stage2_13[42], stage2_13[43], stage2_13[44]},
      {stage2_14[72]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[18],stage3_14[22],stage3_13[39]}
   );
   gpc615_5 gpc8706 (
      {stage2_13[45], stage2_13[46], stage2_13[47], stage2_13[48], stage2_13[49]},
      {stage2_14[73]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[19],stage3_14[23],stage3_13[40]}
   );
   gpc615_5 gpc8707 (
      {stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53], stage2_13[54]},
      {stage2_14[74]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[20],stage3_14[24],stage3_13[41]}
   );
   gpc615_5 gpc8708 (
      {stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_14[75]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[21],stage3_14[25],stage3_13[42]}
   );
   gpc615_5 gpc8709 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64]},
      {stage2_14[76]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[22],stage3_14[26],stage3_13[43]}
   );
   gpc615_5 gpc8710 (
      {stage2_13[65], stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69]},
      {stage2_14[77]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[23],stage3_14[27],stage3_13[44]}
   );
   gpc606_5 gpc8711 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[18],stage3_15[24],stage3_14[28]}
   );
   gpc606_5 gpc8712 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[19],stage3_15[25],stage3_14[29]}
   );
   gpc615_5 gpc8713 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94]},
      {stage2_15[36]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[20],stage3_15[26],stage3_14[30]}
   );
   gpc615_5 gpc8714 (
      {stage2_14[95], stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99]},
      {stage2_15[37]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[21],stage3_15[27],stage3_14[31]}
   );
   gpc615_5 gpc8715 (
      {stage2_14[100], stage2_14[101], stage2_14[102], stage2_14[103], stage2_14[104]},
      {stage2_15[38]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[22],stage3_15[28],stage3_14[32]}
   );
   gpc615_5 gpc8716 (
      {stage2_14[105], stage2_14[106], stage2_14[107], stage2_14[108], stage2_14[109]},
      {stage2_15[39]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[23],stage3_15[29],stage3_14[33]}
   );
   gpc615_5 gpc8717 (
      {stage2_14[110], stage2_14[111], stage2_14[112], stage2_14[113], stage2_14[114]},
      {stage2_15[40]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[24],stage3_15[30],stage3_14[34]}
   );
   gpc207_4 gpc8718 (
      {stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[7],stage3_17[13],stage3_16[25],stage3_15[31]}
   );
   gpc615_5 gpc8719 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[42]},
      {stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7]},
      {stage3_19[0],stage3_18[8],stage3_17[14],stage3_16[26],stage3_15[32]}
   );
   gpc615_5 gpc8720 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[43]},
      {stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13]},
      {stage3_19[1],stage3_18[9],stage3_17[15],stage3_16[27],stage3_15[33]}
   );
   gpc615_5 gpc8721 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[44]},
      {stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19]},
      {stage3_19[2],stage3_18[10],stage3_17[16],stage3_16[28],stage3_15[34]}
   );
   gpc615_5 gpc8722 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[45]},
      {stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25]},
      {stage3_19[3],stage3_18[11],stage3_17[17],stage3_16[29],stage3_15[35]}
   );
   gpc615_5 gpc8723 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[46]},
      {stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31]},
      {stage3_19[4],stage3_18[12],stage3_17[18],stage3_16[30],stage3_15[36]}
   );
   gpc615_5 gpc8724 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[47]},
      {stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37]},
      {stage3_19[5],stage3_18[13],stage3_17[19],stage3_16[31],stage3_15[37]}
   );
   gpc615_5 gpc8725 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[48]},
      {stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43]},
      {stage3_19[6],stage3_18[14],stage3_17[20],stage3_16[32],stage3_15[38]}
   );
   gpc615_5 gpc8726 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[49]},
      {stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49]},
      {stage3_19[7],stage3_18[15],stage3_17[21],stage3_16[33],stage3_15[39]}
   );
   gpc615_5 gpc8727 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[50]},
      {stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55]},
      {stage3_19[8],stage3_18[16],stage3_17[22],stage3_16[34],stage3_15[40]}
   );
   gpc615_5 gpc8728 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[51]},
      {stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61]},
      {stage3_19[9],stage3_18[17],stage3_17[23],stage3_16[35],stage3_15[41]}
   );
   gpc615_5 gpc8729 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[52]},
      {stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67]},
      {stage3_19[10],stage3_18[18],stage3_17[24],stage3_16[36],stage3_15[42]}
   );
   gpc615_5 gpc8730 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[53]},
      {stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73]},
      {stage3_19[11],stage3_18[19],stage3_17[25],stage3_16[37],stage3_15[43]}
   );
   gpc606_5 gpc8731 (
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[12],stage3_18[20],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc8732 (
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[13],stage3_18[21],stage3_17[27],stage3_16[39]}
   );
   gpc606_5 gpc8733 (
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[14],stage3_18[22],stage3_17[28],stage3_16[40]}
   );
   gpc606_5 gpc8734 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[15],stage3_18[23],stage3_17[29],stage3_16[41]}
   );
   gpc606_5 gpc8735 (
      {stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[16],stage3_18[24],stage3_17[30],stage3_16[42]}
   );
   gpc606_5 gpc8736 (
      {stage2_16[84], stage2_16[85], stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89]},
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage3_20[5],stage3_19[17],stage3_18[25],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc8737 (
      {stage2_16[90], stage2_16[91], stage2_16[92], stage2_16[93], stage2_16[94], stage2_16[95]},
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41]},
      {stage3_20[6],stage3_19[18],stage3_18[26],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc8738 (
      {stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[7],stage3_19[19],stage3_18[27],stage3_17[33]}
   );
   gpc2135_5 gpc8739 (
      {stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[1],stage3_20[8],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc8740 (
      {stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50], stage2_18[51]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[2],stage3_20[9],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc8741 (
      {stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55], stage2_18[56]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[3],stage3_20[10],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc8742 (
      {stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60], stage2_18[61]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[4],stage3_20[11],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc8743 (
      {stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[5],stage3_20[12],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc8744 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[6],stage3_20[13],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc8745 (
      {stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75], stage2_18[76]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[7],stage3_20[14],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc8746 (
      {stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80], stage2_18[81]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[8],stage3_20[15],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc8747 (
      {stage2_18[82], stage2_18[83], stage2_18[84], stage2_18[85], stage2_18[86]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[9],stage3_20[16],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc8748 (
      {stage2_18[87], stage2_18[88], stage2_18[89], stage2_18[90], stage2_18[91]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[10],stage3_20[17],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc8749 (
      {stage2_18[92], stage2_18[93], stage2_18[94], stage2_18[95], stage2_18[96]},
      {stage2_19[36], stage2_19[37], stage2_19[38]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[11],stage3_20[18],stage3_19[30],stage3_18[38]}
   );
   gpc2135_5 gpc8750 (
      {stage2_18[97], stage2_18[98], stage2_18[99], stage2_18[100], stage2_18[101]},
      {stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[12],stage3_20[19],stage3_19[31],stage3_18[39]}
   );
   gpc2135_5 gpc8751 (
      {stage2_18[102], stage2_18[103], stage2_18[104], stage2_18[105], stage2_18[106]},
      {stage2_19[42], stage2_19[43], stage2_19[44]},
      {stage2_20[12]},
      {stage2_21[24], stage2_21[25]},
      {stage3_22[12],stage3_21[13],stage3_20[20],stage3_19[32],stage3_18[40]}
   );
   gpc2135_5 gpc8752 (
      {stage2_18[107], stage2_18[108], stage2_18[109], stage2_18[110], stage2_18[111]},
      {stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[13]},
      {stage2_21[26], stage2_21[27]},
      {stage3_22[13],stage3_21[14],stage3_20[21],stage3_19[33],stage3_18[41]}
   );
   gpc2135_5 gpc8753 (
      {stage2_18[112], stage2_18[113], stage2_18[114], stage2_18[115], stage2_18[116]},
      {stage2_19[48], stage2_19[49], stage2_19[50]},
      {stage2_20[14]},
      {stage2_21[28], stage2_21[29]},
      {stage3_22[14],stage3_21[15],stage3_20[22],stage3_19[34],stage3_18[42]}
   );
   gpc2135_5 gpc8754 (
      {stage2_18[117], stage2_18[118], stage2_18[119], stage2_18[120], stage2_18[121]},
      {stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_20[15]},
      {stage2_21[30], stage2_21[31]},
      {stage3_22[15],stage3_21[16],stage3_20[23],stage3_19[35],stage3_18[43]}
   );
   gpc2135_5 gpc8755 (
      {stage2_18[122], stage2_18[123], stage2_18[124], stage2_18[125], stage2_18[126]},
      {stage2_19[54], stage2_19[55], stage2_19[56]},
      {stage2_20[16]},
      {stage2_21[32], stage2_21[33]},
      {stage3_22[16],stage3_21[17],stage3_20[24],stage3_19[36],stage3_18[44]}
   );
   gpc2135_5 gpc8756 (
      {stage2_18[127], stage2_18[128], stage2_18[129], stage2_18[130], stage2_18[131]},
      {stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage2_20[17]},
      {stage2_21[34], stage2_21[35]},
      {stage3_22[17],stage3_21[18],stage3_20[25],stage3_19[37],stage3_18[45]}
   );
   gpc2135_5 gpc8757 (
      {stage2_18[132], stage2_18[133], stage2_18[134], stage2_18[135], stage2_18[136]},
      {stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[18]},
      {stage2_21[36], stage2_21[37]},
      {stage3_22[18],stage3_21[19],stage3_20[26],stage3_19[38],stage3_18[46]}
   );
   gpc2135_5 gpc8758 (
      {stage2_18[137], stage2_18[138], stage2_18[139], stage2_18[140], stage2_18[141]},
      {stage2_19[63], stage2_19[64], stage2_19[65]},
      {stage2_20[19]},
      {stage2_21[38], stage2_21[39]},
      {stage3_22[19],stage3_21[20],stage3_20[27],stage3_19[39],stage3_18[47]}
   );
   gpc2135_5 gpc8759 (
      {stage2_18[142], stage2_18[143], stage2_18[144], stage2_18[145], stage2_18[146]},
      {stage2_19[66], stage2_19[67], stage2_19[68]},
      {stage2_20[20]},
      {stage2_21[40], stage2_21[41]},
      {stage3_22[20],stage3_21[21],stage3_20[28],stage3_19[40],stage3_18[48]}
   );
   gpc615_5 gpc8760 (
      {stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72], stage2_19[73]},
      {stage2_20[21]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[0],stage3_22[21],stage3_21[22],stage3_20[29],stage3_19[41]}
   );
   gpc615_5 gpc8761 (
      {stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77], stage2_19[78]},
      {stage2_20[22]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[1],stage3_22[22],stage3_21[23],stage3_20[30],stage3_19[42]}
   );
   gpc615_5 gpc8762 (
      {stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82], stage2_19[83]},
      {stage2_20[23]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[2],stage3_22[23],stage3_21[24],stage3_20[31],stage3_19[43]}
   );
   gpc615_5 gpc8763 (
      {stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87], stage2_19[88]},
      {stage2_20[24]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[3],stage3_22[24],stage3_21[25],stage3_20[32],stage3_19[44]}
   );
   gpc615_5 gpc8764 (
      {stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92], stage2_19[93]},
      {stage2_20[25]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[4],stage3_22[25],stage3_21[26],stage3_20[33],stage3_19[45]}
   );
   gpc606_5 gpc8765 (
      {stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30], stage2_20[31]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[26],stage3_21[27],stage3_20[34]}
   );
   gpc606_5 gpc8766 (
      {stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35], stage2_20[36], stage2_20[37]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[27],stage3_21[28],stage3_20[35]}
   );
   gpc606_5 gpc8767 (
      {stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[28],stage3_21[29],stage3_20[36]}
   );
   gpc606_5 gpc8768 (
      {stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47], stage2_20[48], stage2_20[49]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[8],stage3_22[29],stage3_21[30],stage3_20[37]}
   );
   gpc606_5 gpc8769 (
      {stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53], stage2_20[54], stage2_20[55]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[9],stage3_22[30],stage3_21[31],stage3_20[38]}
   );
   gpc606_5 gpc8770 (
      {stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59], stage2_20[60], stage2_20[61]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[10],stage3_22[31],stage3_21[32],stage3_20[39]}
   );
   gpc615_5 gpc8771 (
      {stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65], stage2_20[66]},
      {stage2_21[72]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[11],stage3_22[32],stage3_21[33],stage3_20[40]}
   );
   gpc615_5 gpc8772 (
      {stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage2_21[73]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage3_24[7],stage3_23[12],stage3_22[33],stage3_21[34],stage3_20[41]}
   );
   gpc606_5 gpc8773 (
      {stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77], stage2_21[78], stage2_21[79]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[8],stage3_23[13],stage3_22[34],stage3_21[35]}
   );
   gpc606_5 gpc8774 (
      {stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83], stage2_21[84], stage2_21[85]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[9],stage3_23[14],stage3_22[35],stage3_21[36]}
   );
   gpc615_5 gpc8775 (
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[10],stage3_23[15],stage3_22[36]}
   );
   gpc615_5 gpc8776 (
      {stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[11],stage3_23[16],stage3_22[37]}
   );
   gpc615_5 gpc8777 (
      {stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61], stage2_22[62]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[12],stage3_23[17],stage3_22[38]}
   );
   gpc615_5 gpc8778 (
      {stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66], stage2_22[67]},
      {stage2_23[15]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[5],stage3_24[13],stage3_23[18],stage3_22[39]}
   );
   gpc615_5 gpc8779 (
      {stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71], stage2_22[72]},
      {stage2_23[16]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[6],stage3_24[14],stage3_23[19],stage3_22[40]}
   );
   gpc615_5 gpc8780 (
      {stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76], stage2_22[77]},
      {stage2_23[17]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[7],stage3_24[15],stage3_23[20],stage3_22[41]}
   );
   gpc615_5 gpc8781 (
      {stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81], stage2_22[82]},
      {stage2_23[18]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[8],stage3_24[16],stage3_23[21],stage3_22[42]}
   );
   gpc615_5 gpc8782 (
      {stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86], stage2_22[87]},
      {stage2_23[19]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[9],stage3_24[17],stage3_23[22],stage3_22[43]}
   );
   gpc615_5 gpc8783 (
      {stage2_22[88], stage2_22[89], stage2_22[90], stage2_22[91], stage2_22[92]},
      {stage2_23[20]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[10],stage3_24[18],stage3_23[23],stage3_22[44]}
   );
   gpc615_5 gpc8784 (
      {stage2_22[93], stage2_22[94], stage2_22[95], stage2_22[96], stage2_22[97]},
      {stage2_23[21]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[11],stage3_24[19],stage3_23[24],stage3_22[45]}
   );
   gpc615_5 gpc8785 (
      {stage2_22[98], stage2_22[99], stage2_22[100], stage2_22[101], stage2_22[102]},
      {stage2_23[22]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[12],stage3_24[20],stage3_23[25],stage3_22[46]}
   );
   gpc615_5 gpc8786 (
      {stage2_22[103], stage2_22[104], stage2_22[105], stage2_22[106], stage2_22[107]},
      {stage2_23[23]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[13],stage3_24[21],stage3_23[26],stage3_22[47]}
   );
   gpc615_5 gpc8787 (
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28]},
      {stage2_24[72]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[12],stage3_25[14],stage3_24[22],stage3_23[27]}
   );
   gpc615_5 gpc8788 (
      {stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33]},
      {stage2_24[73]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[13],stage3_25[15],stage3_24[23],stage3_23[28]}
   );
   gpc615_5 gpc8789 (
      {stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage2_24[74]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[14],stage3_25[16],stage3_24[24],stage3_23[29]}
   );
   gpc615_5 gpc8790 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43]},
      {stage2_24[75]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[15],stage3_25[17],stage3_24[25],stage3_23[30]}
   );
   gpc615_5 gpc8791 (
      {stage2_23[44], stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48]},
      {stage2_24[76]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[16],stage3_25[18],stage3_24[26],stage3_23[31]}
   );
   gpc615_5 gpc8792 (
      {stage2_23[49], stage2_23[50], stage2_23[51], stage2_23[52], stage2_23[53]},
      {stage2_24[77]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[17],stage3_25[19],stage3_24[27],stage3_23[32]}
   );
   gpc615_5 gpc8793 (
      {stage2_23[54], stage2_23[55], stage2_23[56], stage2_23[57], stage2_23[58]},
      {stage2_24[78]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[18],stage3_25[20],stage3_24[28],stage3_23[33]}
   );
   gpc615_5 gpc8794 (
      {stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62], stage2_23[63]},
      {stage2_24[79]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[19],stage3_25[21],stage3_24[29],stage3_23[34]}
   );
   gpc615_5 gpc8795 (
      {stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_24[80]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[20],stage3_25[22],stage3_24[30],stage3_23[35]}
   );
   gpc615_5 gpc8796 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73]},
      {stage2_24[81]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[21],stage3_25[23],stage3_24[31],stage3_23[36]}
   );
   gpc615_5 gpc8797 (
      {stage2_23[74], stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78]},
      {stage2_24[82]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[22],stage3_25[24],stage3_24[32],stage3_23[37]}
   );
   gpc615_5 gpc8798 (
      {stage2_23[79], stage2_23[80], stage2_23[81], stage2_23[82], stage2_23[83]},
      {stage2_24[83]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[23],stage3_25[25],stage3_24[33],stage3_23[38]}
   );
   gpc615_5 gpc8799 (
      {stage2_23[84], stage2_23[85], stage2_23[86], stage2_23[87], stage2_23[88]},
      {stage2_24[84]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[24],stage3_25[26],stage3_24[34],stage3_23[39]}
   );
   gpc606_5 gpc8800 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[13],stage3_26[25],stage3_25[27]}
   );
   gpc606_5 gpc8801 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[1],stage3_27[14],stage3_26[26],stage3_25[28]}
   );
   gpc606_5 gpc8802 (
      {stage2_25[90], stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[2],stage3_27[15],stage3_26[27],stage3_25[29]}
   );
   gpc606_5 gpc8803 (
      {stage2_25[96], stage2_25[97], stage2_25[98], stage2_25[99], stage2_25[100], stage2_25[101]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[3],stage3_27[16],stage3_26[28],stage3_25[30]}
   );
   gpc117_4 gpc8804 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6]},
      {stage2_27[24]},
      {stage2_28[0]},
      {stage3_29[4],stage3_28[4],stage3_27[17],stage3_26[29]}
   );
   gpc117_4 gpc8805 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12], stage2_26[13]},
      {stage2_27[25]},
      {stage2_28[1]},
      {stage3_29[5],stage3_28[5],stage3_27[18],stage3_26[30]}
   );
   gpc117_4 gpc8806 (
      {stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_27[26]},
      {stage2_28[2]},
      {stage3_29[6],stage3_28[6],stage3_27[19],stage3_26[31]}
   );
   gpc117_4 gpc8807 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[27]},
      {stage2_28[3]},
      {stage3_29[7],stage3_28[7],stage3_27[20],stage3_26[32]}
   );
   gpc117_4 gpc8808 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34]},
      {stage2_27[28]},
      {stage2_28[4]},
      {stage3_29[8],stage3_28[8],stage3_27[21],stage3_26[33]}
   );
   gpc117_4 gpc8809 (
      {stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage2_27[29]},
      {stage2_28[5]},
      {stage3_29[9],stage3_28[9],stage3_27[22],stage3_26[34]}
   );
   gpc117_4 gpc8810 (
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48]},
      {stage2_27[30]},
      {stage2_28[6]},
      {stage3_29[10],stage3_28[10],stage3_27[23],stage3_26[35]}
   );
   gpc117_4 gpc8811 (
      {stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55]},
      {stage2_27[31]},
      {stage2_28[7]},
      {stage3_29[11],stage3_28[11],stage3_27[24],stage3_26[36]}
   );
   gpc117_4 gpc8812 (
      {stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[32]},
      {stage2_28[8]},
      {stage3_29[12],stage3_28[12],stage3_27[25],stage3_26[37]}
   );
   gpc117_4 gpc8813 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69]},
      {stage2_27[33]},
      {stage2_28[9]},
      {stage3_29[13],stage3_28[13],stage3_27[26],stage3_26[38]}
   );
   gpc117_4 gpc8814 (
      {stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76]},
      {stage2_27[34]},
      {stage2_28[10]},
      {stage3_29[14],stage3_28[14],stage3_27[27],stage3_26[39]}
   );
   gpc117_4 gpc8815 (
      {stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage2_27[35]},
      {stage2_28[11]},
      {stage3_29[15],stage3_28[15],stage3_27[28],stage3_26[40]}
   );
   gpc117_4 gpc8816 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88], stage2_26[89], stage2_26[90]},
      {stage2_27[36]},
      {stage2_28[12]},
      {stage3_29[16],stage3_28[16],stage3_27[29],stage3_26[41]}
   );
   gpc117_4 gpc8817 (
      {stage2_26[91], stage2_26[92], stage2_26[93], stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97]},
      {stage2_27[37]},
      {stage2_28[13]},
      {stage3_29[17],stage3_28[17],stage3_27[30],stage3_26[42]}
   );
   gpc117_4 gpc8818 (
      {stage2_26[98], stage2_26[99], stage2_26[100], stage2_26[101], stage2_26[102], stage2_26[103], stage2_26[104]},
      {stage2_27[38]},
      {stage2_28[14]},
      {stage3_29[18],stage3_28[18],stage3_27[31],stage3_26[43]}
   );
   gpc117_4 gpc8819 (
      {stage2_26[105], stage2_26[106], stage2_26[107], stage2_26[108], stage2_26[109], stage2_26[110], stage2_26[111]},
      {stage2_27[39]},
      {stage2_28[15]},
      {stage3_29[19],stage3_28[19],stage3_27[32],stage3_26[44]}
   );
   gpc117_4 gpc8820 (
      {stage2_26[112], stage2_26[113], stage2_26[114], stage2_26[115], stage2_26[116], stage2_26[117], stage2_26[118]},
      {stage2_27[40]},
      {stage2_28[16]},
      {stage3_29[20],stage3_28[20],stage3_27[33],stage3_26[45]}
   );
   gpc117_4 gpc8821 (
      {stage2_26[119], stage2_26[120], stage2_26[121], stage2_26[122], stage2_26[123], stage2_26[124], stage2_26[125]},
      {stage2_27[41]},
      {stage2_28[17]},
      {stage3_29[21],stage3_28[21],stage3_27[34],stage3_26[46]}
   );
   gpc7_3 gpc8822 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48]},
      {stage3_29[22],stage3_28[22],stage3_27[35]}
   );
   gpc7_3 gpc8823 (
      {stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55]},
      {stage3_29[23],stage3_28[23],stage3_27[36]}
   );
   gpc207_4 gpc8824 (
      {stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_29[0], stage2_29[1]},
      {stage3_30[0],stage3_29[24],stage3_28[24],stage3_27[37]}
   );
   gpc207_4 gpc8825 (
      {stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_29[2], stage2_29[3]},
      {stage3_30[1],stage3_29[25],stage3_28[25],stage3_27[38]}
   );
   gpc606_5 gpc8826 (
      {stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73], stage2_27[74], stage2_27[75]},
      {stage2_29[4], stage2_29[5], stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9]},
      {stage3_31[0],stage3_30[2],stage3_29[26],stage3_28[26],stage3_27[39]}
   );
   gpc606_5 gpc8827 (
      {stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80], stage2_27[81]},
      {stage2_29[10], stage2_29[11], stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15]},
      {stage3_31[1],stage3_30[3],stage3_29[27],stage3_28[27],stage3_27[40]}
   );
   gpc615_5 gpc8828 (
      {stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], 1'b0},
      {stage2_28[18]},
      {stage2_29[16], stage2_29[17], stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage3_31[2],stage3_30[4],stage3_29[28],stage3_28[28],stage3_27[41]}
   );
   gpc615_5 gpc8829 (
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_29[22]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[5],stage3_29[29],stage3_28[29]}
   );
   gpc615_5 gpc8830 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[23]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[6],stage3_29[30],stage3_28[30]}
   );
   gpc615_5 gpc8831 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[24]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[7],stage3_29[31],stage3_28[31]}
   );
   gpc615_5 gpc8832 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[25]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[8],stage3_29[32],stage3_28[32]}
   );
   gpc615_5 gpc8833 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[26]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[7],stage3_30[9],stage3_29[33],stage3_28[33]}
   );
   gpc1163_5 gpc8834 (
      {stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[5],stage3_31[8],stage3_30[10],stage3_29[34]}
   );
   gpc1163_5 gpc8835 (
      {stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[6],stage3_31[9],stage3_30[11],stage3_29[35]}
   );
   gpc1163_5 gpc8836 (
      {stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[7],stage3_31[10],stage3_30[12],stage3_29[36]}
   );
   gpc1163_5 gpc8837 (
      {stage2_29[36], stage2_29[37], stage2_29[38]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[8],stage3_31[11],stage3_30[13],stage3_29[37]}
   );
   gpc1163_5 gpc8838 (
      {stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[9],stage3_31[12],stage3_30[14],stage3_29[38]}
   );
   gpc606_5 gpc8839 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[10],stage3_31[13],stage3_30[15],stage3_29[39]}
   );
   gpc606_5 gpc8840 (
      {stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[11],stage3_31[14],stage3_30[16],stage3_29[40]}
   );
   gpc606_5 gpc8841 (
      {stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[12],stage3_31[15],stage3_30[17],stage3_29[41]}
   );
   gpc606_5 gpc8842 (
      {stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[13],stage3_31[16],stage3_30[18],stage3_29[42]}
   );
   gpc606_5 gpc8843 (
      {stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[14],stage3_31[17],stage3_30[19],stage3_29[43]}
   );
   gpc606_5 gpc8844 (
      {stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[15],stage3_31[18],stage3_30[20],stage3_29[44]}
   );
   gpc606_5 gpc8845 (
      {stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[16],stage3_31[19],stage3_30[21],stage3_29[45]}
   );
   gpc606_5 gpc8846 (
      {stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[17],stage3_31[20],stage3_30[22],stage3_29[46]}
   );
   gpc606_5 gpc8847 (
      {stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[18],stage3_31[21],stage3_30[23],stage3_29[47]}
   );
   gpc606_5 gpc8848 (
      {stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101]},
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage3_33[14],stage3_32[19],stage3_31[22],stage3_30[24],stage3_29[48]}
   );
   gpc1163_5 gpc8849 (
      {stage2_30[60], stage2_30[61], stage2_30[62]},
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_32[5]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[15],stage3_32[20],stage3_31[23],stage3_30[25]}
   );
   gpc615_5 gpc8850 (
      {stage2_30[63], stage2_30[64], stage2_30[65], stage2_30[66], stage2_30[67]},
      {stage2_31[71]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[16],stage3_32[21],stage3_31[24],stage3_30[26]}
   );
   gpc615_5 gpc8851 (
      {stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71], stage2_30[72]},
      {stage2_31[72]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[17],stage3_32[22],stage3_31[25],stage3_30[27]}
   );
   gpc615_5 gpc8852 (
      {stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[73]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[18],stage3_32[23],stage3_31[26],stage3_30[28]}
   );
   gpc615_5 gpc8853 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82]},
      {stage2_31[74]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[19],stage3_32[24],stage3_31[27],stage3_30[29]}
   );
   gpc615_5 gpc8854 (
      {stage2_30[83], stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87]},
      {stage2_31[75]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[20],stage3_32[25],stage3_31[28],stage3_30[30]}
   );
   gpc615_5 gpc8855 (
      {stage2_30[88], stage2_30[89], stage2_30[90], stage2_30[91], stage2_30[92]},
      {stage2_31[76]},
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40], stage2_32[41]},
      {stage3_34[6],stage3_33[21],stage3_32[26],stage3_31[29],stage3_30[31]}
   );
   gpc606_5 gpc8856 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[0],stage3_34[7],stage3_33[22],stage3_32[27],stage3_31[30]}
   );
   gpc606_5 gpc8857 (
      {stage2_31[83], stage2_31[84], stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88]},
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12]},
      {stage3_35[1],stage3_34[8],stage3_33[23],stage3_32[28],stage3_31[31]}
   );
   gpc606_5 gpc8858 (
      {stage2_31[89], stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18]},
      {stage3_35[2],stage3_34[9],stage3_33[24],stage3_32[29],stage3_31[32]}
   );
   gpc606_5 gpc8859 (
      {stage2_31[95], stage2_31[96], stage2_31[97], stage2_31[98], stage2_31[99], stage2_31[100]},
      {stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24]},
      {stage3_35[3],stage3_34[10],stage3_33[25],stage3_32[30],stage3_31[33]}
   );
   gpc606_5 gpc8860 (
      {stage2_31[101], stage2_31[102], stage2_31[103], stage2_31[104], stage2_31[105], stage2_31[106]},
      {stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29], stage2_33[30]},
      {stage3_35[4],stage3_34[11],stage3_33[26],stage3_32[31],stage3_31[34]}
   );
   gpc606_5 gpc8861 (
      {stage2_31[107], stage2_31[108], stage2_31[109], stage2_31[110], stage2_31[111], stage2_31[112]},
      {stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35], stage2_33[36]},
      {stage3_35[5],stage3_34[12],stage3_33[27],stage3_32[32],stage3_31[35]}
   );
   gpc606_5 gpc8862 (
      {stage2_31[113], stage2_31[114], stage2_31[115], stage2_31[116], stage2_31[117], stage2_31[118]},
      {stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41], stage2_33[42]},
      {stage3_35[6],stage3_34[13],stage3_33[28],stage3_32[33],stage3_31[36]}
   );
   gpc615_5 gpc8863 (
      {stage2_31[119], stage2_31[120], stage2_31[121], stage2_31[122], stage2_31[123]},
      {stage2_32[42]},
      {stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48]},
      {stage3_35[7],stage3_34[14],stage3_33[29],stage3_32[34],stage3_31[37]}
   );
   gpc1163_5 gpc8864 (
      {stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54]},
      {stage2_34[0]},
      {stage2_35[0]},
      {stage3_36[0],stage3_35[8],stage3_34[15],stage3_33[30],stage3_32[35]}
   );
   gpc1163_5 gpc8865 (
      {stage2_32[46], stage2_32[47], stage2_32[48]},
      {stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59], stage2_33[60]},
      {stage2_34[1]},
      {stage2_35[1]},
      {stage3_36[1],stage3_35[9],stage3_34[16],stage3_33[31],stage3_32[36]}
   );
   gpc1163_5 gpc8866 (
      {stage2_32[49], stage2_32[50], stage2_32[51]},
      {stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65], stage2_33[66]},
      {stage2_34[2]},
      {stage2_35[2]},
      {stage3_36[2],stage3_35[10],stage3_34[17],stage3_33[32],stage3_32[37]}
   );
   gpc1163_5 gpc8867 (
      {stage2_32[52], stage2_32[53], stage2_32[54]},
      {stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71], stage2_33[72]},
      {stage2_34[3]},
      {stage2_35[3]},
      {stage3_36[3],stage3_35[11],stage3_34[18],stage3_33[33],stage3_32[38]}
   );
   gpc1163_5 gpc8868 (
      {stage2_32[55], stage2_32[56], stage2_32[57]},
      {stage2_33[73], stage2_33[74], stage2_33[75], stage2_33[76], stage2_33[77], stage2_33[78]},
      {stage2_34[4]},
      {stage2_35[4]},
      {stage3_36[4],stage3_35[12],stage3_34[19],stage3_33[34],stage3_32[39]}
   );
   gpc1163_5 gpc8869 (
      {stage2_32[58], stage2_32[59], stage2_32[60]},
      {stage2_33[79], stage2_33[80], stage2_33[81], stage2_33[82], stage2_33[83], stage2_33[84]},
      {stage2_34[5]},
      {stage2_35[5]},
      {stage3_36[5],stage3_35[13],stage3_34[20],stage3_33[35],stage3_32[40]}
   );
   gpc1163_5 gpc8870 (
      {stage2_32[61], stage2_32[62], stage2_32[63]},
      {stage2_33[85], stage2_33[86], stage2_33[87], stage2_33[88], stage2_33[89], stage2_33[90]},
      {stage2_34[6]},
      {stage2_35[6]},
      {stage3_36[6],stage3_35[14],stage3_34[21],stage3_33[36],stage3_32[41]}
   );
   gpc606_5 gpc8871 (
      {stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68], stage2_32[69]},
      {stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11], stage2_34[12]},
      {stage3_36[7],stage3_35[15],stage3_34[22],stage3_33[37],stage3_32[42]}
   );
   gpc606_5 gpc8872 (
      {stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74], stage2_32[75]},
      {stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17], stage2_34[18]},
      {stage3_36[8],stage3_35[16],stage3_34[23],stage3_33[38],stage3_32[43]}
   );
   gpc606_5 gpc8873 (
      {stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80], stage2_32[81]},
      {stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23], stage2_34[24]},
      {stage3_36[9],stage3_35[17],stage3_34[24],stage3_33[39],stage3_32[44]}
   );
   gpc606_5 gpc8874 (
      {stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86], stage2_32[87]},
      {stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29], stage2_34[30]},
      {stage3_36[10],stage3_35[18],stage3_34[25],stage3_33[40],stage3_32[45]}
   );
   gpc606_5 gpc8875 (
      {stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92], stage2_32[93]},
      {stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35], stage2_34[36]},
      {stage3_36[11],stage3_35[19],stage3_34[26],stage3_33[41],stage3_32[46]}
   );
   gpc606_5 gpc8876 (
      {stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98], stage2_32[99]},
      {stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41], stage2_34[42]},
      {stage3_36[12],stage3_35[20],stage3_34[27],stage3_33[42],stage3_32[47]}
   );
   gpc606_5 gpc8877 (
      {stage2_32[100], stage2_32[101], stage2_32[102], stage2_32[103], stage2_32[104], stage2_32[105]},
      {stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47], stage2_34[48]},
      {stage3_36[13],stage3_35[21],stage3_34[28],stage3_33[43],stage3_32[48]}
   );
   gpc606_5 gpc8878 (
      {stage2_32[106], stage2_32[107], stage2_32[108], stage2_32[109], stage2_32[110], stage2_32[111]},
      {stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53], stage2_34[54]},
      {stage3_36[14],stage3_35[22],stage3_34[29],stage3_33[44],stage3_32[49]}
   );
   gpc615_5 gpc8879 (
      {stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage2_35[7]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[15],stage3_35[23],stage3_34[30]}
   );
   gpc615_5 gpc8880 (
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64]},
      {stage2_35[8]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[1],stage3_36[16],stage3_35[24],stage3_34[31]}
   );
   gpc615_5 gpc8881 (
      {stage2_34[65], stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69]},
      {stage2_35[9]},
      {stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage3_38[2],stage3_37[2],stage3_36[17],stage3_35[25],stage3_34[32]}
   );
   gpc615_5 gpc8882 (
      {stage2_34[70], stage2_34[71], stage2_34[72], stage2_34[73], stage2_34[74]},
      {stage2_35[10]},
      {stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21], stage2_36[22], stage2_36[23]},
      {stage3_38[3],stage3_37[3],stage3_36[18],stage3_35[26],stage3_34[33]}
   );
   gpc615_5 gpc8883 (
      {stage2_34[75], stage2_34[76], stage2_34[77], stage2_34[78], stage2_34[79]},
      {stage2_35[11]},
      {stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27], stage2_36[28], stage2_36[29]},
      {stage3_38[4],stage3_37[4],stage3_36[19],stage3_35[27],stage3_34[34]}
   );
   gpc615_5 gpc8884 (
      {stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83], stage2_34[84]},
      {stage2_35[12]},
      {stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35]},
      {stage3_38[5],stage3_37[5],stage3_36[20],stage3_35[28],stage3_34[35]}
   );
   gpc615_5 gpc8885 (
      {stage2_34[85], stage2_34[86], stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[13]},
      {stage2_36[36], stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41]},
      {stage3_38[6],stage3_37[6],stage3_36[21],stage3_35[29],stage3_34[36]}
   );
   gpc615_5 gpc8886 (
      {stage2_34[90], stage2_34[91], stage2_34[92], stage2_34[93], stage2_34[94]},
      {stage2_35[14]},
      {stage2_36[42], stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47]},
      {stage3_38[7],stage3_37[7],stage3_36[22],stage3_35[30],stage3_34[37]}
   );
   gpc615_5 gpc8887 (
      {stage2_34[95], stage2_34[96], stage2_34[97], stage2_34[98], stage2_34[99]},
      {stage2_35[15]},
      {stage2_36[48], stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53]},
      {stage3_38[8],stage3_37[8],stage3_36[23],stage3_35[31],stage3_34[38]}
   );
   gpc615_5 gpc8888 (
      {stage2_34[100], stage2_34[101], stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[16]},
      {stage2_36[54], stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59]},
      {stage3_38[9],stage3_37[9],stage3_36[24],stage3_35[32],stage3_34[39]}
   );
   gpc615_5 gpc8889 (
      {stage2_34[105], stage2_34[106], stage2_34[107], stage2_34[108], stage2_34[109]},
      {stage2_35[17]},
      {stage2_36[60], stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65]},
      {stage3_38[10],stage3_37[10],stage3_36[25],stage3_35[33],stage3_34[40]}
   );
   gpc615_5 gpc8890 (
      {stage2_34[110], stage2_34[111], stage2_34[112], stage2_34[113], stage2_34[114]},
      {stage2_35[18]},
      {stage2_36[66], stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71]},
      {stage3_38[11],stage3_37[11],stage3_36[26],stage3_35[34],stage3_34[41]}
   );
   gpc615_5 gpc8891 (
      {stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118], stage2_34[119]},
      {stage2_35[19]},
      {stage2_36[72], stage2_36[73], stage2_36[74], stage2_36[75], stage2_36[76], stage2_36[77]},
      {stage3_38[12],stage3_37[12],stage3_36[27],stage3_35[35],stage3_34[42]}
   );
   gpc615_5 gpc8892 (
      {stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123], stage2_34[124]},
      {stage2_35[20]},
      {stage2_36[78], stage2_36[79], stage2_36[80], stage2_36[81], stage2_36[82], stage2_36[83]},
      {stage3_38[13],stage3_37[13],stage3_36[28],stage3_35[36],stage3_34[43]}
   );
   gpc615_5 gpc8893 (
      {stage2_34[125], stage2_34[126], stage2_34[127], 1'b0, 1'b0},
      {stage2_35[21]},
      {stage2_36[84], stage2_36[85], stage2_36[86], stage2_36[87], stage2_36[88], stage2_36[89]},
      {stage3_38[14],stage3_37[14],stage3_36[29],stage3_35[37],stage3_34[44]}
   );
   gpc606_5 gpc8894 (
      {stage2_35[22], stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[15],stage3_37[15],stage3_36[30],stage3_35[38]}
   );
   gpc615_5 gpc8895 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[90]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[16],stage3_37[16],stage3_36[31],stage3_35[39]}
   );
   gpc615_5 gpc8896 (
      {stage2_35[33], stage2_35[34], stage2_35[35], stage2_35[36], stage2_35[37]},
      {stage2_36[91]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[17],stage3_37[17],stage3_36[32],stage3_35[40]}
   );
   gpc615_5 gpc8897 (
      {stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41], stage2_35[42]},
      {stage2_36[92]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[18],stage3_37[18],stage3_36[33],stage3_35[41]}
   );
   gpc615_5 gpc8898 (
      {stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[93]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[19],stage3_37[19],stage3_36[34],stage3_35[42]}
   );
   gpc615_5 gpc8899 (
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52]},
      {stage2_36[94]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[20],stage3_37[20],stage3_36[35],stage3_35[43]}
   );
   gpc615_5 gpc8900 (
      {stage2_35[53], stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57]},
      {stage2_36[95]},
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage3_39[6],stage3_38[21],stage3_37[21],stage3_36[36],stage3_35[44]}
   );
   gpc615_5 gpc8901 (
      {stage2_35[58], stage2_35[59], stage2_35[60], stage2_35[61], stage2_35[62]},
      {stage2_36[96]},
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage3_39[7],stage3_38[22],stage3_37[22],stage3_36[37],stage3_35[45]}
   );
   gpc615_5 gpc8902 (
      {stage2_35[63], stage2_35[64], stage2_35[65], stage2_35[66], stage2_35[67]},
      {stage2_36[97]},
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage3_39[8],stage3_38[23],stage3_37[23],stage3_36[38],stage3_35[46]}
   );
   gpc615_5 gpc8903 (
      {stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71], stage2_35[72]},
      {stage2_36[98]},
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58], stage2_37[59]},
      {stage3_39[9],stage3_38[24],stage3_37[24],stage3_36[39],stage3_35[47]}
   );
   gpc615_5 gpc8904 (
      {stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[99]},
      {stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63], stage2_37[64], stage2_37[65]},
      {stage3_39[10],stage3_38[25],stage3_37[25],stage3_36[40],stage3_35[48]}
   );
   gpc615_5 gpc8905 (
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82]},
      {stage2_36[100]},
      {stage2_37[66], stage2_37[67], stage2_37[68], stage2_37[69], stage2_37[70], stage2_37[71]},
      {stage3_39[11],stage3_38[26],stage3_37[26],stage3_36[41],stage3_35[49]}
   );
   gpc615_5 gpc8906 (
      {stage2_35[83], stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87]},
      {stage2_36[101]},
      {stage2_37[72], stage2_37[73], stage2_37[74], stage2_37[75], stage2_37[76], stage2_37[77]},
      {stage3_39[12],stage3_38[27],stage3_37[27],stage3_36[42],stage3_35[50]}
   );
   gpc615_5 gpc8907 (
      {stage2_35[88], stage2_35[89], stage2_35[90], stage2_35[91], stage2_35[92]},
      {stage2_36[102]},
      {stage2_37[78], stage2_37[79], stage2_37[80], stage2_37[81], stage2_37[82], stage2_37[83]},
      {stage3_39[13],stage3_38[28],stage3_37[28],stage3_36[43],stage3_35[51]}
   );
   gpc615_5 gpc8908 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97]},
      {stage2_36[103]},
      {stage2_37[84], stage2_37[85], stage2_37[86], stage2_37[87], stage2_37[88], stage2_37[89]},
      {stage3_39[14],stage3_38[29],stage3_37[29],stage3_36[44],stage3_35[52]}
   );
   gpc615_5 gpc8909 (
      {stage2_35[98], stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102]},
      {stage2_36[104]},
      {stage2_37[90], stage2_37[91], stage2_37[92], stage2_37[93], stage2_37[94], stage2_37[95]},
      {stage3_39[15],stage3_38[30],stage3_37[30],stage3_36[45],stage3_35[53]}
   );
   gpc615_5 gpc8910 (
      {stage2_35[103], stage2_35[104], stage2_35[105], stage2_35[106], stage2_35[107]},
      {stage2_36[105]},
      {stage2_37[96], stage2_37[97], stage2_37[98], stage2_37[99], stage2_37[100], stage2_37[101]},
      {stage3_39[16],stage3_38[31],stage3_37[31],stage3_36[46],stage3_35[54]}
   );
   gpc615_5 gpc8911 (
      {stage2_35[108], stage2_35[109], stage2_35[110], stage2_35[111], stage2_35[112]},
      {stage2_36[106]},
      {stage2_37[102], stage2_37[103], stage2_37[104], stage2_37[105], stage2_37[106], stage2_37[107]},
      {stage3_39[17],stage3_38[32],stage3_37[32],stage3_36[47],stage3_35[55]}
   );
   gpc615_5 gpc8912 (
      {stage2_35[113], stage2_35[114], stage2_35[115], stage2_35[116], stage2_35[117]},
      {stage2_36[107]},
      {stage2_37[108], stage2_37[109], stage2_37[110], stage2_37[111], stage2_37[112], stage2_37[113]},
      {stage3_39[18],stage3_38[33],stage3_37[33],stage3_36[48],stage3_35[56]}
   );
   gpc606_5 gpc8913 (
      {stage2_36[108], stage2_36[109], stage2_36[110], stage2_36[111], stage2_36[112], stage2_36[113]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[19],stage3_38[34],stage3_37[34],stage3_36[49]}
   );
   gpc615_5 gpc8914 (
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10]},
      {stage2_39[0]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[1],stage3_39[20],stage3_38[35]}
   );
   gpc615_5 gpc8915 (
      {stage2_38[11], stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15]},
      {stage2_39[1]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[1],stage3_40[2],stage3_39[21],stage3_38[36]}
   );
   gpc615_5 gpc8916 (
      {stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_39[2]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[2],stage3_40[3],stage3_39[22],stage3_38[37]}
   );
   gpc615_5 gpc8917 (
      {stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage2_39[3]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[3],stage3_40[4],stage3_39[23],stage3_38[38]}
   );
   gpc615_5 gpc8918 (
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30]},
      {stage2_39[4]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[4],stage3_40[5],stage3_39[24],stage3_38[39]}
   );
   gpc615_5 gpc8919 (
      {stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage2_39[5]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[5],stage3_40[6],stage3_39[25],stage3_38[40]}
   );
   gpc615_5 gpc8920 (
      {stage2_38[36], stage2_38[37], stage2_38[38], stage2_38[39], stage2_38[40]},
      {stage2_39[6]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[6],stage3_40[7],stage3_39[26],stage3_38[41]}
   );
   gpc615_5 gpc8921 (
      {stage2_38[41], stage2_38[42], stage2_38[43], stage2_38[44], stage2_38[45]},
      {stage2_39[7]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[7],stage3_40[8],stage3_39[27],stage3_38[42]}
   );
   gpc615_5 gpc8922 (
      {stage2_38[46], stage2_38[47], stage2_38[48], stage2_38[49], stage2_38[50]},
      {stage2_39[8]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[8],stage3_40[9],stage3_39[28],stage3_38[43]}
   );
   gpc615_5 gpc8923 (
      {stage2_38[51], stage2_38[52], stage2_38[53], stage2_38[54], stage2_38[55]},
      {stage2_39[9]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[9],stage3_40[10],stage3_39[29],stage3_38[44]}
   );
   gpc615_5 gpc8924 (
      {stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59], stage2_38[60]},
      {stage2_39[10]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[10],stage3_40[11],stage3_39[30],stage3_38[45]}
   );
   gpc615_5 gpc8925 (
      {stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_39[11]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[11],stage3_40[12],stage3_39[31],stage3_38[46]}
   );
   gpc615_5 gpc8926 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70]},
      {stage2_39[12]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[12],stage3_40[13],stage3_39[32],stage3_38[47]}
   );
   gpc615_5 gpc8927 (
      {stage2_38[71], stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75]},
      {stage2_39[13]},
      {stage2_40[78], stage2_40[79], stage2_40[80], stage2_40[81], stage2_40[82], stage2_40[83]},
      {stage3_42[13],stage3_41[13],stage3_40[14],stage3_39[33],stage3_38[48]}
   );
   gpc615_5 gpc8928 (
      {stage2_38[76], stage2_38[77], stage2_38[78], stage2_38[79], stage2_38[80]},
      {stage2_39[14]},
      {stage2_40[84], stage2_40[85], stage2_40[86], stage2_40[87], stage2_40[88], stage2_40[89]},
      {stage3_42[14],stage3_41[14],stage3_40[15],stage3_39[34],stage3_38[49]}
   );
   gpc615_5 gpc8929 (
      {stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_40[90]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[15],stage3_41[15],stage3_40[16],stage3_39[35]}
   );
   gpc615_5 gpc8930 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24]},
      {stage2_40[91]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[16],stage3_41[16],stage3_40[17],stage3_39[36]}
   );
   gpc615_5 gpc8931 (
      {stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage2_40[92]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[17],stage3_41[17],stage3_40[18],stage3_39[37]}
   );
   gpc615_5 gpc8932 (
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34]},
      {stage2_40[93]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[18],stage3_41[18],stage3_40[19],stage3_39[38]}
   );
   gpc615_5 gpc8933 (
      {stage2_39[35], stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39]},
      {stage2_40[94]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[19],stage3_41[19],stage3_40[20],stage3_39[39]}
   );
   gpc615_5 gpc8934 (
      {stage2_39[40], stage2_39[41], stage2_39[42], stage2_39[43], stage2_39[44]},
      {stage2_40[95]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[20],stage3_41[20],stage3_40[21],stage3_39[40]}
   );
   gpc615_5 gpc8935 (
      {stage2_39[45], stage2_39[46], stage2_39[47], stage2_39[48], stage2_39[49]},
      {stage2_40[96]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[21],stage3_41[21],stage3_40[22],stage3_39[41]}
   );
   gpc615_5 gpc8936 (
      {stage2_39[50], stage2_39[51], stage2_39[52], stage2_39[53], stage2_39[54]},
      {stage2_40[97]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[22],stage3_41[22],stage3_40[23],stage3_39[42]}
   );
   gpc615_5 gpc8937 (
      {stage2_39[55], stage2_39[56], stage2_39[57], stage2_39[58], stage2_39[59]},
      {stage2_40[98]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[23],stage3_41[23],stage3_40[24],stage3_39[43]}
   );
   gpc615_5 gpc8938 (
      {stage2_39[60], stage2_39[61], stage2_39[62], stage2_39[63], stage2_39[64]},
      {stage2_40[99]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[24],stage3_41[24],stage3_40[25],stage3_39[44]}
   );
   gpc615_5 gpc8939 (
      {stage2_39[65], stage2_39[66], stage2_39[67], stage2_39[68], stage2_39[69]},
      {stage2_40[100]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[25],stage3_41[25],stage3_40[26],stage3_39[45]}
   );
   gpc615_5 gpc8940 (
      {stage2_39[70], stage2_39[71], stage2_39[72], stage2_39[73], stage2_39[74]},
      {stage2_40[101]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[26],stage3_41[26],stage3_40[27],stage3_39[46]}
   );
   gpc615_5 gpc8941 (
      {stage2_39[75], stage2_39[76], stage2_39[77], stage2_39[78], stage2_39[79]},
      {stage2_40[102]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[27],stage3_41[27],stage3_40[28],stage3_39[47]}
   );
   gpc615_5 gpc8942 (
      {stage2_39[80], stage2_39[81], stage2_39[82], stage2_39[83], stage2_39[84]},
      {stage2_40[103]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[28],stage3_41[28],stage3_40[29],stage3_39[48]}
   );
   gpc615_5 gpc8943 (
      {stage2_39[85], stage2_39[86], stage2_39[87], stage2_39[88], stage2_39[89]},
      {stage2_40[104]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[29],stage3_41[29],stage3_40[30],stage3_39[49]}
   );
   gpc615_5 gpc8944 (
      {stage2_39[90], stage2_39[91], stage2_39[92], stage2_39[93], stage2_39[94]},
      {stage2_40[105]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[30],stage3_41[30],stage3_40[31],stage3_39[50]}
   );
   gpc615_5 gpc8945 (
      {stage2_39[95], stage2_39[96], stage2_39[97], stage2_39[98], stage2_39[99]},
      {stage2_40[106]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[31],stage3_41[31],stage3_40[32],stage3_39[51]}
   );
   gpc606_5 gpc8946 (
      {stage2_40[107], stage2_40[108], stage2_40[109], stage2_40[110], stage2_40[111], stage2_40[112]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[32],stage3_41[32],stage3_40[33]}
   );
   gpc606_5 gpc8947 (
      {stage2_40[113], stage2_40[114], stage2_40[115], stage2_40[116], stage2_40[117], stage2_40[118]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[33],stage3_41[33],stage3_40[34]}
   );
   gpc606_5 gpc8948 (
      {stage2_40[119], stage2_40[120], stage2_40[121], stage2_40[122], stage2_40[123], stage2_40[124]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[19],stage3_42[34],stage3_41[34],stage3_40[35]}
   );
   gpc606_5 gpc8949 (
      {stage2_40[125], stage2_40[126], stage2_40[127], stage2_40[128], stage2_40[129], stage2_40[130]},
      {stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21], stage2_42[22], stage2_42[23]},
      {stage3_44[3],stage3_43[20],stage3_42[35],stage3_41[35],stage3_40[36]}
   );
   gpc615_5 gpc8950 (
      {stage2_42[24], stage2_42[25], stage2_42[26], stage2_42[27], stage2_42[28]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[21],stage3_42[36]}
   );
   gpc615_5 gpc8951 (
      {stage2_42[29], stage2_42[30], stage2_42[31], stage2_42[32], stage2_42[33]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[22],stage3_42[37]}
   );
   gpc615_5 gpc8952 (
      {stage2_42[34], stage2_42[35], stage2_42[36], stage2_42[37], stage2_42[38]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[6],stage3_43[23],stage3_42[38]}
   );
   gpc615_5 gpc8953 (
      {stage2_42[39], stage2_42[40], stage2_42[41], stage2_42[42], stage2_42[43]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[7],stage3_43[24],stage3_42[39]}
   );
   gpc615_5 gpc8954 (
      {stage2_42[44], stage2_42[45], stage2_42[46], stage2_42[47], stage2_42[48]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[8],stage3_43[25],stage3_42[40]}
   );
   gpc615_5 gpc8955 (
      {stage2_42[49], stage2_42[50], stage2_42[51], stage2_42[52], stage2_42[53]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[9],stage3_43[26],stage3_42[41]}
   );
   gpc615_5 gpc8956 (
      {stage2_42[54], stage2_42[55], stage2_42[56], stage2_42[57], stage2_42[58]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[10],stage3_43[27],stage3_42[42]}
   );
   gpc615_5 gpc8957 (
      {stage2_42[59], stage2_42[60], stage2_42[61], stage2_42[62], stage2_42[63]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[11],stage3_43[28],stage3_42[43]}
   );
   gpc615_5 gpc8958 (
      {stage2_42[64], stage2_42[65], stage2_42[66], stage2_42[67], stage2_42[68]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[12],stage3_43[29],stage3_42[44]}
   );
   gpc615_5 gpc8959 (
      {stage2_42[69], stage2_42[70], stage2_42[71], stage2_42[72], stage2_42[73]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[13],stage3_43[30],stage3_42[45]}
   );
   gpc606_5 gpc8960 (
      {stage2_43[10], stage2_43[11], stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[10],stage3_45[10],stage3_44[14],stage3_43[31]}
   );
   gpc606_5 gpc8961 (
      {stage2_43[16], stage2_43[17], stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[11],stage3_45[11],stage3_44[15],stage3_43[32]}
   );
   gpc606_5 gpc8962 (
      {stage2_43[22], stage2_43[23], stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[12],stage3_45[12],stage3_44[16],stage3_43[33]}
   );
   gpc606_5 gpc8963 (
      {stage2_43[28], stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[13],stage3_45[13],stage3_44[17],stage3_43[34]}
   );
   gpc606_5 gpc8964 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38], stage2_43[39]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[14],stage3_45[14],stage3_44[18],stage3_43[35]}
   );
   gpc606_5 gpc8965 (
      {stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[15],stage3_45[15],stage3_44[19],stage3_43[36]}
   );
   gpc606_5 gpc8966 (
      {stage2_43[46], stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[16],stage3_45[16],stage3_44[20],stage3_43[37]}
   );
   gpc606_5 gpc8967 (
      {stage2_43[52], stage2_43[53], stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[17],stage3_45[17],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc8968 (
      {stage2_43[58], stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62]},
      {stage2_44[60]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[18],stage3_45[18],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc8969 (
      {stage2_43[63], stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67]},
      {stage2_44[61]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[19],stage3_45[19],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc8970 (
      {stage2_43[68], stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72]},
      {stage2_44[62]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[20],stage3_45[20],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc8971 (
      {stage2_43[73], stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77]},
      {stage2_44[63]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[21],stage3_45[21],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc8972 (
      {stage2_43[78], stage2_43[79], stage2_43[80], stage2_43[81], stage2_43[82]},
      {stage2_44[64]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[22],stage3_45[22],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc8973 (
      {stage2_43[83], stage2_43[84], stage2_43[85], stage2_43[86], stage2_43[87]},
      {stage2_44[65]},
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage3_47[13],stage3_46[23],stage3_45[23],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc8974 (
      {stage2_43[88], stage2_43[89], stage2_43[90], stage2_43[91], stage2_43[92]},
      {stage2_44[66]},
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage3_47[14],stage3_46[24],stage3_45[24],stage3_44[28],stage3_43[45]}
   );
   gpc615_5 gpc8975 (
      {stage2_43[93], stage2_43[94], stage2_43[95], stage2_43[96], stage2_43[97]},
      {stage2_44[67]},
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage3_47[15],stage3_46[25],stage3_45[25],stage3_44[29],stage3_43[46]}
   );
   gpc606_5 gpc8976 (
      {stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71], stage2_44[72], stage2_44[73]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[16],stage3_46[26],stage3_45[26],stage3_44[30]}
   );
   gpc606_5 gpc8977 (
      {stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77], stage2_44[78], stage2_44[79]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[17],stage3_46[27],stage3_45[27],stage3_44[31]}
   );
   gpc606_5 gpc8978 (
      {stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83], stage2_44[84], stage2_44[85]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[18],stage3_46[28],stage3_45[28],stage3_44[32]}
   );
   gpc606_5 gpc8979 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[3],stage3_47[19],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc8980 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[4],stage3_47[20],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc8981 (
      {stage2_45[108], stage2_45[109], stage2_45[110], stage2_45[111], stage2_45[112], stage2_45[113]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[5],stage3_47[21],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc8982 (
      {stage2_45[114], stage2_45[115], stage2_45[116], stage2_45[117], stage2_45[118], stage2_45[119]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[6],stage3_47[22],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc8983 (
      {stage2_45[120], stage2_45[121], stage2_45[122], stage2_45[123], stage2_45[124], stage2_45[125]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[7],stage3_47[23],stage3_46[33],stage3_45[33]}
   );
   gpc615_5 gpc8984 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[30]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[5],stage3_48[8],stage3_47[24],stage3_46[34]}
   );
   gpc615_5 gpc8985 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[31]},
      {stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage3_50[1],stage3_49[6],stage3_48[9],stage3_47[25],stage3_46[35]}
   );
   gpc615_5 gpc8986 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[32]},
      {stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17]},
      {stage3_50[2],stage3_49[7],stage3_48[10],stage3_47[26],stage3_46[36]}
   );
   gpc615_5 gpc8987 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[33]},
      {stage2_48[18], stage2_48[19], stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23]},
      {stage3_50[3],stage3_49[8],stage3_48[11],stage3_47[27],stage3_46[37]}
   );
   gpc615_5 gpc8988 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[34]},
      {stage2_48[24], stage2_48[25], stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29]},
      {stage3_50[4],stage3_49[9],stage3_48[12],stage3_47[28],stage3_46[38]}
   );
   gpc615_5 gpc8989 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[35]},
      {stage2_48[30], stage2_48[31], stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35]},
      {stage3_50[5],stage3_49[10],stage3_48[13],stage3_47[29],stage3_46[39]}
   );
   gpc615_5 gpc8990 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[36]},
      {stage2_48[36], stage2_48[37], stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41]},
      {stage3_50[6],stage3_49[11],stage3_48[14],stage3_47[30],stage3_46[40]}
   );
   gpc615_5 gpc8991 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[37]},
      {stage2_48[42], stage2_48[43], stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47]},
      {stage3_50[7],stage3_49[12],stage3_48[15],stage3_47[31],stage3_46[41]}
   );
   gpc615_5 gpc8992 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[38]},
      {stage2_48[48], stage2_48[49], stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53]},
      {stage3_50[8],stage3_49[13],stage3_48[16],stage3_47[32],stage3_46[42]}
   );
   gpc615_5 gpc8993 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[39]},
      {stage2_48[54], stage2_48[55], stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59]},
      {stage3_50[9],stage3_49[14],stage3_48[17],stage3_47[33],stage3_46[43]}
   );
   gpc615_5 gpc8994 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[40]},
      {stage2_48[60], stage2_48[61], stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65]},
      {stage3_50[10],stage3_49[15],stage3_48[18],stage3_47[34],stage3_46[44]}
   );
   gpc615_5 gpc8995 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[41]},
      {stage2_48[66], stage2_48[67], stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71]},
      {stage3_50[11],stage3_49[16],stage3_48[19],stage3_47[35],stage3_46[45]}
   );
   gpc615_5 gpc8996 (
      {stage2_46[78], stage2_46[79], stage2_46[80], stage2_46[81], stage2_46[82]},
      {stage2_47[42]},
      {stage2_48[72], stage2_48[73], stage2_48[74], stage2_48[75], stage2_48[76], stage2_48[77]},
      {stage3_50[12],stage3_49[17],stage3_48[20],stage3_47[36],stage3_46[46]}
   );
   gpc615_5 gpc8997 (
      {stage2_46[83], stage2_46[84], stage2_46[85], stage2_46[86], stage2_46[87]},
      {stage2_47[43]},
      {stage2_48[78], stage2_48[79], stage2_48[80], stage2_48[81], stage2_48[82], stage2_48[83]},
      {stage3_50[13],stage3_49[18],stage3_48[21],stage3_47[37],stage3_46[47]}
   );
   gpc615_5 gpc8998 (
      {stage2_46[88], stage2_46[89], stage2_46[90], stage2_46[91], stage2_46[92]},
      {stage2_47[44]},
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage3_50[14],stage3_49[19],stage3_48[22],stage3_47[38],stage3_46[48]}
   );
   gpc1163_5 gpc8999 (
      {stage2_47[45], stage2_47[46], stage2_47[47]},
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_49[0]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[15],stage3_49[20],stage3_48[23],stage3_47[39]}
   );
   gpc1163_5 gpc9000 (
      {stage2_47[48], stage2_47[49], stage2_47[50]},
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_49[1]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[16],stage3_49[21],stage3_48[24],stage3_47[40]}
   );
   gpc1163_5 gpc9001 (
      {stage2_47[51], stage2_47[52], stage2_47[53]},
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_49[2]},
      {stage2_50[2]},
      {stage3_51[2],stage3_50[17],stage3_49[22],stage3_48[25],stage3_47[41]}
   );
   gpc1163_5 gpc9002 (
      {stage2_47[54], stage2_47[55], stage2_47[56]},
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_49[3]},
      {stage2_50[3]},
      {stage3_51[3],stage3_50[18],stage3_49[23],stage3_48[26],stage3_47[42]}
   );
   gpc1163_5 gpc9003 (
      {stage2_47[57], stage2_47[58], stage2_47[59]},
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_49[4]},
      {stage2_50[4]},
      {stage3_51[4],stage3_50[19],stage3_49[24],stage3_48[27],stage3_47[43]}
   );
   gpc1163_5 gpc9004 (
      {stage2_47[60], stage2_47[61], stage2_47[62]},
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_49[5]},
      {stage2_50[5]},
      {stage3_51[5],stage3_50[20],stage3_49[25],stage3_48[28],stage3_47[44]}
   );
   gpc615_5 gpc9005 (
      {stage2_47[63], stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67]},
      {stage2_48[126]},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[6],stage3_50[21],stage3_49[26],stage3_48[29],stage3_47[45]}
   );
   gpc615_5 gpc9006 (
      {stage2_47[68], stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72]},
      {stage2_48[127]},
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage3_51[7],stage3_50[22],stage3_49[27],stage3_48[30],stage3_47[46]}
   );
   gpc615_5 gpc9007 (
      {stage2_47[73], stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77]},
      {stage2_48[128]},
      {stage2_49[18], stage2_49[19], stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23]},
      {stage3_51[8],stage3_50[23],stage3_49[28],stage3_48[31],stage3_47[47]}
   );
   gpc615_5 gpc9008 (
      {stage2_47[78], stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82]},
      {stage2_48[129]},
      {stage2_49[24], stage2_49[25], stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29]},
      {stage3_51[9],stage3_50[24],stage3_49[29],stage3_48[32],stage3_47[48]}
   );
   gpc606_5 gpc9009 (
      {stage2_48[130], stage2_48[131], stage2_48[132], stage2_48[133], stage2_48[134], stage2_48[135]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[0],stage3_51[10],stage3_50[25],stage3_49[30],stage3_48[33]}
   );
   gpc606_5 gpc9010 (
      {stage2_48[136], stage2_48[137], stage2_48[138], stage2_48[139], stage2_48[140], stage2_48[141]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[1],stage3_51[11],stage3_50[26],stage3_49[31],stage3_48[34]}
   );
   gpc606_5 gpc9011 (
      {stage2_48[142], stage2_48[143], stage2_48[144], stage2_48[145], stage2_48[146], stage2_48[147]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[2],stage3_51[12],stage3_50[27],stage3_49[32],stage3_48[35]}
   );
   gpc606_5 gpc9012 (
      {stage2_48[148], stage2_48[149], stage2_48[150], stage2_48[151], stage2_48[152], stage2_48[153]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[3],stage3_51[13],stage3_50[28],stage3_49[33],stage3_48[36]}
   );
   gpc606_5 gpc9013 (
      {stage2_49[30], stage2_49[31], stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[4],stage3_51[14],stage3_50[29],stage3_49[34]}
   );
   gpc606_5 gpc9014 (
      {stage2_49[36], stage2_49[37], stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[5],stage3_51[15],stage3_50[30],stage3_49[35]}
   );
   gpc606_5 gpc9015 (
      {stage2_49[42], stage2_49[43], stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[6],stage3_51[16],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc9016 (
      {stage2_49[48], stage2_49[49], stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[7],stage3_51[17],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc9017 (
      {stage2_49[54], stage2_49[55], stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[8],stage3_51[18],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc9018 (
      {stage2_49[60], stage2_49[61], stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[9],stage3_51[19],stage3_50[34],stage3_49[39]}
   );
   gpc606_5 gpc9019 (
      {stage2_49[66], stage2_49[67], stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71]},
      {stage2_51[36], stage2_51[37], stage2_51[38], stage2_51[39], stage2_51[40], stage2_51[41]},
      {stage3_53[6],stage3_52[10],stage3_51[20],stage3_50[35],stage3_49[40]}
   );
   gpc606_5 gpc9020 (
      {stage2_49[72], stage2_49[73], stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77]},
      {stage2_51[42], stage2_51[43], stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47]},
      {stage3_53[7],stage3_52[11],stage3_51[21],stage3_50[36],stage3_49[41]}
   );
   gpc606_5 gpc9021 (
      {stage2_49[78], stage2_49[79], stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83]},
      {stage2_51[48], stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage3_53[8],stage3_52[12],stage3_51[22],stage3_50[37],stage3_49[42]}
   );
   gpc606_5 gpc9022 (
      {stage2_49[84], stage2_49[85], stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89]},
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58], stage2_51[59]},
      {stage3_53[9],stage3_52[13],stage3_51[23],stage3_50[38],stage3_49[43]}
   );
   gpc606_5 gpc9023 (
      {stage2_49[90], stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_51[60], stage2_51[61], stage2_51[62], stage2_51[63], stage2_51[64], stage2_51[65]},
      {stage3_53[10],stage3_52[14],stage3_51[24],stage3_50[39],stage3_49[44]}
   );
   gpc2135_5 gpc9024 (
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34]},
      {stage2_51[66], stage2_51[67], stage2_51[68]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[11],stage3_52[15],stage3_51[25],stage3_50[40]}
   );
   gpc1406_5 gpc9025 (
      {stage2_50[35], stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40]},
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4]},
      {stage2_53[2]},
      {stage3_54[1],stage3_53[12],stage3_52[16],stage3_51[26],stage3_50[41]}
   );
   gpc1406_5 gpc9026 (
      {stage2_50[41], stage2_50[42], stage2_50[43], stage2_50[44], stage2_50[45], stage2_50[46]},
      {stage2_52[5], stage2_52[6], stage2_52[7], stage2_52[8]},
      {stage2_53[3]},
      {stage3_54[2],stage3_53[13],stage3_52[17],stage3_51[27],stage3_50[42]}
   );
   gpc1406_5 gpc9027 (
      {stage2_50[47], stage2_50[48], stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52]},
      {stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12]},
      {stage2_53[4]},
      {stage3_54[3],stage3_53[14],stage3_52[18],stage3_51[28],stage3_50[43]}
   );
   gpc606_5 gpc9028 (
      {stage2_50[53], stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17], stage2_52[18]},
      {stage3_54[4],stage3_53[15],stage3_52[19],stage3_51[29],stage3_50[44]}
   );
   gpc606_5 gpc9029 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63], stage2_50[64]},
      {stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23], stage2_52[24]},
      {stage3_54[5],stage3_53[16],stage3_52[20],stage3_51[30],stage3_50[45]}
   );
   gpc606_5 gpc9030 (
      {stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68], stage2_50[69], stage2_50[70]},
      {stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29], stage2_52[30]},
      {stage3_54[6],stage3_53[17],stage3_52[21],stage3_51[31],stage3_50[46]}
   );
   gpc606_5 gpc9031 (
      {stage2_50[71], stage2_50[72], stage2_50[73], stage2_50[74], stage2_50[75], stage2_50[76]},
      {stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35], stage2_52[36]},
      {stage3_54[7],stage3_53[18],stage3_52[22],stage3_51[32],stage3_50[47]}
   );
   gpc606_5 gpc9032 (
      {stage2_50[77], stage2_50[78], stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82]},
      {stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41], stage2_52[42]},
      {stage3_54[8],stage3_53[19],stage3_52[23],stage3_51[33],stage3_50[48]}
   );
   gpc606_5 gpc9033 (
      {stage2_50[83], stage2_50[84], stage2_50[85], stage2_50[86], stage2_50[87], stage2_50[88]},
      {stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47], stage2_52[48]},
      {stage3_54[9],stage3_53[20],stage3_52[24],stage3_51[34],stage3_50[49]}
   );
   gpc606_5 gpc9034 (
      {stage2_50[89], stage2_50[90], stage2_50[91], stage2_50[92], stage2_50[93], stage2_50[94]},
      {stage2_52[49], stage2_52[50], stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54]},
      {stage3_54[10],stage3_53[21],stage3_52[25],stage3_51[35],stage3_50[50]}
   );
   gpc606_5 gpc9035 (
      {stage2_50[95], stage2_50[96], stage2_50[97], stage2_50[98], stage2_50[99], stage2_50[100]},
      {stage2_52[55], stage2_52[56], stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60]},
      {stage3_54[11],stage3_53[22],stage3_52[26],stage3_51[36],stage3_50[51]}
   );
   gpc606_5 gpc9036 (
      {stage2_50[101], stage2_50[102], stage2_50[103], stage2_50[104], stage2_50[105], stage2_50[106]},
      {stage2_52[61], stage2_52[62], stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66]},
      {stage3_54[12],stage3_53[23],stage3_52[27],stage3_51[37],stage3_50[52]}
   );
   gpc606_5 gpc9037 (
      {stage2_50[107], stage2_50[108], stage2_50[109], stage2_50[110], stage2_50[111], stage2_50[112]},
      {stage2_52[67], stage2_52[68], stage2_52[69], stage2_52[70], stage2_52[71], stage2_52[72]},
      {stage3_54[13],stage3_53[24],stage3_52[28],stage3_51[38],stage3_50[53]}
   );
   gpc606_5 gpc9038 (
      {stage2_50[113], stage2_50[114], stage2_50[115], stage2_50[116], stage2_50[117], stage2_50[118]},
      {stage2_52[73], stage2_52[74], stage2_52[75], stage2_52[76], stage2_52[77], stage2_52[78]},
      {stage3_54[14],stage3_53[25],stage3_52[29],stage3_51[39],stage3_50[54]}
   );
   gpc606_5 gpc9039 (
      {stage2_50[119], stage2_50[120], stage2_50[121], stage2_50[122], stage2_50[123], stage2_50[124]},
      {stage2_52[79], stage2_52[80], stage2_52[81], stage2_52[82], stage2_52[83], stage2_52[84]},
      {stage3_54[15],stage3_53[26],stage3_52[30],stage3_51[40],stage3_50[55]}
   );
   gpc606_5 gpc9040 (
      {stage2_50[125], stage2_50[126], stage2_50[127], stage2_50[128], stage2_50[129], stage2_50[130]},
      {stage2_52[85], stage2_52[86], stage2_52[87], stage2_52[88], stage2_52[89], stage2_52[90]},
      {stage3_54[16],stage3_53[27],stage3_52[31],stage3_51[41],stage3_50[56]}
   );
   gpc606_5 gpc9041 (
      {stage2_50[131], stage2_50[132], stage2_50[133], stage2_50[134], stage2_50[135], stage2_50[136]},
      {stage2_52[91], stage2_52[92], stage2_52[93], stage2_52[94], stage2_52[95], stage2_52[96]},
      {stage3_54[17],stage3_53[28],stage3_52[32],stage3_51[42],stage3_50[57]}
   );
   gpc606_5 gpc9042 (
      {stage2_50[137], stage2_50[138], stage2_50[139], stage2_50[140], stage2_50[141], stage2_50[142]},
      {stage2_52[97], stage2_52[98], stage2_52[99], stage2_52[100], stage2_52[101], stage2_52[102]},
      {stage3_54[18],stage3_53[29],stage3_52[33],stage3_51[43],stage3_50[58]}
   );
   gpc606_5 gpc9043 (
      {stage2_50[143], stage2_50[144], stage2_50[145], stage2_50[146], stage2_50[147], stage2_50[148]},
      {stage2_52[103], stage2_52[104], stage2_52[105], stage2_52[106], stage2_52[107], stage2_52[108]},
      {stage3_54[19],stage3_53[30],stage3_52[34],stage3_51[44],stage3_50[59]}
   );
   gpc606_5 gpc9044 (
      {stage2_51[69], stage2_51[70], stage2_51[71], stage2_51[72], stage2_51[73], stage2_51[74]},
      {stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10]},
      {stage3_55[0],stage3_54[20],stage3_53[31],stage3_52[35],stage3_51[45]}
   );
   gpc606_5 gpc9045 (
      {stage2_51[75], stage2_51[76], stage2_51[77], stage2_51[78], stage2_51[79], stage2_51[80]},
      {stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16]},
      {stage3_55[1],stage3_54[21],stage3_53[32],stage3_52[36],stage3_51[46]}
   );
   gpc606_5 gpc9046 (
      {stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[2],stage3_54[22],stage3_53[33]}
   );
   gpc606_5 gpc9047 (
      {stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[3],stage3_54[23],stage3_53[34]}
   );
   gpc606_5 gpc9048 (
      {stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[4],stage3_54[24],stage3_53[35]}
   );
   gpc606_5 gpc9049 (
      {stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[3],stage3_55[5],stage3_54[25],stage3_53[36]}
   );
   gpc606_5 gpc9050 (
      {stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[4],stage3_55[6],stage3_54[26],stage3_53[37]}
   );
   gpc606_5 gpc9051 (
      {stage2_53[47], stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[5],stage3_55[7],stage3_54[27],stage3_53[38]}
   );
   gpc606_5 gpc9052 (
      {stage2_53[53], stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[6],stage3_55[8],stage3_54[28],stage3_53[39]}
   );
   gpc606_5 gpc9053 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63], stage2_53[64]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[7],stage3_55[9],stage3_54[29],stage3_53[40]}
   );
   gpc606_5 gpc9054 (
      {stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68], stage2_53[69], stage2_53[70]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[8],stage3_55[10],stage3_54[30],stage3_53[41]}
   );
   gpc606_5 gpc9055 (
      {stage2_53[71], stage2_53[72], stage2_53[73], stage2_53[74], stage2_53[75], stage2_53[76]},
      {stage2_55[54], stage2_55[55], stage2_55[56], stage2_55[57], stage2_55[58], stage2_55[59]},
      {stage3_57[9],stage3_56[9],stage3_55[11],stage3_54[31],stage3_53[42]}
   );
   gpc606_5 gpc9056 (
      {stage2_53[77], stage2_53[78], stage2_53[79], stage2_53[80], stage2_53[81], stage2_53[82]},
      {stage2_55[60], stage2_55[61], stage2_55[62], stage2_55[63], stage2_55[64], stage2_55[65]},
      {stage3_57[10],stage3_56[10],stage3_55[12],stage3_54[32],stage3_53[43]}
   );
   gpc606_5 gpc9057 (
      {stage2_53[83], stage2_53[84], stage2_53[85], stage2_53[86], stage2_53[87], stage2_53[88]},
      {stage2_55[66], stage2_55[67], stage2_55[68], stage2_55[69], stage2_55[70], stage2_55[71]},
      {stage3_57[11],stage3_56[11],stage3_55[13],stage3_54[33],stage3_53[44]}
   );
   gpc606_5 gpc9058 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[12],stage3_56[12],stage3_55[14],stage3_54[34]}
   );
   gpc606_5 gpc9059 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[13],stage3_56[13],stage3_55[15],stage3_54[35]}
   );
   gpc606_5 gpc9060 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[14],stage3_56[14],stage3_55[16],stage3_54[36]}
   );
   gpc606_5 gpc9061 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22], stage2_54[23]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[15],stage3_56[15],stage3_55[17],stage3_54[37]}
   );
   gpc606_5 gpc9062 (
      {stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[16],stage3_56[16],stage3_55[18],stage3_54[38]}
   );
   gpc606_5 gpc9063 (
      {stage2_54[30], stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[17],stage3_56[17],stage3_55[19],stage3_54[39]}
   );
   gpc606_5 gpc9064 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40], stage2_54[41]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[18],stage3_56[18],stage3_55[20],stage3_54[40]}
   );
   gpc606_5 gpc9065 (
      {stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45], stage2_54[46], stage2_54[47]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[19],stage3_56[19],stage3_55[21],stage3_54[41]}
   );
   gpc606_5 gpc9066 (
      {stage2_54[48], stage2_54[49], stage2_54[50], stage2_54[51], stage2_54[52], stage2_54[53]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[20],stage3_56[20],stage3_55[22],stage3_54[42]}
   );
   gpc606_5 gpc9067 (
      {stage2_54[54], stage2_54[55], stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[21],stage3_56[21],stage3_55[23],stage3_54[43]}
   );
   gpc606_5 gpc9068 (
      {stage2_54[60], stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[22],stage3_56[22],stage3_55[24],stage3_54[44]}
   );
   gpc606_5 gpc9069 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70], stage2_54[71]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[23],stage3_56[23],stage3_55[25],stage3_54[45]}
   );
   gpc606_5 gpc9070 (
      {stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75], stage2_54[76], stage2_54[77]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[24],stage3_56[24],stage3_55[26],stage3_54[46]}
   );
   gpc606_5 gpc9071 (
      {stage2_54[78], stage2_54[79], stage2_54[80], stage2_54[81], stage2_54[82], stage2_54[83]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[25],stage3_56[25],stage3_55[27],stage3_54[47]}
   );
   gpc606_5 gpc9072 (
      {stage2_54[84], stage2_54[85], stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[26],stage3_56[26],stage3_55[28],stage3_54[48]}
   );
   gpc606_5 gpc9073 (
      {stage2_54[90], stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[27],stage3_56[27],stage3_55[29],stage3_54[49]}
   );
   gpc606_5 gpc9074 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], stage2_54[100], stage2_54[101]},
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100], stage2_56[101]},
      {stage3_58[16],stage3_57[28],stage3_56[28],stage3_55[30],stage3_54[50]}
   );
   gpc606_5 gpc9075 (
      {stage2_54[102], stage2_54[103], stage2_54[104], stage2_54[105], stage2_54[106], stage2_54[107]},
      {stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105], stage2_56[106], stage2_56[107]},
      {stage3_58[17],stage3_57[29],stage3_56[29],stage3_55[31],stage3_54[51]}
   );
   gpc606_5 gpc9076 (
      {stage2_54[108], stage2_54[109], stage2_54[110], stage2_54[111], stage2_54[112], stage2_54[113]},
      {stage2_56[108], stage2_56[109], stage2_56[110], stage2_56[111], stage2_56[112], stage2_56[113]},
      {stage3_58[18],stage3_57[30],stage3_56[30],stage3_55[32],stage3_54[52]}
   );
   gpc606_5 gpc9077 (
      {stage2_55[72], stage2_55[73], stage2_55[74], stage2_55[75], stage2_55[76], stage2_55[77]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[19],stage3_57[31],stage3_56[31],stage3_55[33]}
   );
   gpc606_5 gpc9078 (
      {stage2_55[78], stage2_55[79], stage2_55[80], stage2_55[81], stage2_55[82], stage2_55[83]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[20],stage3_57[32],stage3_56[32],stage3_55[34]}
   );
   gpc606_5 gpc9079 (
      {stage2_55[84], stage2_55[85], stage2_55[86], stage2_55[87], stage2_55[88], stage2_55[89]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[21],stage3_57[33],stage3_56[33],stage3_55[35]}
   );
   gpc606_5 gpc9080 (
      {stage2_55[90], stage2_55[91], stage2_55[92], stage2_55[93], stage2_55[94], stage2_55[95]},
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage3_59[3],stage3_58[22],stage3_57[34],stage3_56[34],stage3_55[36]}
   );
   gpc606_5 gpc9081 (
      {stage2_55[96], stage2_55[97], stage2_55[98], stage2_55[99], stage2_55[100], stage2_55[101]},
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage3_59[4],stage3_58[23],stage3_57[35],stage3_56[35],stage3_55[37]}
   );
   gpc606_5 gpc9082 (
      {stage2_56[114], stage2_56[115], stage2_56[116], stage2_56[117], stage2_56[118], stage2_56[119]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[5],stage3_58[24],stage3_57[36],stage3_56[36]}
   );
   gpc606_5 gpc9083 (
      {stage2_56[120], stage2_56[121], stage2_56[122], stage2_56[123], stage2_56[124], stage2_56[125]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[6],stage3_58[25],stage3_57[37],stage3_56[37]}
   );
   gpc606_5 gpc9084 (
      {stage2_56[126], stage2_56[127], stage2_56[128], stage2_56[129], stage2_56[130], stage2_56[131]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[7],stage3_58[26],stage3_57[38],stage3_56[38]}
   );
   gpc606_5 gpc9085 (
      {stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33], stage2_57[34], stage2_57[35]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[3],stage3_59[8],stage3_58[27],stage3_57[39]}
   );
   gpc606_5 gpc9086 (
      {stage2_57[36], stage2_57[37], stage2_57[38], stage2_57[39], stage2_57[40], stage2_57[41]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[4],stage3_59[9],stage3_58[28],stage3_57[40]}
   );
   gpc606_5 gpc9087 (
      {stage2_57[42], stage2_57[43], stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[5],stage3_59[10],stage3_58[29],stage3_57[41]}
   );
   gpc606_5 gpc9088 (
      {stage2_57[48], stage2_57[49], stage2_57[50], stage2_57[51], stage2_57[52], stage2_57[53]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[6],stage3_59[11],stage3_58[30],stage3_57[42]}
   );
   gpc606_5 gpc9089 (
      {stage2_57[54], stage2_57[55], stage2_57[56], stage2_57[57], stage2_57[58], stage2_57[59]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[7],stage3_59[12],stage3_58[31],stage3_57[43]}
   );
   gpc606_5 gpc9090 (
      {stage2_57[60], stage2_57[61], stage2_57[62], stage2_57[63], stage2_57[64], stage2_57[65]},
      {stage2_59[30], stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35]},
      {stage3_61[5],stage3_60[8],stage3_59[13],stage3_58[32],stage3_57[44]}
   );
   gpc606_5 gpc9091 (
      {stage2_57[66], stage2_57[67], stage2_57[68], stage2_57[69], stage2_57[70], stage2_57[71]},
      {stage2_59[36], stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41]},
      {stage3_61[6],stage3_60[9],stage3_59[14],stage3_58[33],stage3_57[45]}
   );
   gpc207_4 gpc9092 (
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23], stage2_58[24]},
      {stage2_60[0], stage2_60[1]},
      {stage3_61[7],stage3_60[10],stage3_59[15],stage3_58[34]}
   );
   gpc207_4 gpc9093 (
      {stage2_58[25], stage2_58[26], stage2_58[27], stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31]},
      {stage2_60[2], stage2_60[3]},
      {stage3_61[8],stage3_60[11],stage3_59[16],stage3_58[35]}
   );
   gpc207_4 gpc9094 (
      {stage2_58[32], stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37], stage2_58[38]},
      {stage2_60[4], stage2_60[5]},
      {stage3_61[9],stage3_60[12],stage3_59[17],stage3_58[36]}
   );
   gpc207_4 gpc9095 (
      {stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42], stage2_58[43], stage2_58[44], stage2_58[45]},
      {stage2_60[6], stage2_60[7]},
      {stage3_61[10],stage3_60[13],stage3_59[18],stage3_58[37]}
   );
   gpc207_4 gpc9096 (
      {stage2_58[46], stage2_58[47], stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_60[8], stage2_60[9]},
      {stage3_61[11],stage3_60[14],stage3_59[19],stage3_58[38]}
   );
   gpc207_4 gpc9097 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57], stage2_58[58], stage2_58[59]},
      {stage2_60[10], stage2_60[11]},
      {stage3_61[12],stage3_60[15],stage3_59[20],stage3_58[39]}
   );
   gpc207_4 gpc9098 (
      {stage2_58[60], stage2_58[61], stage2_58[62], stage2_58[63], stage2_58[64], stage2_58[65], stage2_58[66]},
      {stage2_60[12], stage2_60[13]},
      {stage3_61[13],stage3_60[16],stage3_59[21],stage3_58[40]}
   );
   gpc207_4 gpc9099 (
      {stage2_58[67], stage2_58[68], stage2_58[69], stage2_58[70], stage2_58[71], stage2_58[72], stage2_58[73]},
      {stage2_60[14], stage2_60[15]},
      {stage3_61[14],stage3_60[17],stage3_59[22],stage3_58[41]}
   );
   gpc615_5 gpc9100 (
      {stage2_58[74], stage2_58[75], stage2_58[76], stage2_58[77], stage2_58[78]},
      {stage2_59[42]},
      {stage2_60[16], stage2_60[17], stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21]},
      {stage3_62[0],stage3_61[15],stage3_60[18],stage3_59[23],stage3_58[42]}
   );
   gpc606_5 gpc9101 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[1],stage3_61[16],stage3_60[19],stage3_59[24]}
   );
   gpc606_5 gpc9102 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[2],stage3_61[17],stage3_60[20],stage3_59[25]}
   );
   gpc606_5 gpc9103 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59], stage2_59[60]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[3],stage3_61[18],stage3_60[21],stage3_59[26]}
   );
   gpc606_5 gpc9104 (
      {stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64], stage2_59[65], stage2_59[66]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[4],stage3_61[19],stage3_60[22],stage3_59[27]}
   );
   gpc606_5 gpc9105 (
      {stage2_59[67], stage2_59[68], stage2_59[69], stage2_59[70], stage2_59[71], stage2_59[72]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[5],stage3_61[20],stage3_60[23],stage3_59[28]}
   );
   gpc606_5 gpc9106 (
      {stage2_59[73], stage2_59[74], stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[6],stage3_61[21],stage3_60[24],stage3_59[29]}
   );
   gpc606_5 gpc9107 (
      {stage2_59[79], stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[7],stage3_61[22],stage3_60[25],stage3_59[30]}
   );
   gpc606_5 gpc9108 (
      {stage2_59[85], stage2_59[86], stage2_59[87], stage2_59[88], stage2_59[89], stage2_59[90]},
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage3_63[7],stage3_62[8],stage3_61[23],stage3_60[26],stage3_59[31]}
   );
   gpc606_5 gpc9109 (
      {stage2_59[91], stage2_59[92], stage2_59[93], stage2_59[94], stage2_59[95], stage2_59[96]},
      {stage2_61[48], stage2_61[49], stage2_61[50], stage2_61[51], stage2_61[52], stage2_61[53]},
      {stage3_63[8],stage3_62[9],stage3_61[24],stage3_60[27],stage3_59[32]}
   );
   gpc606_5 gpc9110 (
      {stage2_59[97], stage2_59[98], stage2_59[99], stage2_59[100], stage2_59[101], stage2_59[102]},
      {stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58], stage2_61[59]},
      {stage3_63[9],stage3_62[10],stage3_61[25],stage3_60[28],stage3_59[33]}
   );
   gpc606_5 gpc9111 (
      {stage2_59[103], stage2_59[104], stage2_59[105], stage2_59[106], stage2_59[107], stage2_59[108]},
      {stage2_61[60], stage2_61[61], stage2_61[62], stage2_61[63], stage2_61[64], stage2_61[65]},
      {stage3_63[10],stage3_62[11],stage3_61[26],stage3_60[29],stage3_59[34]}
   );
   gpc606_5 gpc9112 (
      {stage2_59[109], stage2_59[110], stage2_59[111], stage2_59[112], stage2_59[113], stage2_59[114]},
      {stage2_61[66], stage2_61[67], stage2_61[68], stage2_61[69], stage2_61[70], stage2_61[71]},
      {stage3_63[11],stage3_62[12],stage3_61[27],stage3_60[30],stage3_59[35]}
   );
   gpc606_5 gpc9113 (
      {stage2_59[115], stage2_59[116], stage2_59[117], stage2_59[118], stage2_59[119], stage2_59[120]},
      {stage2_61[72], stage2_61[73], stage2_61[74], stage2_61[75], stage2_61[76], stage2_61[77]},
      {stage3_63[12],stage3_62[13],stage3_61[28],stage3_60[31],stage3_59[36]}
   );
   gpc606_5 gpc9114 (
      {stage2_59[121], stage2_59[122], stage2_59[123], stage2_59[124], stage2_59[125], stage2_59[126]},
      {stage2_61[78], stage2_61[79], stage2_61[80], stage2_61[81], stage2_61[82], stage2_61[83]},
      {stage3_63[13],stage3_62[14],stage3_61[29],stage3_60[32],stage3_59[37]}
   );
   gpc606_5 gpc9115 (
      {stage2_59[127], stage2_59[128], stage2_59[129], stage2_59[130], stage2_59[131], stage2_59[132]},
      {stage2_61[84], stage2_61[85], stage2_61[86], stage2_61[87], stage2_61[88], stage2_61[89]},
      {stage3_63[14],stage3_62[15],stage3_61[30],stage3_60[33],stage3_59[38]}
   );
   gpc606_5 gpc9116 (
      {stage2_60[22], stage2_60[23], stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[15],stage3_62[16],stage3_61[31],stage3_60[34]}
   );
   gpc606_5 gpc9117 (
      {stage2_60[28], stage2_60[29], stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[16],stage3_62[17],stage3_61[32],stage3_60[35]}
   );
   gpc606_5 gpc9118 (
      {stage2_60[34], stage2_60[35], stage2_60[36], stage2_60[37], stage2_60[38], stage2_60[39]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[17],stage3_62[18],stage3_61[33],stage3_60[36]}
   );
   gpc606_5 gpc9119 (
      {stage2_60[40], stage2_60[41], stage2_60[42], stage2_60[43], stage2_60[44], stage2_60[45]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[18],stage3_62[19],stage3_61[34],stage3_60[37]}
   );
   gpc606_5 gpc9120 (
      {stage2_60[46], stage2_60[47], stage2_60[48], stage2_60[49], stage2_60[50], stage2_60[51]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[19],stage3_62[20],stage3_61[35],stage3_60[38]}
   );
   gpc606_5 gpc9121 (
      {stage2_60[52], stage2_60[53], stage2_60[54], stage2_60[55], stage2_60[56], stage2_60[57]},
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34], stage2_62[35]},
      {stage3_64[5],stage3_63[20],stage3_62[21],stage3_61[36],stage3_60[39]}
   );
   gpc606_5 gpc9122 (
      {stage2_60[58], stage2_60[59], stage2_60[60], stage2_60[61], stage2_60[62], stage2_60[63]},
      {stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39], stage2_62[40], stage2_62[41]},
      {stage3_64[6],stage3_63[21],stage3_62[22],stage3_61[37],stage3_60[40]}
   );
   gpc606_5 gpc9123 (
      {stage2_60[64], stage2_60[65], stage2_60[66], stage2_60[67], stage2_60[68], stage2_60[69]},
      {stage2_62[42], stage2_62[43], stage2_62[44], stage2_62[45], stage2_62[46], stage2_62[47]},
      {stage3_64[7],stage3_63[22],stage3_62[23],stage3_61[38],stage3_60[41]}
   );
   gpc606_5 gpc9124 (
      {stage2_60[70], stage2_60[71], stage2_60[72], stage2_60[73], stage2_60[74], stage2_60[75]},
      {stage2_62[48], stage2_62[49], stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53]},
      {stage3_64[8],stage3_63[23],stage3_62[24],stage3_61[39],stage3_60[42]}
   );
   gpc606_5 gpc9125 (
      {stage2_60[76], stage2_60[77], stage2_60[78], stage2_60[79], stage2_60[80], stage2_60[81]},
      {stage2_62[54], stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage3_64[9],stage3_63[24],stage3_62[25],stage3_61[40],stage3_60[43]}
   );
   gpc606_5 gpc9126 (
      {stage2_60[82], stage2_60[83], stage2_60[84], stage2_60[85], stage2_60[86], stage2_60[87]},
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64], stage2_62[65]},
      {stage3_64[10],stage3_63[25],stage3_62[26],stage3_61[41],stage3_60[44]}
   );
   gpc606_5 gpc9127 (
      {stage2_60[88], stage2_60[89], stage2_60[90], stage2_60[91], stage2_60[92], stage2_60[93]},
      {stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69], stage2_62[70], stage2_62[71]},
      {stage3_64[11],stage3_63[26],stage3_62[27],stage3_61[42],stage3_60[45]}
   );
   gpc606_5 gpc9128 (
      {stage2_60[94], stage2_60[95], stage2_60[96], stage2_60[97], stage2_60[98], stage2_60[99]},
      {stage2_62[72], stage2_62[73], stage2_62[74], stage2_62[75], stage2_62[76], stage2_62[77]},
      {stage3_64[12],stage3_63[27],stage3_62[28],stage3_61[43],stage3_60[46]}
   );
   gpc606_5 gpc9129 (
      {stage2_60[100], stage2_60[101], stage2_60[102], stage2_60[103], stage2_60[104], stage2_60[105]},
      {stage2_62[78], stage2_62[79], stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83]},
      {stage3_64[13],stage3_63[28],stage3_62[29],stage3_61[44],stage3_60[47]}
   );
   gpc606_5 gpc9130 (
      {stage2_62[84], stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[0],stage3_64[14],stage3_63[29],stage3_62[30]}
   );
   gpc606_5 gpc9131 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94], stage2_62[95]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[1],stage3_64[15],stage3_63[30],stage3_62[31]}
   );
   gpc606_5 gpc9132 (
      {stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99], stage2_62[100], stage2_62[101]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[2],stage3_64[16],stage3_63[31],stage3_62[32]}
   );
   gpc606_5 gpc9133 (
      {stage2_62[102], stage2_62[103], stage2_62[104], stage2_62[105], stage2_62[106], stage2_62[107]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[3],stage3_64[17],stage3_63[32],stage3_62[33]}
   );
   gpc606_5 gpc9134 (
      {stage2_62[108], stage2_62[109], stage2_62[110], stage2_62[111], stage2_62[112], stage2_62[113]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[4],stage3_64[18],stage3_63[33],stage3_62[34]}
   );
   gpc606_5 gpc9135 (
      {stage2_62[114], stage2_62[115], stage2_62[116], stage2_62[117], stage2_62[118], stage2_62[119]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[5],stage3_64[19],stage3_63[34],stage3_62[35]}
   );
   gpc606_5 gpc9136 (
      {stage2_62[120], stage2_62[121], stage2_62[122], stage2_62[123], stage2_62[124], stage2_62[125]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[6],stage3_64[20],stage3_63[35],stage3_62[36]}
   );
   gpc606_5 gpc9137 (
      {stage2_62[126], stage2_62[127], stage2_62[128], stage2_62[129], stage2_62[130], stage2_62[131]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[7],stage3_64[21],stage3_63[36],stage3_62[37]}
   );
   gpc606_5 gpc9138 (
      {stage2_62[132], stage2_62[133], stage2_62[134], stage2_62[135], stage2_62[136], stage2_62[137]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[8],stage3_64[22],stage3_63[37],stage3_62[38]}
   );
   gpc606_5 gpc9139 (
      {stage2_62[138], stage2_62[139], stage2_62[140], stage2_62[141], stage2_62[142], stage2_62[143]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[9],stage3_64[23],stage3_63[38],stage3_62[39]}
   );
   gpc117_4 gpc9140 (
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage2_64[60]},
      {stage2_65[0]},
      {stage3_66[10],stage3_65[10],stage3_64[24],stage3_63[39]}
   );
   gpc117_4 gpc9141 (
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12], stage2_63[13]},
      {stage2_64[61]},
      {stage2_65[1]},
      {stage3_66[11],stage3_65[11],stage3_64[25],stage3_63[40]}
   );
   gpc117_4 gpc9142 (
      {stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18], stage2_63[19], stage2_63[20]},
      {stage2_64[62]},
      {stage2_65[2]},
      {stage3_66[12],stage3_65[12],stage3_64[26],stage3_63[41]}
   );
   gpc117_4 gpc9143 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[63]},
      {stage2_65[3]},
      {stage3_66[13],stage3_65[13],stage3_64[27],stage3_63[42]}
   );
   gpc117_4 gpc9144 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[64]},
      {stage2_65[4]},
      {stage3_66[14],stage3_65[14],stage3_64[28],stage3_63[43]}
   );
   gpc606_5 gpc9145 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40]},
      {stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9], stage2_65[10]},
      {stage3_67[0],stage3_66[15],stage3_65[15],stage3_64[29],stage3_63[44]}
   );
   gpc606_5 gpc9146 (
      {stage2_63[41], stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46]},
      {stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14], stage2_65[15], stage2_65[16]},
      {stage3_67[1],stage3_66[16],stage3_65[16],stage3_64[30],stage3_63[45]}
   );
   gpc606_5 gpc9147 (
      {stage2_63[47], stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52]},
      {stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20], stage2_65[21], stage2_65[22]},
      {stage3_67[2],stage3_66[17],stage3_65[17],stage3_64[31],stage3_63[46]}
   );
   gpc606_5 gpc9148 (
      {stage2_63[53], stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58]},
      {stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26], stage2_65[27], stage2_65[28]},
      {stage3_67[3],stage3_66[18],stage3_65[18],stage3_64[32],stage3_63[47]}
   );
   gpc606_5 gpc9149 (
      {stage2_63[59], stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64]},
      {stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32], stage2_65[33], stage2_65[34]},
      {stage3_67[4],stage3_66[19],stage3_65[19],stage3_64[33],stage3_63[48]}
   );
   gpc606_5 gpc9150 (
      {stage2_63[65], stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70]},
      {stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38], stage2_65[39], stage2_65[40]},
      {stage3_67[5],stage3_66[20],stage3_65[20],stage3_64[34],stage3_63[49]}
   );
   gpc606_5 gpc9151 (
      {stage2_63[71], stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76]},
      {stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44], stage2_65[45], stage2_65[46]},
      {stage3_67[6],stage3_66[21],stage3_65[21],stage3_64[35],stage3_63[50]}
   );
   gpc606_5 gpc9152 (
      {stage2_63[77], stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82]},
      {stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50], stage2_65[51], stage2_65[52]},
      {stage3_67[7],stage3_66[22],stage3_65[22],stage3_64[36],stage3_63[51]}
   );
   gpc606_5 gpc9153 (
      {stage2_63[83], stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88]},
      {stage2_65[53], stage2_65[54], stage2_65[55], stage2_65[56], stage2_65[57], stage2_65[58]},
      {stage3_67[8],stage3_66[23],stage3_65[23],stage3_64[37],stage3_63[52]}
   );
   gpc606_5 gpc9154 (
      {stage2_63[89], stage2_63[90], stage2_63[91], stage2_63[92], stage2_63[93], stage2_63[94]},
      {stage2_65[59], stage2_65[60], stage2_65[61], stage2_65[62], stage2_65[63], stage2_65[64]},
      {stage3_67[9],stage3_66[24],stage3_65[24],stage3_64[38],stage3_63[53]}
   );
   gpc606_5 gpc9155 (
      {stage2_64[65], stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[10],stage3_66[25],stage3_65[25],stage3_64[39]}
   );
   gpc606_5 gpc9156 (
      {stage2_64[71], stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[11],stage3_66[26],stage3_65[26],stage3_64[40]}
   );
   gpc606_5 gpc9157 (
      {stage2_64[77], stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[12],stage3_66[27],stage3_65[27],stage3_64[41]}
   );
   gpc606_5 gpc9158 (
      {stage2_64[83], stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[13],stage3_66[28],stage3_65[28],stage3_64[42]}
   );
   gpc606_5 gpc9159 (
      {stage2_64[89], stage2_64[90], stage2_64[91], stage2_64[92], stage2_64[93], stage2_64[94]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[14],stage3_66[29],stage3_65[29],stage3_64[43]}
   );
   gpc1_1 gpc9160 (
      {stage2_0[29]},
      {stage3_0[6]}
   );
   gpc1_1 gpc9161 (
      {stage2_0[30]},
      {stage3_0[7]}
   );
   gpc1_1 gpc9162 (
      {stage2_0[31]},
      {stage3_0[8]}
   );
   gpc1_1 gpc9163 (
      {stage2_0[32]},
      {stage3_0[9]}
   );
   gpc1_1 gpc9164 (
      {stage2_0[33]},
      {stage3_0[10]}
   );
   gpc1_1 gpc9165 (
      {stage2_1[22]},
      {stage3_1[9]}
   );
   gpc1_1 gpc9166 (
      {stage2_1[23]},
      {stage3_1[10]}
   );
   gpc1_1 gpc9167 (
      {stage2_1[24]},
      {stage3_1[11]}
   );
   gpc1_1 gpc9168 (
      {stage2_1[25]},
      {stage3_1[12]}
   );
   gpc1_1 gpc9169 (
      {stage2_1[26]},
      {stage3_1[13]}
   );
   gpc1_1 gpc9170 (
      {stage2_1[27]},
      {stage3_1[14]}
   );
   gpc1_1 gpc9171 (
      {stage2_1[28]},
      {stage3_1[15]}
   );
   gpc1_1 gpc9172 (
      {stage2_1[29]},
      {stage3_1[16]}
   );
   gpc1_1 gpc9173 (
      {stage2_1[30]},
      {stage3_1[17]}
   );
   gpc1_1 gpc9174 (
      {stage2_1[31]},
      {stage3_1[18]}
   );
   gpc1_1 gpc9175 (
      {stage2_1[32]},
      {stage3_1[19]}
   );
   gpc1_1 gpc9176 (
      {stage2_1[33]},
      {stage3_1[20]}
   );
   gpc1_1 gpc9177 (
      {stage2_1[34]},
      {stage3_1[21]}
   );
   gpc1_1 gpc9178 (
      {stage2_1[35]},
      {stage3_1[22]}
   );
   gpc1_1 gpc9179 (
      {stage2_1[36]},
      {stage3_1[23]}
   );
   gpc1_1 gpc9180 (
      {stage2_1[37]},
      {stage3_1[24]}
   );
   gpc1_1 gpc9181 (
      {stage2_1[38]},
      {stage3_1[25]}
   );
   gpc1_1 gpc9182 (
      {stage2_7[85]},
      {stage3_7[43]}
   );
   gpc1_1 gpc9183 (
      {stage2_7[86]},
      {stage3_7[44]}
   );
   gpc1_1 gpc9184 (
      {stage2_7[87]},
      {stage3_7[45]}
   );
   gpc1_1 gpc9185 (
      {stage2_7[88]},
      {stage3_7[46]}
   );
   gpc1_1 gpc9186 (
      {stage2_7[89]},
      {stage3_7[47]}
   );
   gpc1_1 gpc9187 (
      {stage2_7[90]},
      {stage3_7[48]}
   );
   gpc1_1 gpc9188 (
      {stage2_7[91]},
      {stage3_7[49]}
   );
   gpc1_1 gpc9189 (
      {stage2_7[92]},
      {stage3_7[50]}
   );
   gpc1_1 gpc9190 (
      {stage2_7[93]},
      {stage3_7[51]}
   );
   gpc1_1 gpc9191 (
      {stage2_7[94]},
      {stage3_7[52]}
   );
   gpc1_1 gpc9192 (
      {stage2_7[95]},
      {stage3_7[53]}
   );
   gpc1_1 gpc9193 (
      {stage2_7[96]},
      {stage3_7[54]}
   );
   gpc1_1 gpc9194 (
      {stage2_10[125]},
      {stage3_10[59]}
   );
   gpc1_1 gpc9195 (
      {stage2_10[126]},
      {stage3_10[60]}
   );
   gpc1_1 gpc9196 (
      {stage2_10[127]},
      {stage3_10[61]}
   );
   gpc1_1 gpc9197 (
      {stage2_10[128]},
      {stage3_10[62]}
   );
   gpc1_1 gpc9198 (
      {stage2_10[129]},
      {stage3_10[63]}
   );
   gpc1_1 gpc9199 (
      {stage2_10[130]},
      {stage3_10[64]}
   );
   gpc1_1 gpc9200 (
      {stage2_10[131]},
      {stage3_10[65]}
   );
   gpc1_1 gpc9201 (
      {stage2_10[132]},
      {stage3_10[66]}
   );
   gpc1_1 gpc9202 (
      {stage2_10[133]},
      {stage3_10[67]}
   );
   gpc1_1 gpc9203 (
      {stage2_11[125]},
      {stage3_11[50]}
   );
   gpc1_1 gpc9204 (
      {stage2_11[126]},
      {stage3_11[51]}
   );
   gpc1_1 gpc9205 (
      {stage2_11[127]},
      {stage3_11[52]}
   );
   gpc1_1 gpc9206 (
      {stage2_11[128]},
      {stage3_11[53]}
   );
   gpc1_1 gpc9207 (
      {stage2_11[129]},
      {stage3_11[54]}
   );
   gpc1_1 gpc9208 (
      {stage2_11[130]},
      {stage3_11[55]}
   );
   gpc1_1 gpc9209 (
      {stage2_11[131]},
      {stage3_11[56]}
   );
   gpc1_1 gpc9210 (
      {stage2_11[132]},
      {stage3_11[57]}
   );
   gpc1_1 gpc9211 (
      {stage2_11[133]},
      {stage3_11[58]}
   );
   gpc1_1 gpc9212 (
      {stage2_11[134]},
      {stage3_11[59]}
   );
   gpc1_1 gpc9213 (
      {stage2_11[135]},
      {stage3_11[60]}
   );
   gpc1_1 gpc9214 (
      {stage2_12[98]},
      {stage3_12[51]}
   );
   gpc1_1 gpc9215 (
      {stage2_12[99]},
      {stage3_12[52]}
   );
   gpc1_1 gpc9216 (
      {stage2_12[100]},
      {stage3_12[53]}
   );
   gpc1_1 gpc9217 (
      {stage2_12[101]},
      {stage3_12[54]}
   );
   gpc1_1 gpc9218 (
      {stage2_12[102]},
      {stage3_12[55]}
   );
   gpc1_1 gpc9219 (
      {stage2_12[103]},
      {stage3_12[56]}
   );
   gpc1_1 gpc9220 (
      {stage2_12[104]},
      {stage3_12[57]}
   );
   gpc1_1 gpc9221 (
      {stage2_12[105]},
      {stage3_12[58]}
   );
   gpc1_1 gpc9222 (
      {stage2_12[106]},
      {stage3_12[59]}
   );
   gpc1_1 gpc9223 (
      {stage2_12[107]},
      {stage3_12[60]}
   );
   gpc1_1 gpc9224 (
      {stage2_12[108]},
      {stage3_12[61]}
   );
   gpc1_1 gpc9225 (
      {stage2_12[109]},
      {stage3_12[62]}
   );
   gpc1_1 gpc9226 (
      {stage2_12[110]},
      {stage3_12[63]}
   );
   gpc1_1 gpc9227 (
      {stage2_12[111]},
      {stage3_12[64]}
   );
   gpc1_1 gpc9228 (
      {stage2_12[112]},
      {stage3_12[65]}
   );
   gpc1_1 gpc9229 (
      {stage2_12[113]},
      {stage3_12[66]}
   );
   gpc1_1 gpc9230 (
      {stage2_12[114]},
      {stage3_12[67]}
   );
   gpc1_1 gpc9231 (
      {stage2_12[115]},
      {stage3_12[68]}
   );
   gpc1_1 gpc9232 (
      {stage2_12[116]},
      {stage3_12[69]}
   );
   gpc1_1 gpc9233 (
      {stage2_12[117]},
      {stage3_12[70]}
   );
   gpc1_1 gpc9234 (
      {stage2_12[118]},
      {stage3_12[71]}
   );
   gpc1_1 gpc9235 (
      {stage2_12[119]},
      {stage3_12[72]}
   );
   gpc1_1 gpc9236 (
      {stage2_12[120]},
      {stage3_12[73]}
   );
   gpc1_1 gpc9237 (
      {stage2_12[121]},
      {stage3_12[74]}
   );
   gpc1_1 gpc9238 (
      {stage2_12[122]},
      {stage3_12[75]}
   );
   gpc1_1 gpc9239 (
      {stage2_12[123]},
      {stage3_12[76]}
   );
   gpc1_1 gpc9240 (
      {stage2_12[124]},
      {stage3_12[77]}
   );
   gpc1_1 gpc9241 (
      {stage2_12[125]},
      {stage3_12[78]}
   );
   gpc1_1 gpc9242 (
      {stage2_12[126]},
      {stage3_12[79]}
   );
   gpc1_1 gpc9243 (
      {stage2_12[127]},
      {stage3_12[80]}
   );
   gpc1_1 gpc9244 (
      {stage2_13[70]},
      {stage3_13[45]}
   );
   gpc1_1 gpc9245 (
      {stage2_13[71]},
      {stage3_13[46]}
   );
   gpc1_1 gpc9246 (
      {stage2_15[108]},
      {stage3_15[44]}
   );
   gpc1_1 gpc9247 (
      {stage2_15[109]},
      {stage3_15[45]}
   );
   gpc1_1 gpc9248 (
      {stage2_15[110]},
      {stage3_15[46]}
   );
   gpc1_1 gpc9249 (
      {stage2_15[111]},
      {stage3_15[47]}
   );
   gpc1_1 gpc9250 (
      {stage2_15[112]},
      {stage3_15[48]}
   );
   gpc1_1 gpc9251 (
      {stage2_15[113]},
      {stage3_15[49]}
   );
   gpc1_1 gpc9252 (
      {stage2_15[114]},
      {stage3_15[50]}
   );
   gpc1_1 gpc9253 (
      {stage2_16[96]},
      {stage3_16[45]}
   );
   gpc1_1 gpc9254 (
      {stage2_16[97]},
      {stage3_16[46]}
   );
   gpc1_1 gpc9255 (
      {stage2_16[98]},
      {stage3_16[47]}
   );
   gpc1_1 gpc9256 (
      {stage2_16[99]},
      {stage3_16[48]}
   );
   gpc1_1 gpc9257 (
      {stage2_16[100]},
      {stage3_16[49]}
   );
   gpc1_1 gpc9258 (
      {stage2_16[101]},
      {stage3_16[50]}
   );
   gpc1_1 gpc9259 (
      {stage2_16[102]},
      {stage3_16[51]}
   );
   gpc1_1 gpc9260 (
      {stage2_16[103]},
      {stage3_16[52]}
   );
   gpc1_1 gpc9261 (
      {stage2_16[104]},
      {stage3_16[53]}
   );
   gpc1_1 gpc9262 (
      {stage2_16[105]},
      {stage3_16[54]}
   );
   gpc1_1 gpc9263 (
      {stage2_16[106]},
      {stage3_16[55]}
   );
   gpc1_1 gpc9264 (
      {stage2_16[107]},
      {stage3_16[56]}
   );
   gpc1_1 gpc9265 (
      {stage2_16[108]},
      {stage3_16[57]}
   );
   gpc1_1 gpc9266 (
      {stage2_16[109]},
      {stage3_16[58]}
   );
   gpc1_1 gpc9267 (
      {stage2_17[80]},
      {stage3_17[34]}
   );
   gpc1_1 gpc9268 (
      {stage2_17[81]},
      {stage3_17[35]}
   );
   gpc1_1 gpc9269 (
      {stage2_17[82]},
      {stage3_17[36]}
   );
   gpc1_1 gpc9270 (
      {stage2_17[83]},
      {stage3_17[37]}
   );
   gpc1_1 gpc9271 (
      {stage2_17[84]},
      {stage3_17[38]}
   );
   gpc1_1 gpc9272 (
      {stage2_17[85]},
      {stage3_17[39]}
   );
   gpc1_1 gpc9273 (
      {stage2_17[86]},
      {stage3_17[40]}
   );
   gpc1_1 gpc9274 (
      {stage2_17[87]},
      {stage3_17[41]}
   );
   gpc1_1 gpc9275 (
      {stage2_17[88]},
      {stage3_17[42]}
   );
   gpc1_1 gpc9276 (
      {stage2_17[89]},
      {stage3_17[43]}
   );
   gpc1_1 gpc9277 (
      {stage2_18[147]},
      {stage3_18[49]}
   );
   gpc1_1 gpc9278 (
      {stage2_18[148]},
      {stage3_18[50]}
   );
   gpc1_1 gpc9279 (
      {stage2_18[149]},
      {stage3_18[51]}
   );
   gpc1_1 gpc9280 (
      {stage2_18[150]},
      {stage3_18[52]}
   );
   gpc1_1 gpc9281 (
      {stage2_18[151]},
      {stage3_18[53]}
   );
   gpc1_1 gpc9282 (
      {stage2_18[152]},
      {stage3_18[54]}
   );
   gpc1_1 gpc9283 (
      {stage2_18[153]},
      {stage3_18[55]}
   );
   gpc1_1 gpc9284 (
      {stage2_18[154]},
      {stage3_18[56]}
   );
   gpc1_1 gpc9285 (
      {stage2_18[155]},
      {stage3_18[57]}
   );
   gpc1_1 gpc9286 (
      {stage2_18[156]},
      {stage3_18[58]}
   );
   gpc1_1 gpc9287 (
      {stage2_18[157]},
      {stage3_18[59]}
   );
   gpc1_1 gpc9288 (
      {stage2_18[158]},
      {stage3_18[60]}
   );
   gpc1_1 gpc9289 (
      {stage2_18[159]},
      {stage3_18[61]}
   );
   gpc1_1 gpc9290 (
      {stage2_18[160]},
      {stage3_18[62]}
   );
   gpc1_1 gpc9291 (
      {stage2_18[161]},
      {stage3_18[63]}
   );
   gpc1_1 gpc9292 (
      {stage2_20[72]},
      {stage3_20[42]}
   );
   gpc1_1 gpc9293 (
      {stage2_20[73]},
      {stage3_20[43]}
   );
   gpc1_1 gpc9294 (
      {stage2_20[74]},
      {stage3_20[44]}
   );
   gpc1_1 gpc9295 (
      {stage2_20[75]},
      {stage3_20[45]}
   );
   gpc1_1 gpc9296 (
      {stage2_20[76]},
      {stage3_20[46]}
   );
   gpc1_1 gpc9297 (
      {stage2_20[77]},
      {stage3_20[47]}
   );
   gpc1_1 gpc9298 (
      {stage2_20[78]},
      {stage3_20[48]}
   );
   gpc1_1 gpc9299 (
      {stage2_20[79]},
      {stage3_20[49]}
   );
   gpc1_1 gpc9300 (
      {stage2_20[80]},
      {stage3_20[50]}
   );
   gpc1_1 gpc9301 (
      {stage2_20[81]},
      {stage3_20[51]}
   );
   gpc1_1 gpc9302 (
      {stage2_20[82]},
      {stage3_20[52]}
   );
   gpc1_1 gpc9303 (
      {stage2_20[83]},
      {stage3_20[53]}
   );
   gpc1_1 gpc9304 (
      {stage2_20[84]},
      {stage3_20[54]}
   );
   gpc1_1 gpc9305 (
      {stage2_20[85]},
      {stage3_20[55]}
   );
   gpc1_1 gpc9306 (
      {stage2_20[86]},
      {stage3_20[56]}
   );
   gpc1_1 gpc9307 (
      {stage2_20[87]},
      {stage3_20[57]}
   );
   gpc1_1 gpc9308 (
      {stage2_21[86]},
      {stage3_21[37]}
   );
   gpc1_1 gpc9309 (
      {stage2_21[87]},
      {stage3_21[38]}
   );
   gpc1_1 gpc9310 (
      {stage2_21[88]},
      {stage3_21[39]}
   );
   gpc1_1 gpc9311 (
      {stage2_21[89]},
      {stage3_21[40]}
   );
   gpc1_1 gpc9312 (
      {stage2_21[90]},
      {stage3_21[41]}
   );
   gpc1_1 gpc9313 (
      {stage2_21[91]},
      {stage3_21[42]}
   );
   gpc1_1 gpc9314 (
      {stage2_21[92]},
      {stage3_21[43]}
   );
   gpc1_1 gpc9315 (
      {stage2_21[93]},
      {stage3_21[44]}
   );
   gpc1_1 gpc9316 (
      {stage2_21[94]},
      {stage3_21[45]}
   );
   gpc1_1 gpc9317 (
      {stage2_21[95]},
      {stage3_21[46]}
   );
   gpc1_1 gpc9318 (
      {stage2_21[96]},
      {stage3_21[47]}
   );
   gpc1_1 gpc9319 (
      {stage2_21[97]},
      {stage3_21[48]}
   );
   gpc1_1 gpc9320 (
      {stage2_21[98]},
      {stage3_21[49]}
   );
   gpc1_1 gpc9321 (
      {stage2_21[99]},
      {stage3_21[50]}
   );
   gpc1_1 gpc9322 (
      {stage2_21[100]},
      {stage3_21[51]}
   );
   gpc1_1 gpc9323 (
      {stage2_21[101]},
      {stage3_21[52]}
   );
   gpc1_1 gpc9324 (
      {stage2_21[102]},
      {stage3_21[53]}
   );
   gpc1_1 gpc9325 (
      {stage2_21[103]},
      {stage3_21[54]}
   );
   gpc1_1 gpc9326 (
      {stage2_21[104]},
      {stage3_21[55]}
   );
   gpc1_1 gpc9327 (
      {stage2_21[105]},
      {stage3_21[56]}
   );
   gpc1_1 gpc9328 (
      {stage2_21[106]},
      {stage3_21[57]}
   );
   gpc1_1 gpc9329 (
      {stage2_21[107]},
      {stage3_21[58]}
   );
   gpc1_1 gpc9330 (
      {stage2_21[108]},
      {stage3_21[59]}
   );
   gpc1_1 gpc9331 (
      {stage2_21[109]},
      {stage3_21[60]}
   );
   gpc1_1 gpc9332 (
      {stage2_21[110]},
      {stage3_21[61]}
   );
   gpc1_1 gpc9333 (
      {stage2_21[111]},
      {stage3_21[62]}
   );
   gpc1_1 gpc9334 (
      {stage2_22[108]},
      {stage3_22[48]}
   );
   gpc1_1 gpc9335 (
      {stage2_22[109]},
      {stage3_22[49]}
   );
   gpc1_1 gpc9336 (
      {stage2_23[89]},
      {stage3_23[40]}
   );
   gpc1_1 gpc9337 (
      {stage2_23[90]},
      {stage3_23[41]}
   );
   gpc1_1 gpc9338 (
      {stage2_23[91]},
      {stage3_23[42]}
   );
   gpc1_1 gpc9339 (
      {stage2_23[92]},
      {stage3_23[43]}
   );
   gpc1_1 gpc9340 (
      {stage2_23[93]},
      {stage3_23[44]}
   );
   gpc1_1 gpc9341 (
      {stage2_23[94]},
      {stage3_23[45]}
   );
   gpc1_1 gpc9342 (
      {stage2_23[95]},
      {stage3_23[46]}
   );
   gpc1_1 gpc9343 (
      {stage2_23[96]},
      {stage3_23[47]}
   );
   gpc1_1 gpc9344 (
      {stage2_23[97]},
      {stage3_23[48]}
   );
   gpc1_1 gpc9345 (
      {stage2_25[102]},
      {stage3_25[31]}
   );
   gpc1_1 gpc9346 (
      {stage2_25[103]},
      {stage3_25[32]}
   );
   gpc1_1 gpc9347 (
      {stage2_25[104]},
      {stage3_25[33]}
   );
   gpc1_1 gpc9348 (
      {stage2_25[105]},
      {stage3_25[34]}
   );
   gpc1_1 gpc9349 (
      {stage2_25[106]},
      {stage3_25[35]}
   );
   gpc1_1 gpc9350 (
      {stage2_25[107]},
      {stage3_25[36]}
   );
   gpc1_1 gpc9351 (
      {stage2_25[108]},
      {stage3_25[37]}
   );
   gpc1_1 gpc9352 (
      {stage2_25[109]},
      {stage3_25[38]}
   );
   gpc1_1 gpc9353 (
      {stage2_25[110]},
      {stage3_25[39]}
   );
   gpc1_1 gpc9354 (
      {stage2_25[111]},
      {stage3_25[40]}
   );
   gpc1_1 gpc9355 (
      {stage2_25[112]},
      {stage3_25[41]}
   );
   gpc1_1 gpc9356 (
      {stage2_25[113]},
      {stage3_25[42]}
   );
   gpc1_1 gpc9357 (
      {stage2_25[114]},
      {stage3_25[43]}
   );
   gpc1_1 gpc9358 (
      {stage2_25[115]},
      {stage3_25[44]}
   );
   gpc1_1 gpc9359 (
      {stage2_25[116]},
      {stage3_25[45]}
   );
   gpc1_1 gpc9360 (
      {stage2_25[117]},
      {stage3_25[46]}
   );
   gpc1_1 gpc9361 (
      {stage2_25[118]},
      {stage3_25[47]}
   );
   gpc1_1 gpc9362 (
      {stage2_25[119]},
      {stage3_25[48]}
   );
   gpc1_1 gpc9363 (
      {stage2_25[120]},
      {stage3_25[49]}
   );
   gpc1_1 gpc9364 (
      {stage2_25[121]},
      {stage3_25[50]}
   );
   gpc1_1 gpc9365 (
      {stage2_25[122]},
      {stage3_25[51]}
   );
   gpc1_1 gpc9366 (
      {stage2_26[126]},
      {stage3_26[47]}
   );
   gpc1_1 gpc9367 (
      {stage2_26[127]},
      {stage3_26[48]}
   );
   gpc1_1 gpc9368 (
      {stage2_26[128]},
      {stage3_26[49]}
   );
   gpc1_1 gpc9369 (
      {stage2_26[129]},
      {stage3_26[50]}
   );
   gpc1_1 gpc9370 (
      {stage2_26[130]},
      {stage3_26[51]}
   );
   gpc1_1 gpc9371 (
      {stage2_28[44]},
      {stage3_28[34]}
   );
   gpc1_1 gpc9372 (
      {stage2_28[45]},
      {stage3_28[35]}
   );
   gpc1_1 gpc9373 (
      {stage2_28[46]},
      {stage3_28[36]}
   );
   gpc1_1 gpc9374 (
      {stage2_28[47]},
      {stage3_28[37]}
   );
   gpc1_1 gpc9375 (
      {stage2_28[48]},
      {stage3_28[38]}
   );
   gpc1_1 gpc9376 (
      {stage2_28[49]},
      {stage3_28[39]}
   );
   gpc1_1 gpc9377 (
      {stage2_28[50]},
      {stage3_28[40]}
   );
   gpc1_1 gpc9378 (
      {stage2_28[51]},
      {stage3_28[41]}
   );
   gpc1_1 gpc9379 (
      {stage2_28[52]},
      {stage3_28[42]}
   );
   gpc1_1 gpc9380 (
      {stage2_28[53]},
      {stage3_28[43]}
   );
   gpc1_1 gpc9381 (
      {stage2_28[54]},
      {stage3_28[44]}
   );
   gpc1_1 gpc9382 (
      {stage2_28[55]},
      {stage3_28[45]}
   );
   gpc1_1 gpc9383 (
      {stage2_28[56]},
      {stage3_28[46]}
   );
   gpc1_1 gpc9384 (
      {stage2_28[57]},
      {stage3_28[47]}
   );
   gpc1_1 gpc9385 (
      {stage2_28[58]},
      {stage3_28[48]}
   );
   gpc1_1 gpc9386 (
      {stage2_28[59]},
      {stage3_28[49]}
   );
   gpc1_1 gpc9387 (
      {stage2_28[60]},
      {stage3_28[50]}
   );
   gpc1_1 gpc9388 (
      {stage2_28[61]},
      {stage3_28[51]}
   );
   gpc1_1 gpc9389 (
      {stage2_28[62]},
      {stage3_28[52]}
   );
   gpc1_1 gpc9390 (
      {stage2_28[63]},
      {stage3_28[53]}
   );
   gpc1_1 gpc9391 (
      {stage2_28[64]},
      {stage3_28[54]}
   );
   gpc1_1 gpc9392 (
      {stage2_28[65]},
      {stage3_28[55]}
   );
   gpc1_1 gpc9393 (
      {stage2_28[66]},
      {stage3_28[56]}
   );
   gpc1_1 gpc9394 (
      {stage2_28[67]},
      {stage3_28[57]}
   );
   gpc1_1 gpc9395 (
      {stage2_28[68]},
      {stage3_28[58]}
   );
   gpc1_1 gpc9396 (
      {stage2_28[69]},
      {stage3_28[59]}
   );
   gpc1_1 gpc9397 (
      {stage2_28[70]},
      {stage3_28[60]}
   );
   gpc1_1 gpc9398 (
      {stage2_28[71]},
      {stage3_28[61]}
   );
   gpc1_1 gpc9399 (
      {stage2_28[72]},
      {stage3_28[62]}
   );
   gpc1_1 gpc9400 (
      {stage2_28[73]},
      {stage3_28[63]}
   );
   gpc1_1 gpc9401 (
      {stage2_28[74]},
      {stage3_28[64]}
   );
   gpc1_1 gpc9402 (
      {stage2_28[75]},
      {stage3_28[65]}
   );
   gpc1_1 gpc9403 (
      {stage2_28[76]},
      {stage3_28[66]}
   );
   gpc1_1 gpc9404 (
      {stage2_28[77]},
      {stage3_28[67]}
   );
   gpc1_1 gpc9405 (
      {stage2_28[78]},
      {stage3_28[68]}
   );
   gpc1_1 gpc9406 (
      {stage2_28[79]},
      {stage3_28[69]}
   );
   gpc1_1 gpc9407 (
      {stage2_29[102]},
      {stage3_29[49]}
   );
   gpc1_1 gpc9408 (
      {stage2_29[103]},
      {stage3_29[50]}
   );
   gpc1_1 gpc9409 (
      {stage2_29[104]},
      {stage3_29[51]}
   );
   gpc1_1 gpc9410 (
      {stage2_29[105]},
      {stage3_29[52]}
   );
   gpc1_1 gpc9411 (
      {stage2_29[106]},
      {stage3_29[53]}
   );
   gpc1_1 gpc9412 (
      {stage2_29[107]},
      {stage3_29[54]}
   );
   gpc1_1 gpc9413 (
      {stage2_29[108]},
      {stage3_29[55]}
   );
   gpc1_1 gpc9414 (
      {stage2_29[109]},
      {stage3_29[56]}
   );
   gpc1_1 gpc9415 (
      {stage2_29[110]},
      {stage3_29[57]}
   );
   gpc1_1 gpc9416 (
      {stage2_29[111]},
      {stage3_29[58]}
   );
   gpc1_1 gpc9417 (
      {stage2_30[93]},
      {stage3_30[32]}
   );
   gpc1_1 gpc9418 (
      {stage2_30[94]},
      {stage3_30[33]}
   );
   gpc1_1 gpc9419 (
      {stage2_30[95]},
      {stage3_30[34]}
   );
   gpc1_1 gpc9420 (
      {stage2_30[96]},
      {stage3_30[35]}
   );
   gpc1_1 gpc9421 (
      {stage2_30[97]},
      {stage3_30[36]}
   );
   gpc1_1 gpc9422 (
      {stage2_30[98]},
      {stage3_30[37]}
   );
   gpc1_1 gpc9423 (
      {stage2_30[99]},
      {stage3_30[38]}
   );
   gpc1_1 gpc9424 (
      {stage2_31[124]},
      {stage3_31[38]}
   );
   gpc1_1 gpc9425 (
      {stage2_31[125]},
      {stage3_31[39]}
   );
   gpc1_1 gpc9426 (
      {stage2_31[126]},
      {stage3_31[40]}
   );
   gpc1_1 gpc9427 (
      {stage2_31[127]},
      {stage3_31[41]}
   );
   gpc1_1 gpc9428 (
      {stage2_32[112]},
      {stage3_32[50]}
   );
   gpc1_1 gpc9429 (
      {stage2_32[113]},
      {stage3_32[51]}
   );
   gpc1_1 gpc9430 (
      {stage2_32[114]},
      {stage3_32[52]}
   );
   gpc1_1 gpc9431 (
      {stage2_32[115]},
      {stage3_32[53]}
   );
   gpc1_1 gpc9432 (
      {stage2_32[116]},
      {stage3_32[54]}
   );
   gpc1_1 gpc9433 (
      {stage2_32[117]},
      {stage3_32[55]}
   );
   gpc1_1 gpc9434 (
      {stage2_33[91]},
      {stage3_33[45]}
   );
   gpc1_1 gpc9435 (
      {stage2_33[92]},
      {stage3_33[46]}
   );
   gpc1_1 gpc9436 (
      {stage2_33[93]},
      {stage3_33[47]}
   );
   gpc1_1 gpc9437 (
      {stage2_33[94]},
      {stage3_33[48]}
   );
   gpc1_1 gpc9438 (
      {stage2_33[95]},
      {stage3_33[49]}
   );
   gpc1_1 gpc9439 (
      {stage2_33[96]},
      {stage3_33[50]}
   );
   gpc1_1 gpc9440 (
      {stage2_33[97]},
      {stage3_33[51]}
   );
   gpc1_1 gpc9441 (
      {stage2_33[98]},
      {stage3_33[52]}
   );
   gpc1_1 gpc9442 (
      {stage2_33[99]},
      {stage3_33[53]}
   );
   gpc1_1 gpc9443 (
      {stage2_33[100]},
      {stage3_33[54]}
   );
   gpc1_1 gpc9444 (
      {stage2_33[101]},
      {stage3_33[55]}
   );
   gpc1_1 gpc9445 (
      {stage2_33[102]},
      {stage3_33[56]}
   );
   gpc1_1 gpc9446 (
      {stage2_33[103]},
      {stage3_33[57]}
   );
   gpc1_1 gpc9447 (
      {stage2_33[104]},
      {stage3_33[58]}
   );
   gpc1_1 gpc9448 (
      {stage2_33[105]},
      {stage3_33[59]}
   );
   gpc1_1 gpc9449 (
      {stage2_33[106]},
      {stage3_33[60]}
   );
   gpc1_1 gpc9450 (
      {stage2_33[107]},
      {stage3_33[61]}
   );
   gpc1_1 gpc9451 (
      {stage2_33[108]},
      {stage3_33[62]}
   );
   gpc1_1 gpc9452 (
      {stage2_36[114]},
      {stage3_36[50]}
   );
   gpc1_1 gpc9453 (
      {stage2_36[115]},
      {stage3_36[51]}
   );
   gpc1_1 gpc9454 (
      {stage2_36[116]},
      {stage3_36[52]}
   );
   gpc1_1 gpc9455 (
      {stage2_36[117]},
      {stage3_36[53]}
   );
   gpc1_1 gpc9456 (
      {stage2_36[118]},
      {stage3_36[54]}
   );
   gpc1_1 gpc9457 (
      {stage2_36[119]},
      {stage3_36[55]}
   );
   gpc1_1 gpc9458 (
      {stage2_38[81]},
      {stage3_38[50]}
   );
   gpc1_1 gpc9459 (
      {stage2_38[82]},
      {stage3_38[51]}
   );
   gpc1_1 gpc9460 (
      {stage2_38[83]},
      {stage3_38[52]}
   );
   gpc1_1 gpc9461 (
      {stage2_38[84]},
      {stage3_38[53]}
   );
   gpc1_1 gpc9462 (
      {stage2_38[85]},
      {stage3_38[54]}
   );
   gpc1_1 gpc9463 (
      {stage2_38[86]},
      {stage3_38[55]}
   );
   gpc1_1 gpc9464 (
      {stage2_38[87]},
      {stage3_38[56]}
   );
   gpc1_1 gpc9465 (
      {stage2_38[88]},
      {stage3_38[57]}
   );
   gpc1_1 gpc9466 (
      {stage2_38[89]},
      {stage3_38[58]}
   );
   gpc1_1 gpc9467 (
      {stage2_38[90]},
      {stage3_38[59]}
   );
   gpc1_1 gpc9468 (
      {stage2_38[91]},
      {stage3_38[60]}
   );
   gpc1_1 gpc9469 (
      {stage2_38[92]},
      {stage3_38[61]}
   );
   gpc1_1 gpc9470 (
      {stage2_38[93]},
      {stage3_38[62]}
   );
   gpc1_1 gpc9471 (
      {stage2_38[94]},
      {stage3_38[63]}
   );
   gpc1_1 gpc9472 (
      {stage2_38[95]},
      {stage3_38[64]}
   );
   gpc1_1 gpc9473 (
      {stage2_38[96]},
      {stage3_38[65]}
   );
   gpc1_1 gpc9474 (
      {stage2_38[97]},
      {stage3_38[66]}
   );
   gpc1_1 gpc9475 (
      {stage2_38[98]},
      {stage3_38[67]}
   );
   gpc1_1 gpc9476 (
      {stage2_38[99]},
      {stage3_38[68]}
   );
   gpc1_1 gpc9477 (
      {stage2_39[100]},
      {stage3_39[52]}
   );
   gpc1_1 gpc9478 (
      {stage2_39[101]},
      {stage3_39[53]}
   );
   gpc1_1 gpc9479 (
      {stage2_39[102]},
      {stage3_39[54]}
   );
   gpc1_1 gpc9480 (
      {stage2_39[103]},
      {stage3_39[55]}
   );
   gpc1_1 gpc9481 (
      {stage2_39[104]},
      {stage3_39[56]}
   );
   gpc1_1 gpc9482 (
      {stage2_39[105]},
      {stage3_39[57]}
   );
   gpc1_1 gpc9483 (
      {stage2_39[106]},
      {stage3_39[58]}
   );
   gpc1_1 gpc9484 (
      {stage2_39[107]},
      {stage3_39[59]}
   );
   gpc1_1 gpc9485 (
      {stage2_40[131]},
      {stage3_40[37]}
   );
   gpc1_1 gpc9486 (
      {stage2_40[132]},
      {stage3_40[38]}
   );
   gpc1_1 gpc9487 (
      {stage2_40[133]},
      {stage3_40[39]}
   );
   gpc1_1 gpc9488 (
      {stage2_40[134]},
      {stage3_40[40]}
   );
   gpc1_1 gpc9489 (
      {stage2_40[135]},
      {stage3_40[41]}
   );
   gpc1_1 gpc9490 (
      {stage2_40[136]},
      {stage3_40[42]}
   );
   gpc1_1 gpc9491 (
      {stage2_40[137]},
      {stage3_40[43]}
   );
   gpc1_1 gpc9492 (
      {stage2_40[138]},
      {stage3_40[44]}
   );
   gpc1_1 gpc9493 (
      {stage2_40[139]},
      {stage3_40[45]}
   );
   gpc1_1 gpc9494 (
      {stage2_41[102]},
      {stage3_41[36]}
   );
   gpc1_1 gpc9495 (
      {stage2_41[103]},
      {stage3_41[37]}
   );
   gpc1_1 gpc9496 (
      {stage2_41[104]},
      {stage3_41[38]}
   );
   gpc1_1 gpc9497 (
      {stage2_41[105]},
      {stage3_41[39]}
   );
   gpc1_1 gpc9498 (
      {stage2_41[106]},
      {stage3_41[40]}
   );
   gpc1_1 gpc9499 (
      {stage2_41[107]},
      {stage3_41[41]}
   );
   gpc1_1 gpc9500 (
      {stage2_41[108]},
      {stage3_41[42]}
   );
   gpc1_1 gpc9501 (
      {stage2_41[109]},
      {stage3_41[43]}
   );
   gpc1_1 gpc9502 (
      {stage2_41[110]},
      {stage3_41[44]}
   );
   gpc1_1 gpc9503 (
      {stage2_41[111]},
      {stage3_41[45]}
   );
   gpc1_1 gpc9504 (
      {stage2_41[112]},
      {stage3_41[46]}
   );
   gpc1_1 gpc9505 (
      {stage2_41[113]},
      {stage3_41[47]}
   );
   gpc1_1 gpc9506 (
      {stage2_41[114]},
      {stage3_41[48]}
   );
   gpc1_1 gpc9507 (
      {stage2_41[115]},
      {stage3_41[49]}
   );
   gpc1_1 gpc9508 (
      {stage2_41[116]},
      {stage3_41[50]}
   );
   gpc1_1 gpc9509 (
      {stage2_41[117]},
      {stage3_41[51]}
   );
   gpc1_1 gpc9510 (
      {stage2_41[118]},
      {stage3_41[52]}
   );
   gpc1_1 gpc9511 (
      {stage2_41[119]},
      {stage3_41[53]}
   );
   gpc1_1 gpc9512 (
      {stage2_41[120]},
      {stage3_41[54]}
   );
   gpc1_1 gpc9513 (
      {stage2_41[121]},
      {stage3_41[55]}
   );
   gpc1_1 gpc9514 (
      {stage2_41[122]},
      {stage3_41[56]}
   );
   gpc1_1 gpc9515 (
      {stage2_42[74]},
      {stage3_42[46]}
   );
   gpc1_1 gpc9516 (
      {stage2_42[75]},
      {stage3_42[47]}
   );
   gpc1_1 gpc9517 (
      {stage2_42[76]},
      {stage3_42[48]}
   );
   gpc1_1 gpc9518 (
      {stage2_42[77]},
      {stage3_42[49]}
   );
   gpc1_1 gpc9519 (
      {stage2_42[78]},
      {stage3_42[50]}
   );
   gpc1_1 gpc9520 (
      {stage2_42[79]},
      {stage3_42[51]}
   );
   gpc1_1 gpc9521 (
      {stage2_42[80]},
      {stage3_42[52]}
   );
   gpc1_1 gpc9522 (
      {stage2_42[81]},
      {stage3_42[53]}
   );
   gpc1_1 gpc9523 (
      {stage2_43[98]},
      {stage3_43[47]}
   );
   gpc1_1 gpc9524 (
      {stage2_43[99]},
      {stage3_43[48]}
   );
   gpc1_1 gpc9525 (
      {stage2_43[100]},
      {stage3_43[49]}
   );
   gpc1_1 gpc9526 (
      {stage2_43[101]},
      {stage3_43[50]}
   );
   gpc1_1 gpc9527 (
      {stage2_43[102]},
      {stage3_43[51]}
   );
   gpc1_1 gpc9528 (
      {stage2_43[103]},
      {stage3_43[52]}
   );
   gpc1_1 gpc9529 (
      {stage2_43[104]},
      {stage3_43[53]}
   );
   gpc1_1 gpc9530 (
      {stage2_43[105]},
      {stage3_43[54]}
   );
   gpc1_1 gpc9531 (
      {stage2_43[106]},
      {stage3_43[55]}
   );
   gpc1_1 gpc9532 (
      {stage2_43[107]},
      {stage3_43[56]}
   );
   gpc1_1 gpc9533 (
      {stage2_43[108]},
      {stage3_43[57]}
   );
   gpc1_1 gpc9534 (
      {stage2_43[109]},
      {stage3_43[58]}
   );
   gpc1_1 gpc9535 (
      {stage2_43[110]},
      {stage3_43[59]}
   );
   gpc1_1 gpc9536 (
      {stage2_44[86]},
      {stage3_44[33]}
   );
   gpc1_1 gpc9537 (
      {stage2_44[87]},
      {stage3_44[34]}
   );
   gpc1_1 gpc9538 (
      {stage2_44[88]},
      {stage3_44[35]}
   );
   gpc1_1 gpc9539 (
      {stage2_44[89]},
      {stage3_44[36]}
   );
   gpc1_1 gpc9540 (
      {stage2_44[90]},
      {stage3_44[37]}
   );
   gpc1_1 gpc9541 (
      {stage2_44[91]},
      {stage3_44[38]}
   );
   gpc1_1 gpc9542 (
      {stage2_44[92]},
      {stage3_44[39]}
   );
   gpc1_1 gpc9543 (
      {stage2_44[93]},
      {stage3_44[40]}
   );
   gpc1_1 gpc9544 (
      {stage2_44[94]},
      {stage3_44[41]}
   );
   gpc1_1 gpc9545 (
      {stage2_44[95]},
      {stage3_44[42]}
   );
   gpc1_1 gpc9546 (
      {stage2_44[96]},
      {stage3_44[43]}
   );
   gpc1_1 gpc9547 (
      {stage2_44[97]},
      {stage3_44[44]}
   );
   gpc1_1 gpc9548 (
      {stage2_44[98]},
      {stage3_44[45]}
   );
   gpc1_1 gpc9549 (
      {stage2_44[99]},
      {stage3_44[46]}
   );
   gpc1_1 gpc9550 (
      {stage2_44[100]},
      {stage3_44[47]}
   );
   gpc1_1 gpc9551 (
      {stage2_44[101]},
      {stage3_44[48]}
   );
   gpc1_1 gpc9552 (
      {stage2_44[102]},
      {stage3_44[49]}
   );
   gpc1_1 gpc9553 (
      {stage2_44[103]},
      {stage3_44[50]}
   );
   gpc1_1 gpc9554 (
      {stage2_44[104]},
      {stage3_44[51]}
   );
   gpc1_1 gpc9555 (
      {stage2_44[105]},
      {stage3_44[52]}
   );
   gpc1_1 gpc9556 (
      {stage2_44[106]},
      {stage3_44[53]}
   );
   gpc1_1 gpc9557 (
      {stage2_44[107]},
      {stage3_44[54]}
   );
   gpc1_1 gpc9558 (
      {stage2_44[108]},
      {stage3_44[55]}
   );
   gpc1_1 gpc9559 (
      {stage2_44[109]},
      {stage3_44[56]}
   );
   gpc1_1 gpc9560 (
      {stage2_44[110]},
      {stage3_44[57]}
   );
   gpc1_1 gpc9561 (
      {stage2_44[111]},
      {stage3_44[58]}
   );
   gpc1_1 gpc9562 (
      {stage2_44[112]},
      {stage3_44[59]}
   );
   gpc1_1 gpc9563 (
      {stage2_44[113]},
      {stage3_44[60]}
   );
   gpc1_1 gpc9564 (
      {stage2_44[114]},
      {stage3_44[61]}
   );
   gpc1_1 gpc9565 (
      {stage2_44[115]},
      {stage3_44[62]}
   );
   gpc1_1 gpc9566 (
      {stage2_44[116]},
      {stage3_44[63]}
   );
   gpc1_1 gpc9567 (
      {stage2_44[117]},
      {stage3_44[64]}
   );
   gpc1_1 gpc9568 (
      {stage2_44[118]},
      {stage3_44[65]}
   );
   gpc1_1 gpc9569 (
      {stage2_44[119]},
      {stage3_44[66]}
   );
   gpc1_1 gpc9570 (
      {stage2_44[120]},
      {stage3_44[67]}
   );
   gpc1_1 gpc9571 (
      {stage2_44[121]},
      {stage3_44[68]}
   );
   gpc1_1 gpc9572 (
      {stage2_44[122]},
      {stage3_44[69]}
   );
   gpc1_1 gpc9573 (
      {stage2_44[123]},
      {stage3_44[70]}
   );
   gpc1_1 gpc9574 (
      {stage2_44[124]},
      {stage3_44[71]}
   );
   gpc1_1 gpc9575 (
      {stage2_44[125]},
      {stage3_44[72]}
   );
   gpc1_1 gpc9576 (
      {stage2_44[126]},
      {stage3_44[73]}
   );
   gpc1_1 gpc9577 (
      {stage2_44[127]},
      {stage3_44[74]}
   );
   gpc1_1 gpc9578 (
      {stage2_44[128]},
      {stage3_44[75]}
   );
   gpc1_1 gpc9579 (
      {stage2_44[129]},
      {stage3_44[76]}
   );
   gpc1_1 gpc9580 (
      {stage2_44[130]},
      {stage3_44[77]}
   );
   gpc1_1 gpc9581 (
      {stage2_44[131]},
      {stage3_44[78]}
   );
   gpc1_1 gpc9582 (
      {stage2_44[132]},
      {stage3_44[79]}
   );
   gpc1_1 gpc9583 (
      {stage2_44[133]},
      {stage3_44[80]}
   );
   gpc1_1 gpc9584 (
      {stage2_44[134]},
      {stage3_44[81]}
   );
   gpc1_1 gpc9585 (
      {stage2_44[135]},
      {stage3_44[82]}
   );
   gpc1_1 gpc9586 (
      {stage2_44[136]},
      {stage3_44[83]}
   );
   gpc1_1 gpc9587 (
      {stage2_44[137]},
      {stage3_44[84]}
   );
   gpc1_1 gpc9588 (
      {stage2_45[126]},
      {stage3_45[34]}
   );
   gpc1_1 gpc9589 (
      {stage2_45[127]},
      {stage3_45[35]}
   );
   gpc1_1 gpc9590 (
      {stage2_45[128]},
      {stage3_45[36]}
   );
   gpc1_1 gpc9591 (
      {stage2_45[129]},
      {stage3_45[37]}
   );
   gpc1_1 gpc9592 (
      {stage2_45[130]},
      {stage3_45[38]}
   );
   gpc1_1 gpc9593 (
      {stage2_45[131]},
      {stage3_45[39]}
   );
   gpc1_1 gpc9594 (
      {stage2_47[83]},
      {stage3_47[49]}
   );
   gpc1_1 gpc9595 (
      {stage2_47[84]},
      {stage3_47[50]}
   );
   gpc1_1 gpc9596 (
      {stage2_47[85]},
      {stage3_47[51]}
   );
   gpc1_1 gpc9597 (
      {stage2_47[86]},
      {stage3_47[52]}
   );
   gpc1_1 gpc9598 (
      {stage2_47[87]},
      {stage3_47[53]}
   );
   gpc1_1 gpc9599 (
      {stage2_47[88]},
      {stage3_47[54]}
   );
   gpc1_1 gpc9600 (
      {stage2_47[89]},
      {stage3_47[55]}
   );
   gpc1_1 gpc9601 (
      {stage2_47[90]},
      {stage3_47[56]}
   );
   gpc1_1 gpc9602 (
      {stage2_47[91]},
      {stage3_47[57]}
   );
   gpc1_1 gpc9603 (
      {stage2_47[92]},
      {stage3_47[58]}
   );
   gpc1_1 gpc9604 (
      {stage2_47[93]},
      {stage3_47[59]}
   );
   gpc1_1 gpc9605 (
      {stage2_47[94]},
      {stage3_47[60]}
   );
   gpc1_1 gpc9606 (
      {stage2_47[95]},
      {stage3_47[61]}
   );
   gpc1_1 gpc9607 (
      {stage2_47[96]},
      {stage3_47[62]}
   );
   gpc1_1 gpc9608 (
      {stage2_47[97]},
      {stage3_47[63]}
   );
   gpc1_1 gpc9609 (
      {stage2_47[98]},
      {stage3_47[64]}
   );
   gpc1_1 gpc9610 (
      {stage2_47[99]},
      {stage3_47[65]}
   );
   gpc1_1 gpc9611 (
      {stage2_47[100]},
      {stage3_47[66]}
   );
   gpc1_1 gpc9612 (
      {stage2_47[101]},
      {stage3_47[67]}
   );
   gpc1_1 gpc9613 (
      {stage2_47[102]},
      {stage3_47[68]}
   );
   gpc1_1 gpc9614 (
      {stage2_47[103]},
      {stage3_47[69]}
   );
   gpc1_1 gpc9615 (
      {stage2_47[104]},
      {stage3_47[70]}
   );
   gpc1_1 gpc9616 (
      {stage2_47[105]},
      {stage3_47[71]}
   );
   gpc1_1 gpc9617 (
      {stage2_47[106]},
      {stage3_47[72]}
   );
   gpc1_1 gpc9618 (
      {stage2_47[107]},
      {stage3_47[73]}
   );
   gpc1_1 gpc9619 (
      {stage2_49[96]},
      {stage3_49[45]}
   );
   gpc1_1 gpc9620 (
      {stage2_49[97]},
      {stage3_49[46]}
   );
   gpc1_1 gpc9621 (
      {stage2_49[98]},
      {stage3_49[47]}
   );
   gpc1_1 gpc9622 (
      {stage2_49[99]},
      {stage3_49[48]}
   );
   gpc1_1 gpc9623 (
      {stage2_49[100]},
      {stage3_49[49]}
   );
   gpc1_1 gpc9624 (
      {stage2_49[101]},
      {stage3_49[50]}
   );
   gpc1_1 gpc9625 (
      {stage2_49[102]},
      {stage3_49[51]}
   );
   gpc1_1 gpc9626 (
      {stage2_49[103]},
      {stage3_49[52]}
   );
   gpc1_1 gpc9627 (
      {stage2_49[104]},
      {stage3_49[53]}
   );
   gpc1_1 gpc9628 (
      {stage2_49[105]},
      {stage3_49[54]}
   );
   gpc1_1 gpc9629 (
      {stage2_49[106]},
      {stage3_49[55]}
   );
   gpc1_1 gpc9630 (
      {stage2_49[107]},
      {stage3_49[56]}
   );
   gpc1_1 gpc9631 (
      {stage2_49[108]},
      {stage3_49[57]}
   );
   gpc1_1 gpc9632 (
      {stage2_49[109]},
      {stage3_49[58]}
   );
   gpc1_1 gpc9633 (
      {stage2_49[110]},
      {stage3_49[59]}
   );
   gpc1_1 gpc9634 (
      {stage2_49[111]},
      {stage3_49[60]}
   );
   gpc1_1 gpc9635 (
      {stage2_49[112]},
      {stage3_49[61]}
   );
   gpc1_1 gpc9636 (
      {stage2_49[113]},
      {stage3_49[62]}
   );
   gpc1_1 gpc9637 (
      {stage2_49[114]},
      {stage3_49[63]}
   );
   gpc1_1 gpc9638 (
      {stage2_49[115]},
      {stage3_49[64]}
   );
   gpc1_1 gpc9639 (
      {stage2_50[149]},
      {stage3_50[60]}
   );
   gpc1_1 gpc9640 (
      {stage2_50[150]},
      {stage3_50[61]}
   );
   gpc1_1 gpc9641 (
      {stage2_50[151]},
      {stage3_50[62]}
   );
   gpc1_1 gpc9642 (
      {stage2_50[152]},
      {stage3_50[63]}
   );
   gpc1_1 gpc9643 (
      {stage2_51[81]},
      {stage3_51[47]}
   );
   gpc1_1 gpc9644 (
      {stage2_51[82]},
      {stage3_51[48]}
   );
   gpc1_1 gpc9645 (
      {stage2_51[83]},
      {stage3_51[49]}
   );
   gpc1_1 gpc9646 (
      {stage2_51[84]},
      {stage3_51[50]}
   );
   gpc1_1 gpc9647 (
      {stage2_51[85]},
      {stage3_51[51]}
   );
   gpc1_1 gpc9648 (
      {stage2_51[86]},
      {stage3_51[52]}
   );
   gpc1_1 gpc9649 (
      {stage2_51[87]},
      {stage3_51[53]}
   );
   gpc1_1 gpc9650 (
      {stage2_52[109]},
      {stage3_52[37]}
   );
   gpc1_1 gpc9651 (
      {stage2_52[110]},
      {stage3_52[38]}
   );
   gpc1_1 gpc9652 (
      {stage2_52[111]},
      {stage3_52[39]}
   );
   gpc1_1 gpc9653 (
      {stage2_52[112]},
      {stage3_52[40]}
   );
   gpc1_1 gpc9654 (
      {stage2_52[113]},
      {stage3_52[41]}
   );
   gpc1_1 gpc9655 (
      {stage2_52[114]},
      {stage3_52[42]}
   );
   gpc1_1 gpc9656 (
      {stage2_52[115]},
      {stage3_52[43]}
   );
   gpc1_1 gpc9657 (
      {stage2_52[116]},
      {stage3_52[44]}
   );
   gpc1_1 gpc9658 (
      {stage2_52[117]},
      {stage3_52[45]}
   );
   gpc1_1 gpc9659 (
      {stage2_52[118]},
      {stage3_52[46]}
   );
   gpc1_1 gpc9660 (
      {stage2_52[119]},
      {stage3_52[47]}
   );
   gpc1_1 gpc9661 (
      {stage2_52[120]},
      {stage3_52[48]}
   );
   gpc1_1 gpc9662 (
      {stage2_52[121]},
      {stage3_52[49]}
   );
   gpc1_1 gpc9663 (
      {stage2_52[122]},
      {stage3_52[50]}
   );
   gpc1_1 gpc9664 (
      {stage2_52[123]},
      {stage3_52[51]}
   );
   gpc1_1 gpc9665 (
      {stage2_52[124]},
      {stage3_52[52]}
   );
   gpc1_1 gpc9666 (
      {stage2_52[125]},
      {stage3_52[53]}
   );
   gpc1_1 gpc9667 (
      {stage2_52[126]},
      {stage3_52[54]}
   );
   gpc1_1 gpc9668 (
      {stage2_52[127]},
      {stage3_52[55]}
   );
   gpc1_1 gpc9669 (
      {stage2_53[89]},
      {stage3_53[45]}
   );
   gpc1_1 gpc9670 (
      {stage2_53[90]},
      {stage3_53[46]}
   );
   gpc1_1 gpc9671 (
      {stage2_53[91]},
      {stage3_53[47]}
   );
   gpc1_1 gpc9672 (
      {stage2_53[92]},
      {stage3_53[48]}
   );
   gpc1_1 gpc9673 (
      {stage2_53[93]},
      {stage3_53[49]}
   );
   gpc1_1 gpc9674 (
      {stage2_53[94]},
      {stage3_53[50]}
   );
   gpc1_1 gpc9675 (
      {stage2_53[95]},
      {stage3_53[51]}
   );
   gpc1_1 gpc9676 (
      {stage2_53[96]},
      {stage3_53[52]}
   );
   gpc1_1 gpc9677 (
      {stage2_54[114]},
      {stage3_54[53]}
   );
   gpc1_1 gpc9678 (
      {stage2_54[115]},
      {stage3_54[54]}
   );
   gpc1_1 gpc9679 (
      {stage2_54[116]},
      {stage3_54[55]}
   );
   gpc1_1 gpc9680 (
      {stage2_54[117]},
      {stage3_54[56]}
   );
   gpc1_1 gpc9681 (
      {stage2_54[118]},
      {stage3_54[57]}
   );
   gpc1_1 gpc9682 (
      {stage2_54[119]},
      {stage3_54[58]}
   );
   gpc1_1 gpc9683 (
      {stage2_54[120]},
      {stage3_54[59]}
   );
   gpc1_1 gpc9684 (
      {stage2_54[121]},
      {stage3_54[60]}
   );
   gpc1_1 gpc9685 (
      {stage2_54[122]},
      {stage3_54[61]}
   );
   gpc1_1 gpc9686 (
      {stage2_54[123]},
      {stage3_54[62]}
   );
   gpc1_1 gpc9687 (
      {stage2_55[102]},
      {stage3_55[38]}
   );
   gpc1_1 gpc9688 (
      {stage2_55[103]},
      {stage3_55[39]}
   );
   gpc1_1 gpc9689 (
      {stage2_55[104]},
      {stage3_55[40]}
   );
   gpc1_1 gpc9690 (
      {stage2_55[105]},
      {stage3_55[41]}
   );
   gpc1_1 gpc9691 (
      {stage2_55[106]},
      {stage3_55[42]}
   );
   gpc1_1 gpc9692 (
      {stage2_55[107]},
      {stage3_55[43]}
   );
   gpc1_1 gpc9693 (
      {stage2_55[108]},
      {stage3_55[44]}
   );
   gpc1_1 gpc9694 (
      {stage2_55[109]},
      {stage3_55[45]}
   );
   gpc1_1 gpc9695 (
      {stage2_55[110]},
      {stage3_55[46]}
   );
   gpc1_1 gpc9696 (
      {stage2_57[72]},
      {stage3_57[46]}
   );
   gpc1_1 gpc9697 (
      {stage2_57[73]},
      {stage3_57[47]}
   );
   gpc1_1 gpc9698 (
      {stage2_57[74]},
      {stage3_57[48]}
   );
   gpc1_1 gpc9699 (
      {stage2_57[75]},
      {stage3_57[49]}
   );
   gpc1_1 gpc9700 (
      {stage2_57[76]},
      {stage3_57[50]}
   );
   gpc1_1 gpc9701 (
      {stage2_57[77]},
      {stage3_57[51]}
   );
   gpc1_1 gpc9702 (
      {stage2_57[78]},
      {stage3_57[52]}
   );
   gpc1_1 gpc9703 (
      {stage2_58[79]},
      {stage3_58[43]}
   );
   gpc1_1 gpc9704 (
      {stage2_58[80]},
      {stage3_58[44]}
   );
   gpc1_1 gpc9705 (
      {stage2_58[81]},
      {stage3_58[45]}
   );
   gpc1_1 gpc9706 (
      {stage2_58[82]},
      {stage3_58[46]}
   );
   gpc1_1 gpc9707 (
      {stage2_58[83]},
      {stage3_58[47]}
   );
   gpc1_1 gpc9708 (
      {stage2_58[84]},
      {stage3_58[48]}
   );
   gpc1_1 gpc9709 (
      {stage2_59[133]},
      {stage3_59[39]}
   );
   gpc1_1 gpc9710 (
      {stage2_59[134]},
      {stage3_59[40]}
   );
   gpc1_1 gpc9711 (
      {stage2_59[135]},
      {stage3_59[41]}
   );
   gpc1_1 gpc9712 (
      {stage2_59[136]},
      {stage3_59[42]}
   );
   gpc1_1 gpc9713 (
      {stage2_59[137]},
      {stage3_59[43]}
   );
   gpc1_1 gpc9714 (
      {stage2_59[138]},
      {stage3_59[44]}
   );
   gpc1_1 gpc9715 (
      {stage2_59[139]},
      {stage3_59[45]}
   );
   gpc1_1 gpc9716 (
      {stage2_60[106]},
      {stage3_60[48]}
   );
   gpc1_1 gpc9717 (
      {stage2_60[107]},
      {stage3_60[49]}
   );
   gpc1_1 gpc9718 (
      {stage2_60[108]},
      {stage3_60[50]}
   );
   gpc1_1 gpc9719 (
      {stage2_60[109]},
      {stage3_60[51]}
   );
   gpc1_1 gpc9720 (
      {stage2_60[110]},
      {stage3_60[52]}
   );
   gpc1_1 gpc9721 (
      {stage2_61[90]},
      {stage3_61[45]}
   );
   gpc1_1 gpc9722 (
      {stage2_61[91]},
      {stage3_61[46]}
   );
   gpc1_1 gpc9723 (
      {stage2_61[92]},
      {stage3_61[47]}
   );
   gpc1_1 gpc9724 (
      {stage2_61[93]},
      {stage3_61[48]}
   );
   gpc1_1 gpc9725 (
      {stage2_61[94]},
      {stage3_61[49]}
   );
   gpc1_1 gpc9726 (
      {stage2_61[95]},
      {stage3_61[50]}
   );
   gpc1_1 gpc9727 (
      {stage2_61[96]},
      {stage3_61[51]}
   );
   gpc1_1 gpc9728 (
      {stage2_61[97]},
      {stage3_61[52]}
   );
   gpc1_1 gpc9729 (
      {stage2_61[98]},
      {stage3_61[53]}
   );
   gpc1_1 gpc9730 (
      {stage2_61[99]},
      {stage3_61[54]}
   );
   gpc1_1 gpc9731 (
      {stage2_61[100]},
      {stage3_61[55]}
   );
   gpc1_1 gpc9732 (
      {stage2_61[101]},
      {stage3_61[56]}
   );
   gpc1_1 gpc9733 (
      {stage2_62[144]},
      {stage3_62[40]}
   );
   gpc1_1 gpc9734 (
      {stage2_63[95]},
      {stage3_63[54]}
   );
   gpc1_1 gpc9735 (
      {stage2_63[96]},
      {stage3_63[55]}
   );
   gpc1_1 gpc9736 (
      {stage2_63[97]},
      {stage3_63[56]}
   );
   gpc1_1 gpc9737 (
      {stage2_63[98]},
      {stage3_63[57]}
   );
   gpc1_1 gpc9738 (
      {stage2_63[99]},
      {stage3_63[58]}
   );
   gpc1_1 gpc9739 (
      {stage2_63[100]},
      {stage3_63[59]}
   );
   gpc1_1 gpc9740 (
      {stage2_63[101]},
      {stage3_63[60]}
   );
   gpc1_1 gpc9741 (
      {stage2_63[102]},
      {stage3_63[61]}
   );
   gpc1_1 gpc9742 (
      {stage2_63[103]},
      {stage3_63[62]}
   );
   gpc1_1 gpc9743 (
      {stage2_63[104]},
      {stage3_63[63]}
   );
   gpc1_1 gpc9744 (
      {stage2_63[105]},
      {stage3_63[64]}
   );
   gpc1_1 gpc9745 (
      {stage2_63[106]},
      {stage3_63[65]}
   );
   gpc1_1 gpc9746 (
      {stage2_63[107]},
      {stage3_63[66]}
   );
   gpc1_1 gpc9747 (
      {stage2_63[108]},
      {stage3_63[67]}
   );
   gpc1_1 gpc9748 (
      {stage2_63[109]},
      {stage3_63[68]}
   );
   gpc1_1 gpc9749 (
      {stage2_63[110]},
      {stage3_63[69]}
   );
   gpc1_1 gpc9750 (
      {stage2_63[111]},
      {stage3_63[70]}
   );
   gpc1_1 gpc9751 (
      {stage2_63[112]},
      {stage3_63[71]}
   );
   gpc1_1 gpc9752 (
      {stage2_64[95]},
      {stage3_64[44]}
   );
   gpc1_1 gpc9753 (
      {stage2_64[96]},
      {stage3_64[45]}
   );
   gpc1_1 gpc9754 (
      {stage2_64[97]},
      {stage3_64[46]}
   );
   gpc1_1 gpc9755 (
      {stage2_64[98]},
      {stage3_64[47]}
   );
   gpc1_1 gpc9756 (
      {stage2_64[99]},
      {stage3_64[48]}
   );
   gpc1_1 gpc9757 (
      {stage2_64[100]},
      {stage3_64[49]}
   );
   gpc1_1 gpc9758 (
      {stage2_64[101]},
      {stage3_64[50]}
   );
   gpc1_1 gpc9759 (
      {stage2_65[65]},
      {stage3_65[30]}
   );
   gpc1_1 gpc9760 (
      {stage2_65[66]},
      {stage3_65[31]}
   );
   gpc1_1 gpc9761 (
      {stage2_65[67]},
      {stage3_65[32]}
   );
   gpc1_1 gpc9762 (
      {stage2_66[30]},
      {stage3_66[30]}
   );
   gpc1_1 gpc9763 (
      {stage2_66[31]},
      {stage3_66[31]}
   );
   gpc1_1 gpc9764 (
      {stage2_66[32]},
      {stage3_66[32]}
   );
   gpc1_1 gpc9765 (
      {stage2_66[33]},
      {stage3_66[33]}
   );
   gpc1_1 gpc9766 (
      {stage2_66[34]},
      {stage3_66[34]}
   );
   gpc1_1 gpc9767 (
      {stage2_66[35]},
      {stage3_66[35]}
   );
   gpc1_1 gpc9768 (
      {stage2_66[36]},
      {stage3_66[36]}
   );
   gpc1_1 gpc9769 (
      {stage2_66[37]},
      {stage3_66[37]}
   );
   gpc1_1 gpc9770 (
      {stage2_66[38]},
      {stage3_66[38]}
   );
   gpc1_1 gpc9771 (
      {stage2_66[39]},
      {stage3_66[39]}
   );
   gpc1_1 gpc9772 (
      {stage2_66[40]},
      {stage3_66[40]}
   );
   gpc1_1 gpc9773 (
      {stage2_66[41]},
      {stage3_66[41]}
   );
   gpc1_1 gpc9774 (
      {stage2_66[42]},
      {stage3_66[42]}
   );
   gpc1_1 gpc9775 (
      {stage2_66[43]},
      {stage3_66[43]}
   );
   gpc1_1 gpc9776 (
      {stage2_66[44]},
      {stage3_66[44]}
   );
   gpc1_1 gpc9777 (
      {stage2_66[45]},
      {stage3_66[45]}
   );
   gpc1_1 gpc9778 (
      {stage2_66[46]},
      {stage3_66[46]}
   );
   gpc1_1 gpc9779 (
      {stage2_66[47]},
      {stage3_66[47]}
   );
   gpc1_1 gpc9780 (
      {stage2_66[48]},
      {stage3_66[48]}
   );
   gpc1_1 gpc9781 (
      {stage2_66[49]},
      {stage3_66[49]}
   );
   gpc1_1 gpc9782 (
      {stage2_66[50]},
      {stage3_66[50]}
   );
   gpc1_1 gpc9783 (
      {stage2_66[51]},
      {stage3_66[51]}
   );
   gpc1_1 gpc9784 (
      {stage2_66[52]},
      {stage3_66[52]}
   );
   gpc1_1 gpc9785 (
      {stage2_66[53]},
      {stage3_66[53]}
   );
   gpc606_5 gpc9786 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc9787 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc9788 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc9789 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc9790 (
      {stage3_1[18], stage3_1[19], stage3_1[20], stage3_1[21], stage3_1[22], stage3_1[23]},
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc9791 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc9792 (
      {stage3_3[24], stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc9793 (
      {stage3_3[29], stage3_3[30], stage3_3[31], stage3_3[32], stage3_3[33]},
      {stage3_4[7]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc9794 (
      {stage3_3[34], stage3_3[35], stage3_3[36], stage3_3[37], stage3_3[38]},
      {stage3_4[8]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[3],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc9795 (
      {stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[4],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc9796 (
      {stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[5],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc9797 (
      {stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[5],stage4_6[6],stage4_5[10],stage4_4[11]}
   );
   gpc606_5 gpc9798 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[3],stage4_7[6],stage4_6[7],stage4_5[11],stage4_4[12]}
   );
   gpc606_5 gpc9799 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[4],stage4_7[7],stage4_6[8],stage4_5[12],stage4_4[13]}
   );
   gpc606_5 gpc9800 (
      {stage3_4[39], stage3_4[40], stage3_4[41], stage3_4[42], stage3_4[43], stage3_4[44]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[5],stage4_7[8],stage4_6[9],stage4_5[13],stage4_4[14]}
   );
   gpc606_5 gpc9801 (
      {stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48], stage3_4[49], stage3_4[50]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[6],stage4_7[9],stage4_6[10],stage4_5[14],stage4_4[15]}
   );
   gpc606_5 gpc9802 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[7],stage4_7[10],stage4_6[11],stage4_5[15]}
   );
   gpc615_5 gpc9803 (
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[8],stage4_7[11],stage4_6[12]}
   );
   gpc615_5 gpc9804 (
      {stage3_6[47], stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[9],stage4_7[12],stage4_6[13]}
   );
   gpc615_5 gpc9805 (
      {stage3_6[52], stage3_6[53], stage3_6[54], stage3_6[55], stage3_6[56]},
      {stage3_7[8]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[10],stage4_7[13],stage4_6[14]}
   );
   gpc615_5 gpc9806 (
      {stage3_6[57], stage3_6[58], stage3_6[59], stage3_6[60], stage3_6[61]},
      {stage3_7[9]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[4],stage4_8[11],stage4_7[14],stage4_6[15]}
   );
   gpc615_5 gpc9807 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[24]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[4],stage4_9[5],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc9808 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[25]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[5],stage4_9[6],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc9809 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[26]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[6],stage4_9[7],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc9810 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[27]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[7],stage4_9[8],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc9811 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[28]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[8],stage4_9[9],stage4_8[16],stage4_7[19]}
   );
   gpc606_5 gpc9812 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[5],stage4_10[9],stage4_9[10]}
   );
   gpc606_5 gpc9813 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[6],stage4_10[10],stage4_9[11]}
   );
   gpc606_5 gpc9814 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[7],stage4_10[11],stage4_9[12]}
   );
   gpc606_5 gpc9815 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], 1'b0},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[8],stage4_10[12],stage4_9[13]}
   );
   gpc615_5 gpc9816 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[24]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[4],stage4_12[4],stage4_11[9],stage4_10[13]}
   );
   gpc615_5 gpc9817 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[25]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[5],stage4_12[5],stage4_11[10],stage4_10[14]}
   );
   gpc615_5 gpc9818 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[26]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[6],stage4_12[6],stage4_11[11],stage4_10[15]}
   );
   gpc615_5 gpc9819 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[27]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[7],stage4_12[7],stage4_11[12],stage4_10[16]}
   );
   gpc615_5 gpc9820 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24]},
      {stage3_11[28]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[8],stage4_12[8],stage4_11[13],stage4_10[17]}
   );
   gpc615_5 gpc9821 (
      {stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29]},
      {stage3_11[29]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[9],stage4_12[9],stage4_11[14],stage4_10[18]}
   );
   gpc615_5 gpc9822 (
      {stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33], stage3_10[34]},
      {stage3_11[30]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[10],stage4_12[10],stage4_11[15],stage4_10[19]}
   );
   gpc615_5 gpc9823 (
      {stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38], stage3_10[39]},
      {stage3_11[31]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[11],stage4_12[11],stage4_11[16],stage4_10[20]}
   );
   gpc615_5 gpc9824 (
      {stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43], stage3_10[44]},
      {stage3_11[32]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[12],stage4_12[12],stage4_11[17],stage4_10[21]}
   );
   gpc615_5 gpc9825 (
      {stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48], stage3_10[49]},
      {stage3_11[33]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[13],stage4_12[13],stage4_11[18],stage4_10[22]}
   );
   gpc615_5 gpc9826 (
      {stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53], stage3_10[54]},
      {stage3_11[34]},
      {stage3_12[60], stage3_12[61], stage3_12[62], stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage4_14[10],stage4_13[14],stage4_12[14],stage4_11[19],stage4_10[23]}
   );
   gpc615_5 gpc9827 (
      {stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58], stage3_10[59]},
      {stage3_11[35]},
      {stage3_12[66], stage3_12[67], stage3_12[68], stage3_12[69], stage3_12[70], stage3_12[71]},
      {stage4_14[11],stage4_13[15],stage4_12[15],stage4_11[20],stage4_10[24]}
   );
   gpc615_5 gpc9828 (
      {stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63], stage3_10[64]},
      {stage3_11[36]},
      {stage3_12[72], stage3_12[73], stage3_12[74], stage3_12[75], stage3_12[76], stage3_12[77]},
      {stage4_14[12],stage4_13[16],stage4_12[16],stage4_11[21],stage4_10[25]}
   );
   gpc615_5 gpc9829 (
      {stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[78]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[13],stage4_13[17],stage4_12[17],stage4_11[22]}
   );
   gpc615_5 gpc9830 (
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46]},
      {stage3_12[79]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[14],stage4_13[18],stage4_12[18],stage4_11[23]}
   );
   gpc615_5 gpc9831 (
      {stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51]},
      {stage3_12[80]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[15],stage4_13[19],stage4_12[19],stage4_11[24]}
   );
   gpc117_4 gpc9832 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[3],stage4_14[16],stage4_13[20]}
   );
   gpc606_5 gpc9833 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6]},
      {stage4_17[0],stage4_16[1],stage4_15[4],stage4_14[17],stage4_13[21]}
   );
   gpc606_5 gpc9834 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage4_17[1],stage4_16[2],stage4_15[5],stage4_14[18],stage4_13[22]}
   );
   gpc606_5 gpc9835 (
      {stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42]},
      {stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18]},
      {stage4_17[2],stage4_16[3],stage4_15[6],stage4_14[19],stage4_13[23]}
   );
   gpc615_5 gpc9836 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_15[19]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[3],stage4_16[4],stage4_15[7],stage4_14[20]}
   );
   gpc615_5 gpc9837 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[20]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[4],stage4_16[5],stage4_15[8],stage4_14[21]}
   );
   gpc615_5 gpc9838 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[21]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[5],stage4_16[6],stage4_15[9],stage4_14[22]}
   );
   gpc615_5 gpc9839 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[22]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[6],stage4_16[7],stage4_15[10],stage4_14[23]}
   );
   gpc615_5 gpc9840 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[23]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[7],stage4_16[8],stage4_15[11],stage4_14[24]}
   );
   gpc615_5 gpc9841 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[24]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[8],stage4_16[9],stage4_15[12],stage4_14[25]}
   );
   gpc615_5 gpc9842 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[9],stage4_16[10],stage4_15[13]}
   );
   gpc615_5 gpc9843 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[37]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[7],stage4_17[10],stage4_16[11],stage4_15[14]}
   );
   gpc615_5 gpc9844 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[38]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[8],stage4_17[11],stage4_16[12],stage4_15[15]}
   );
   gpc615_5 gpc9845 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[39]},
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage4_19[3],stage4_18[9],stage4_17[12],stage4_16[13],stage4_15[16]}
   );
   gpc606_5 gpc9846 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[4],stage4_18[10],stage4_17[13]}
   );
   gpc606_5 gpc9847 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[5],stage4_18[11],stage4_17[14]}
   );
   gpc207_4 gpc9848 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[2],stage4_20[2],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc9849 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[3],stage4_20[3],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc9850 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[4],stage4_20[4],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc9851 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[5],stage4_20[5],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc9852 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[6],stage4_20[6],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc9853 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[7],stage4_20[7],stage4_19[11],stage4_18[17]}
   );
   gpc615_5 gpc9854 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46]},
      {stage3_19[12]},
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage4_22[0],stage4_21[8],stage4_20[8],stage4_19[12],stage4_18[18]}
   );
   gpc615_5 gpc9855 (
      {stage3_18[47], stage3_18[48], stage3_18[49], stage3_18[50], stage3_18[51]},
      {stage3_19[13]},
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage4_22[1],stage4_21[9],stage4_20[9],stage4_19[13],stage4_18[19]}
   );
   gpc606_5 gpc9856 (
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[2],stage4_21[10],stage4_20[10],stage4_19[14]}
   );
   gpc606_5 gpc9857 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[3],stage4_21[11],stage4_20[11],stage4_19[15]}
   );
   gpc615_5 gpc9858 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[24]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[4],stage4_21[12],stage4_20[12],stage4_19[16]}
   );
   gpc615_5 gpc9859 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35]},
      {stage3_20[25]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[5],stage4_21[13],stage4_20[13],stage4_19[17]}
   );
   gpc615_5 gpc9860 (
      {stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40]},
      {stage3_20[26]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[6],stage4_21[14],stage4_20[14],stage4_19[18]}
   );
   gpc615_5 gpc9861 (
      {stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45]},
      {stage3_20[27]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[7],stage4_21[15],stage4_20[15],stage4_19[19]}
   );
   gpc606_5 gpc9862 (
      {stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31], stage3_20[32], stage3_20[33]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[6],stage4_22[8],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc9863 (
      {stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37], stage3_20[38], stage3_20[39]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[7],stage4_22[9],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc9864 (
      {stage3_20[40], stage3_20[41], stage3_20[42], stage3_20[43], stage3_20[44], stage3_20[45]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[8],stage4_22[10],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc9865 (
      {stage3_20[46], stage3_20[47], stage3_20[48], stage3_20[49], stage3_20[50], stage3_20[51]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[9],stage4_22[11],stage4_21[19],stage4_20[19]}
   );
   gpc615_5 gpc9866 (
      {stage3_20[52], stage3_20[53], stage3_20[54], stage3_20[55], stage3_20[56]},
      {stage3_21[36]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[10],stage4_22[12],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc9867 (
      {stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[5],stage4_23[11],stage4_22[13],stage4_21[21]}
   );
   gpc606_5 gpc9868 (
      {stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[6],stage4_23[12],stage4_22[14],stage4_21[22]}
   );
   gpc606_5 gpc9869 (
      {stage3_21[49], stage3_21[50], stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[7],stage4_23[13],stage4_22[15],stage4_21[23]}
   );
   gpc606_5 gpc9870 (
      {stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59], stage3_21[60]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[8],stage4_23[14],stage4_22[16],stage4_21[24]}
   );
   gpc615_5 gpc9871 (
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[9],stage4_23[15],stage4_22[17]}
   );
   gpc615_5 gpc9872 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[10],stage4_23[16],stage4_22[18]}
   );
   gpc615_5 gpc9873 (
      {stage3_22[40], stage3_22[41], stage3_22[42], stage3_22[43], stage3_22[44]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[11],stage4_23[17],stage4_22[19]}
   );
   gpc615_5 gpc9874 (
      {stage3_22[45], stage3_22[46], stage3_22[47], stage3_22[48], stage3_22[49]},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[12],stage4_23[18],stage4_22[20]}
   );
   gpc615_5 gpc9875 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[13],stage4_23[19]}
   );
   gpc615_5 gpc9876 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[14],stage4_23[20]}
   );
   gpc615_5 gpc9877 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[15],stage4_23[21]}
   );
   gpc615_5 gpc9878 (
      {stage3_23[43], stage3_23[44], stage3_23[45], stage3_23[46], stage3_23[47]},
      {stage3_24[27]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[7],stage4_25[11],stage4_24[16],stage4_23[22]}
   );
   gpc615_5 gpc9879 (
      {stage3_23[48], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_24[28]},
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage4_27[4],stage4_26[8],stage4_25[12],stage4_24[17],stage4_23[23]}
   );
   gpc606_5 gpc9880 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[5],stage4_26[9],stage4_25[13]}
   );
   gpc606_5 gpc9881 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[6],stage4_26[10],stage4_25[14]}
   );
   gpc606_5 gpc9882 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46], stage3_25[47]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[7],stage4_26[11],stage4_25[15]}
   );
   gpc606_5 gpc9883 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[3],stage4_28[3],stage4_27[8],stage4_26[12]}
   );
   gpc606_5 gpc9884 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[4],stage4_28[4],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc9885 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[5],stage4_28[5],stage4_27[10],stage4_26[14]}
   );
   gpc606_5 gpc9886 (
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[6],stage4_28[6],stage4_27[11],stage4_26[15]}
   );
   gpc606_5 gpc9887 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage4_30[4],stage4_29[7],stage4_28[7],stage4_27[12],stage4_26[16]}
   );
   gpc606_5 gpc9888 (
      {stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage4_30[5],stage4_29[8],stage4_28[8],stage4_27[13],stage4_26[17]}
   );
   gpc606_5 gpc9889 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40], stage3_26[41]},
      {stage3_28[36], stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41]},
      {stage4_30[6],stage4_29[9],stage4_28[9],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc9890 (
      {stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47]},
      {stage3_28[42], stage3_28[43], stage3_28[44], stage3_28[45], stage3_28[46], stage3_28[47]},
      {stage4_30[7],stage4_29[10],stage4_28[10],stage4_27[15],stage4_26[19]}
   );
   gpc606_5 gpc9891 (
      {stage3_26[48], stage3_26[49], stage3_26[50], stage3_26[51], 1'b0, 1'b0},
      {stage3_28[48], stage3_28[49], stage3_28[50], stage3_28[51], stage3_28[52], stage3_28[53]},
      {stage4_30[8],stage4_29[11],stage4_28[11],stage4_27[16],stage4_26[20]}
   );
   gpc606_5 gpc9892 (
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[9],stage4_29[12],stage4_28[12],stage4_27[17]}
   );
   gpc606_5 gpc9893 (
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[10],stage4_29[13],stage4_28[13],stage4_27[18]}
   );
   gpc606_5 gpc9894 (
      {stage3_27[30], stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[11],stage4_29[14],stage4_28[14],stage4_27[19]}
   );
   gpc606_5 gpc9895 (
      {stage3_27[36], stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[12],stage4_29[15],stage4_28[15],stage4_27[20]}
   );
   gpc1163_5 gpc9896 (
      {stage3_29[24], stage3_29[25], stage3_29[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[4],stage4_30[13],stage4_29[16]}
   );
   gpc1163_5 gpc9897 (
      {stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[5],stage4_30[14],stage4_29[17]}
   );
   gpc1163_5 gpc9898 (
      {stage3_29[30], stage3_29[31], stage3_29[32]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[6],stage4_30[15],stage4_29[18]}
   );
   gpc1163_5 gpc9899 (
      {stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[7],stage4_30[16],stage4_29[19]}
   );
   gpc606_5 gpc9900 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[4],stage4_32[4],stage4_31[8],stage4_30[17],stage4_29[20]}
   );
   gpc606_5 gpc9901 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15]},
      {stage4_33[5],stage4_32[5],stage4_31[9],stage4_30[18],stage4_29[21]}
   );
   gpc606_5 gpc9902 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52], stage3_29[53]},
      {stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21]},
      {stage4_33[6],stage4_32[6],stage4_31[10],stage4_30[19],stage4_29[22]}
   );
   gpc606_5 gpc9903 (
      {stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57], stage3_29[58], 1'b0},
      {stage3_31[22], stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage4_33[7],stage4_32[7],stage4_31[11],stage4_30[20],stage4_29[23]}
   );
   gpc606_5 gpc9904 (
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_32[4], stage3_32[5], stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9]},
      {stage4_34[0],stage4_33[8],stage4_32[8],stage4_31[12],stage4_30[21]}
   );
   gpc606_5 gpc9905 (
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage4_34[1],stage4_33[9],stage4_32[9],stage4_31[13],stage4_30[22]}
   );
   gpc615_5 gpc9906 (
      {stage3_31[28], stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32]},
      {stage3_32[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[10],stage4_32[10],stage4_31[14]}
   );
   gpc615_5 gpc9907 (
      {stage3_31[33], stage3_31[34], stage3_31[35], stage3_31[36], stage3_31[37]},
      {stage3_32[17]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[11],stage4_32[11],stage4_31[15]}
   );
   gpc615_5 gpc9908 (
      {stage3_31[38], stage3_31[39], stage3_31[40], stage3_31[41], 1'b0},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[12],stage4_32[12],stage4_31[16]}
   );
   gpc2116_5 gpc9909 (
      {stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24]},
      {stage3_33[18]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[13],stage4_32[13]}
   );
   gpc2116_5 gpc9910 (
      {stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[19]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc9911 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[20]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc9912 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[21]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[16],stage4_32[16]}
   );
   gpc615_5 gpc9913 (
      {stage3_32[41], stage3_32[42], stage3_32[43], stage3_32[44], stage3_32[45]},
      {stage3_33[22]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[17],stage4_32[17]}
   );
   gpc615_5 gpc9914 (
      {stage3_32[46], stage3_32[47], stage3_32[48], stage3_32[49], stage3_32[50]},
      {stage3_33[23]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[8],stage4_34[10],stage4_33[18],stage4_32[18]}
   );
   gpc215_4 gpc9915 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28]},
      {stage3_34[26]},
      {stage3_35[4], stage3_35[5]},
      {stage4_36[6],stage4_35[9],stage4_34[11],stage4_33[19]}
   );
   gpc606_5 gpc9916 (
      {stage3_33[29], stage3_33[30], stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[7],stage4_35[10],stage4_34[12],stage4_33[20]}
   );
   gpc606_5 gpc9917 (
      {stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38], stage3_33[39], stage3_33[40]},
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage4_37[1],stage4_36[8],stage4_35[11],stage4_34[13],stage4_33[21]}
   );
   gpc606_5 gpc9918 (
      {stage3_33[41], stage3_33[42], stage3_33[43], stage3_33[44], stage3_33[45], stage3_33[46]},
      {stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage4_37[2],stage4_36[9],stage4_35[12],stage4_34[14],stage4_33[22]}
   );
   gpc606_5 gpc9919 (
      {stage3_33[47], stage3_33[48], stage3_33[49], stage3_33[50], stage3_33[51], stage3_33[52]},
      {stage3_35[24], stage3_35[25], stage3_35[26], stage3_35[27], stage3_35[28], stage3_35[29]},
      {stage4_37[3],stage4_36[10],stage4_35[13],stage4_34[15],stage4_33[23]}
   );
   gpc615_5 gpc9920 (
      {stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage3_35[30]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage4_38[0],stage4_37[4],stage4_36[11],stage4_35[14],stage4_34[16]}
   );
   gpc606_5 gpc9921 (
      {stage3_35[31], stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[1],stage4_37[5],stage4_36[12],stage4_35[15]}
   );
   gpc615_5 gpc9922 (
      {stage3_35[37], stage3_35[38], stage3_35[39], stage3_35[40], stage3_35[41]},
      {stage3_36[6]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[2],stage4_37[6],stage4_36[13],stage4_35[16]}
   );
   gpc615_5 gpc9923 (
      {stage3_35[42], stage3_35[43], stage3_35[44], stage3_35[45], stage3_35[46]},
      {stage3_36[7]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[3],stage4_37[7],stage4_36[14],stage4_35[17]}
   );
   gpc615_5 gpc9924 (
      {stage3_35[47], stage3_35[48], stage3_35[49], stage3_35[50], stage3_35[51]},
      {stage3_36[8]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[4],stage4_37[8],stage4_36[15],stage4_35[18]}
   );
   gpc606_5 gpc9925 (
      {stage3_36[9], stage3_36[10], stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[4],stage4_38[5],stage4_37[9],stage4_36[16]}
   );
   gpc606_5 gpc9926 (
      {stage3_36[15], stage3_36[16], stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[5],stage4_38[6],stage4_37[10],stage4_36[17]}
   );
   gpc606_5 gpc9927 (
      {stage3_36[21], stage3_36[22], stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[6],stage4_38[7],stage4_37[11],stage4_36[18]}
   );
   gpc606_5 gpc9928 (
      {stage3_36[27], stage3_36[28], stage3_36[29], stage3_36[30], stage3_36[31], stage3_36[32]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[7],stage4_38[8],stage4_37[12],stage4_36[19]}
   );
   gpc606_5 gpc9929 (
      {stage3_36[33], stage3_36[34], stage3_36[35], stage3_36[36], stage3_36[37], stage3_36[38]},
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28], stage3_38[29]},
      {stage4_40[4],stage4_39[8],stage4_38[9],stage4_37[13],stage4_36[20]}
   );
   gpc606_5 gpc9930 (
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[5],stage4_39[9],stage4_38[10],stage4_37[14]}
   );
   gpc606_5 gpc9931 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], 1'b0},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[6],stage4_39[10],stage4_38[11],stage4_37[15]}
   );
   gpc615_5 gpc9932 (
      {stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33], stage3_38[34]},
      {stage3_39[12]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[2],stage4_40[7],stage4_39[11],stage4_38[12]}
   );
   gpc615_5 gpc9933 (
      {stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38], stage3_38[39]},
      {stage3_39[13]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[3],stage4_40[8],stage4_39[12],stage4_38[13]}
   );
   gpc615_5 gpc9934 (
      {stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43], stage3_38[44]},
      {stage3_39[14]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[4],stage4_40[9],stage4_39[13],stage4_38[14]}
   );
   gpc615_5 gpc9935 (
      {stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48], stage3_38[49]},
      {stage3_39[15]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[5],stage4_40[10],stage4_39[14],stage4_38[15]}
   );
   gpc615_5 gpc9936 (
      {stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53], stage3_38[54]},
      {stage3_39[16]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[6],stage4_40[11],stage4_39[15],stage4_38[16]}
   );
   gpc615_5 gpc9937 (
      {stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58], stage3_38[59]},
      {stage3_39[17]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[7],stage4_40[12],stage4_39[16],stage4_38[17]}
   );
   gpc207_4 gpc9938 (
      {stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22], stage3_39[23], stage3_39[24]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[6],stage4_41[8],stage4_40[13],stage4_39[17]}
   );
   gpc207_4 gpc9939 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[7],stage4_41[9],stage4_40[14],stage4_39[18]}
   );
   gpc207_4 gpc9940 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[8],stage4_41[10],stage4_40[15],stage4_39[19]}
   );
   gpc207_4 gpc9941 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[9],stage4_41[11],stage4_40[16],stage4_39[20]}
   );
   gpc207_4 gpc9942 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[8], stage3_41[9]},
      {stage4_42[10],stage4_41[12],stage4_40[17],stage4_39[21]}
   );
   gpc207_4 gpc9943 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57], stage3_39[58], stage3_39[59]},
      {stage3_41[10], stage3_41[11]},
      {stage4_42[11],stage4_41[13],stage4_40[18],stage4_39[22]}
   );
   gpc606_5 gpc9944 (
      {stage3_41[12], stage3_41[13], stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[12],stage4_41[14]}
   );
   gpc606_5 gpc9945 (
      {stage3_41[18], stage3_41[19], stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[13],stage4_41[15]}
   );
   gpc606_5 gpc9946 (
      {stage3_41[24], stage3_41[25], stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[14],stage4_41[16]}
   );
   gpc606_5 gpc9947 (
      {stage3_41[30], stage3_41[31], stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[15],stage4_41[17]}
   );
   gpc606_5 gpc9948 (
      {stage3_41[36], stage3_41[37], stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41]},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[16],stage4_41[18]}
   );
   gpc606_5 gpc9949 (
      {stage3_41[42], stage3_41[43], stage3_41[44], stage3_41[45], stage3_41[46], stage3_41[47]},
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[17],stage4_41[19]}
   );
   gpc606_5 gpc9950 (
      {stage3_41[48], stage3_41[49], stage3_41[50], stage3_41[51], stage3_41[52], stage3_41[53]},
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage4_45[6],stage4_44[6],stage4_43[6],stage4_42[18],stage4_41[20]}
   );
   gpc207_4 gpc9951 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[7],stage4_44[7],stage4_43[7],stage4_42[19]}
   );
   gpc207_4 gpc9952 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[8],stage4_44[8],stage4_43[8],stage4_42[20]}
   );
   gpc615_5 gpc9953 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18]},
      {stage3_43[42]},
      {stage3_44[4], stage3_44[5], stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[9],stage4_42[21]}
   );
   gpc615_5 gpc9954 (
      {stage3_42[19], stage3_42[20], stage3_42[21], stage3_42[22], stage3_42[23]},
      {stage3_43[43]},
      {stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[10],stage4_42[22]}
   );
   gpc615_5 gpc9955 (
      {stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27], stage3_42[28]},
      {stage3_43[44]},
      {stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21]},
      {stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[11],stage4_42[23]}
   );
   gpc615_5 gpc9956 (
      {stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_43[45]},
      {stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26], stage3_44[27]},
      {stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[12],stage4_42[24]}
   );
   gpc615_5 gpc9957 (
      {stage3_42[34], stage3_42[35], stage3_42[36], stage3_42[37], stage3_42[38]},
      {stage3_43[46]},
      {stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31], stage3_44[32], stage3_44[33]},
      {stage4_46[4],stage4_45[13],stage4_44[13],stage4_43[13],stage4_42[25]}
   );
   gpc615_5 gpc9958 (
      {stage3_42[39], stage3_42[40], stage3_42[41], stage3_42[42], stage3_42[43]},
      {stage3_43[47]},
      {stage3_44[34], stage3_44[35], stage3_44[36], stage3_44[37], stage3_44[38], stage3_44[39]},
      {stage4_46[5],stage4_45[14],stage4_44[14],stage4_43[14],stage4_42[26]}
   );
   gpc615_5 gpc9959 (
      {stage3_42[44], stage3_42[45], stage3_42[46], stage3_42[47], stage3_42[48]},
      {stage3_43[48]},
      {stage3_44[40], stage3_44[41], stage3_44[42], stage3_44[43], stage3_44[44], stage3_44[45]},
      {stage4_46[6],stage4_45[15],stage4_44[15],stage4_43[15],stage4_42[27]}
   );
   gpc615_5 gpc9960 (
      {stage3_42[49], stage3_42[50], stage3_42[51], stage3_42[52], stage3_42[53]},
      {stage3_43[49]},
      {stage3_44[46], stage3_44[47], stage3_44[48], stage3_44[49], stage3_44[50], stage3_44[51]},
      {stage4_46[7],stage4_45[16],stage4_44[16],stage4_43[16],stage4_42[28]}
   );
   gpc615_5 gpc9961 (
      {stage3_43[50], stage3_43[51], stage3_43[52], stage3_43[53], stage3_43[54]},
      {stage3_44[52]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[8],stage4_45[17],stage4_44[17],stage4_43[17]}
   );
   gpc1343_5 gpc9962 (
      {stage3_44[53], stage3_44[54], stage3_44[55]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[1],stage4_46[9],stage4_45[18],stage4_44[18]}
   );
   gpc1343_5 gpc9963 (
      {stage3_44[56], stage3_44[57], stage3_44[58]},
      {stage3_45[10], stage3_45[11], stage3_45[12], stage3_45[13]},
      {stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[1]},
      {stage4_48[1],stage4_47[2],stage4_46[10],stage4_45[19],stage4_44[19]}
   );
   gpc1343_5 gpc9964 (
      {stage3_44[59], stage3_44[60], stage3_44[61]},
      {stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_46[6], stage3_46[7], stage3_46[8]},
      {stage3_47[2]},
      {stage4_48[2],stage4_47[3],stage4_46[11],stage4_45[20],stage4_44[20]}
   );
   gpc623_5 gpc9965 (
      {stage3_44[62], stage3_44[63], stage3_44[64]},
      {stage3_45[18], stage3_45[19]},
      {stage3_46[9], stage3_46[10], stage3_46[11], stage3_46[12], stage3_46[13], stage3_46[14]},
      {stage4_48[3],stage4_47[4],stage4_46[12],stage4_45[21],stage4_44[21]}
   );
   gpc623_5 gpc9966 (
      {stage3_44[65], stage3_44[66], stage3_44[67]},
      {stage3_45[20], stage3_45[21]},
      {stage3_46[15], stage3_46[16], stage3_46[17], stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage4_48[4],stage4_47[5],stage4_46[13],stage4_45[22],stage4_44[22]}
   );
   gpc606_5 gpc9967 (
      {stage3_45[22], stage3_45[23], stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27]},
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8]},
      {stage4_49[0],stage4_48[5],stage4_47[6],stage4_46[14],stage4_45[23]}
   );
   gpc606_5 gpc9968 (
      {stage3_45[28], stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage4_49[1],stage4_48[6],stage4_47[7],stage4_46[15],stage4_45[24]}
   );
   gpc606_5 gpc9969 (
      {stage3_45[34], stage3_45[35], stage3_45[36], stage3_45[37], stage3_45[38], stage3_45[39]},
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage4_49[2],stage4_48[7],stage4_47[8],stage4_46[16],stage4_45[25]}
   );
   gpc615_5 gpc9970 (
      {stage3_46[21], stage3_46[22], stage3_46[23], stage3_46[24], stage3_46[25]},
      {stage3_47[21]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[3],stage4_48[8],stage4_47[9],stage4_46[17]}
   );
   gpc615_5 gpc9971 (
      {stage3_46[26], stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30]},
      {stage3_47[22]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[4],stage4_48[9],stage4_47[10],stage4_46[18]}
   );
   gpc615_5 gpc9972 (
      {stage3_46[31], stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35]},
      {stage3_47[23]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[5],stage4_48[10],stage4_47[11],stage4_46[19]}
   );
   gpc615_5 gpc9973 (
      {stage3_46[36], stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40]},
      {stage3_47[24]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[6],stage4_48[11],stage4_47[12],stage4_46[20]}
   );
   gpc615_5 gpc9974 (
      {stage3_46[41], stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45]},
      {stage3_47[25]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[7],stage4_48[12],stage4_47[13],stage4_46[21]}
   );
   gpc615_5 gpc9975 (
      {stage3_47[26], stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30]},
      {stage3_48[30]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[5],stage4_49[8],stage4_48[13],stage4_47[14]}
   );
   gpc615_5 gpc9976 (
      {stage3_47[31], stage3_47[32], stage3_47[33], stage3_47[34], stage3_47[35]},
      {stage3_48[31]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[6],stage4_49[9],stage4_48[14],stage4_47[15]}
   );
   gpc615_5 gpc9977 (
      {stage3_47[36], stage3_47[37], stage3_47[38], stage3_47[39], stage3_47[40]},
      {stage3_48[32]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[7],stage4_49[10],stage4_48[15],stage4_47[16]}
   );
   gpc615_5 gpc9978 (
      {stage3_47[41], stage3_47[42], stage3_47[43], stage3_47[44], stage3_47[45]},
      {stage3_48[33]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[8],stage4_49[11],stage4_48[16],stage4_47[17]}
   );
   gpc615_5 gpc9979 (
      {stage3_47[46], stage3_47[47], stage3_47[48], stage3_47[49], stage3_47[50]},
      {stage3_48[34]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[9],stage4_49[12],stage4_48[17],stage4_47[18]}
   );
   gpc615_5 gpc9980 (
      {stage3_47[51], stage3_47[52], stage3_47[53], stage3_47[54], stage3_47[55]},
      {stage3_48[35]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[10],stage4_49[13],stage4_48[18],stage4_47[19]}
   );
   gpc615_5 gpc9981 (
      {stage3_47[56], stage3_47[57], stage3_47[58], stage3_47[59], stage3_47[60]},
      {stage3_48[36]},
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage4_51[6],stage4_50[11],stage4_49[14],stage4_48[19],stage4_47[20]}
   );
   gpc615_5 gpc9982 (
      {stage3_47[61], stage3_47[62], stage3_47[63], stage3_47[64], stage3_47[65]},
      {1'b0},
      {stage3_49[42], stage3_49[43], stage3_49[44], stage3_49[45], stage3_49[46], stage3_49[47]},
      {stage4_51[7],stage4_50[12],stage4_49[15],stage4_48[20],stage4_47[21]}
   );
   gpc615_5 gpc9983 (
      {stage3_47[66], stage3_47[67], stage3_47[68], stage3_47[69], stage3_47[70]},
      {1'b0},
      {stage3_49[48], stage3_49[49], stage3_49[50], stage3_49[51], stage3_49[52], stage3_49[53]},
      {stage4_51[8],stage4_50[13],stage4_49[16],stage4_48[21],stage4_47[22]}
   );
   gpc117_4 gpc9984 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[0]},
      {stage3_52[0]},
      {stage4_53[0],stage4_52[0],stage4_51[9],stage4_50[14]}
   );
   gpc117_4 gpc9985 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[1]},
      {stage3_52[1]},
      {stage4_53[1],stage4_52[1],stage4_51[10],stage4_50[15]}
   );
   gpc117_4 gpc9986 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18], stage3_50[19], stage3_50[20]},
      {stage3_51[2]},
      {stage3_52[2]},
      {stage4_53[2],stage4_52[2],stage4_51[11],stage4_50[16]}
   );
   gpc117_4 gpc9987 (
      {stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27]},
      {stage3_51[3]},
      {stage3_52[3]},
      {stage4_53[3],stage4_52[3],stage4_51[12],stage4_50[17]}
   );
   gpc117_4 gpc9988 (
      {stage3_50[28], stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33], stage3_50[34]},
      {stage3_51[4]},
      {stage3_52[4]},
      {stage4_53[4],stage4_52[4],stage4_51[13],stage4_50[18]}
   );
   gpc117_4 gpc9989 (
      {stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38], stage3_50[39], stage3_50[40], stage3_50[41]},
      {stage3_51[5]},
      {stage3_52[5]},
      {stage4_53[5],stage4_52[5],stage4_51[14],stage4_50[19]}
   );
   gpc117_4 gpc9990 (
      {stage3_50[42], stage3_50[43], stage3_50[44], stage3_50[45], stage3_50[46], stage3_50[47], stage3_50[48]},
      {stage3_51[6]},
      {stage3_52[6]},
      {stage4_53[6],stage4_52[6],stage4_51[15],stage4_50[20]}
   );
   gpc117_4 gpc9991 (
      {stage3_50[49], stage3_50[50], stage3_50[51], stage3_50[52], stage3_50[53], stage3_50[54], stage3_50[55]},
      {stage3_51[7]},
      {stage3_52[7]},
      {stage4_53[7],stage4_52[7],stage4_51[16],stage4_50[21]}
   );
   gpc117_4 gpc9992 (
      {stage3_50[56], stage3_50[57], stage3_50[58], stage3_50[59], stage3_50[60], stage3_50[61], stage3_50[62]},
      {stage3_51[8]},
      {stage3_52[8]},
      {stage4_53[8],stage4_52[8],stage4_51[17],stage4_50[22]}
   );
   gpc2135_5 gpc9993 (
      {stage3_51[9], stage3_51[10], stage3_51[11], stage3_51[12], stage3_51[13]},
      {stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[0],stage4_53[9],stage4_52[9],stage4_51[18]}
   );
   gpc2135_5 gpc9994 (
      {stage3_51[14], stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18]},
      {stage3_52[12], stage3_52[13], stage3_52[14]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[1],stage4_53[10],stage4_52[10],stage4_51[19]}
   );
   gpc2135_5 gpc9995 (
      {stage3_51[19], stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23]},
      {stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[2],stage4_53[11],stage4_52[11],stage4_51[20]}
   );
   gpc2135_5 gpc9996 (
      {stage3_51[24], stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28]},
      {stage3_52[18], stage3_52[19], stage3_52[20]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[3],stage4_53[12],stage4_52[12],stage4_51[21]}
   );
   gpc2135_5 gpc9997 (
      {stage3_51[29], stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33]},
      {stage3_52[21], stage3_52[22], stage3_52[23]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[4],stage4_53[13],stage4_52[13],stage4_51[22]}
   );
   gpc2135_5 gpc9998 (
      {stage3_51[34], stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38]},
      {stage3_52[24], stage3_52[25], stage3_52[26]},
      {stage3_53[5]},
      {stage3_54[10], stage3_54[11]},
      {stage4_55[5],stage4_54[5],stage4_53[14],stage4_52[14],stage4_51[23]}
   );
   gpc2135_5 gpc9999 (
      {stage3_51[39], stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43]},
      {stage3_52[27], stage3_52[28], stage3_52[29]},
      {stage3_53[6]},
      {stage3_54[12], stage3_54[13]},
      {stage4_55[6],stage4_54[6],stage4_53[15],stage4_52[15],stage4_51[24]}
   );
   gpc2135_5 gpc10000 (
      {stage3_51[44], stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48]},
      {stage3_52[30], stage3_52[31], stage3_52[32]},
      {stage3_53[7]},
      {stage3_54[14], stage3_54[15]},
      {stage4_55[7],stage4_54[7],stage4_53[16],stage4_52[16],stage4_51[25]}
   );
   gpc2135_5 gpc10001 (
      {stage3_51[49], stage3_51[50], stage3_51[51], stage3_51[52], stage3_51[53]},
      {stage3_52[33], stage3_52[34], stage3_52[35]},
      {stage3_53[8]},
      {stage3_54[16], stage3_54[17]},
      {stage4_55[8],stage4_54[8],stage4_53[17],stage4_52[17],stage4_51[26]}
   );
   gpc606_5 gpc10002 (
      {stage3_52[36], stage3_52[37], stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41]},
      {stage3_54[18], stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage4_56[0],stage4_55[9],stage4_54[9],stage4_53[18],stage4_52[18]}
   );
   gpc606_5 gpc10003 (
      {stage3_52[42], stage3_52[43], stage3_52[44], stage3_52[45], stage3_52[46], stage3_52[47]},
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28], stage3_54[29]},
      {stage4_56[1],stage4_55[10],stage4_54[10],stage4_53[19],stage4_52[19]}
   );
   gpc606_5 gpc10004 (
      {stage3_52[48], stage3_52[49], stage3_52[50], stage3_52[51], stage3_52[52], stage3_52[53]},
      {stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33], stage3_54[34], stage3_54[35]},
      {stage4_56[2],stage4_55[11],stage4_54[11],stage4_53[20],stage4_52[20]}
   );
   gpc1415_5 gpc10005 (
      {stage3_53[9], stage3_53[10], stage3_53[11], stage3_53[12], stage3_53[13]},
      {stage3_54[36]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[3],stage4_55[12],stage4_54[12],stage4_53[21]}
   );
   gpc1415_5 gpc10006 (
      {stage3_53[14], stage3_53[15], stage3_53[16], stage3_53[17], stage3_53[18]},
      {stage3_54[37]},
      {stage3_55[4], stage3_55[5], stage3_55[6], stage3_55[7]},
      {stage3_56[1]},
      {stage4_57[1],stage4_56[4],stage4_55[13],stage4_54[13],stage4_53[22]}
   );
   gpc1415_5 gpc10007 (
      {stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22], stage3_53[23]},
      {stage3_54[38]},
      {stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage3_56[2]},
      {stage4_57[2],stage4_56[5],stage4_55[14],stage4_54[14],stage4_53[23]}
   );
   gpc1415_5 gpc10008 (
      {stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_54[39]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15]},
      {stage3_56[3]},
      {stage4_57[3],stage4_56[6],stage4_55[15],stage4_54[15],stage4_53[24]}
   );
   gpc606_5 gpc10009 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[16], stage3_55[17], stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21]},
      {stage4_57[4],stage4_56[7],stage4_55[16],stage4_54[16],stage4_53[25]}
   );
   gpc606_5 gpc10010 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39], stage3_53[40]},
      {stage3_55[22], stage3_55[23], stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27]},
      {stage4_57[5],stage4_56[8],stage4_55[17],stage4_54[17],stage4_53[26]}
   );
   gpc606_5 gpc10011 (
      {stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44], stage3_53[45], stage3_53[46]},
      {stage3_55[28], stage3_55[29], stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33]},
      {stage4_57[6],stage4_56[9],stage4_55[18],stage4_54[18],stage4_53[27]}
   );
   gpc606_5 gpc10012 (
      {stage3_53[47], stage3_53[48], stage3_53[49], stage3_53[50], stage3_53[51], stage3_53[52]},
      {stage3_55[34], stage3_55[35], stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39]},
      {stage4_57[7],stage4_56[10],stage4_55[19],stage4_54[19],stage4_53[28]}
   );
   gpc207_4 gpc10013 (
      {stage3_54[40], stage3_54[41], stage3_54[42], stage3_54[43], stage3_54[44], stage3_54[45], stage3_54[46]},
      {stage3_56[4], stage3_56[5]},
      {stage4_57[8],stage4_56[11],stage4_55[20],stage4_54[20]}
   );
   gpc207_4 gpc10014 (
      {stage3_54[47], stage3_54[48], stage3_54[49], stage3_54[50], stage3_54[51], stage3_54[52], stage3_54[53]},
      {stage3_56[6], stage3_56[7]},
      {stage4_57[9],stage4_56[12],stage4_55[21],stage4_54[21]}
   );
   gpc606_5 gpc10015 (
      {stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12], stage3_56[13]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[0],stage4_58[0],stage4_57[10],stage4_56[13]}
   );
   gpc606_5 gpc10016 (
      {stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18], stage3_56[19]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[1],stage4_58[1],stage4_57[11],stage4_56[14]}
   );
   gpc606_5 gpc10017 (
      {stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23], stage3_56[24], stage3_56[25]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[2],stage4_58[2],stage4_57[12],stage4_56[15]}
   );
   gpc1163_5 gpc10018 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[3],stage4_59[3],stage4_58[3],stage4_57[13]}
   );
   gpc1163_5 gpc10019 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[4],stage4_59[4],stage4_58[4],stage4_57[14]}
   );
   gpc1163_5 gpc10020 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[5],stage4_59[5],stage4_58[5],stage4_57[15]}
   );
   gpc606_5 gpc10021 (
      {stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7], stage3_59[8]},
      {stage4_61[3],stage4_60[6],stage4_59[6],stage4_58[6],stage4_57[16]}
   );
   gpc606_5 gpc10022 (
      {stage3_57[15], stage3_57[16], stage3_57[17], stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[4],stage4_60[7],stage4_59[7],stage4_58[7],stage4_57[17]}
   );
   gpc606_5 gpc10023 (
      {stage3_57[21], stage3_57[22], stage3_57[23], stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[5],stage4_60[8],stage4_59[8],stage4_58[8],stage4_57[18]}
   );
   gpc606_5 gpc10024 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[6],stage4_60[9],stage4_59[9],stage4_58[9],stage4_57[19]}
   );
   gpc606_5 gpc10025 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[7],stage4_60[10],stage4_59[10],stage4_58[10],stage4_57[20]}
   );
   gpc606_5 gpc10026 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43], stage3_57[44]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[8],stage4_60[11],stage4_59[11],stage4_58[11],stage4_57[21]}
   );
   gpc606_5 gpc10027 (
      {stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48], stage3_57[49], stage3_57[50]},
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43], stage3_59[44]},
      {stage4_61[9],stage4_60[12],stage4_59[12],stage4_58[12],stage4_57[22]}
   );
   gpc1406_5 gpc10028 (
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_60[3], stage3_60[4], stage3_60[5], stage3_60[6]},
      {stage3_61[0]},
      {stage4_62[0],stage4_61[10],stage4_60[13],stage4_59[13],stage4_58[13]}
   );
   gpc606_5 gpc10029 (
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10], stage3_60[11], stage3_60[12]},
      {stage4_62[1],stage4_61[11],stage4_60[14],stage4_59[14],stage4_58[14]}
   );
   gpc1406_5 gpc10030 (
      {stage3_60[13], stage3_60[14], stage3_60[15], stage3_60[16], stage3_60[17], stage3_60[18]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0]},
      {stage4_64[0],stage4_63[0],stage4_62[2],stage4_61[12],stage4_60[15]}
   );
   gpc606_5 gpc10031 (
      {stage3_60[19], stage3_60[20], stage3_60[21], stage3_60[22], stage3_60[23], stage3_60[24]},
      {stage3_62[4], stage3_62[5], stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9]},
      {stage4_64[1],stage4_63[1],stage4_62[3],stage4_61[13],stage4_60[16]}
   );
   gpc606_5 gpc10032 (
      {stage3_60[25], stage3_60[26], stage3_60[27], stage3_60[28], stage3_60[29], stage3_60[30]},
      {stage3_62[10], stage3_62[11], stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15]},
      {stage4_64[2],stage4_63[2],stage4_62[4],stage4_61[14],stage4_60[17]}
   );
   gpc606_5 gpc10033 (
      {stage3_60[31], stage3_60[32], stage3_60[33], stage3_60[34], stage3_60[35], stage3_60[36]},
      {stage3_62[16], stage3_62[17], stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21]},
      {stage4_64[3],stage4_63[3],stage4_62[5],stage4_61[15],stage4_60[18]}
   );
   gpc606_5 gpc10034 (
      {stage3_60[37], stage3_60[38], stage3_60[39], stage3_60[40], stage3_60[41], stage3_60[42]},
      {stage3_62[22], stage3_62[23], stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27]},
      {stage4_64[4],stage4_63[4],stage4_62[6],stage4_61[16],stage4_60[19]}
   );
   gpc606_5 gpc10035 (
      {stage3_60[43], stage3_60[44], stage3_60[45], stage3_60[46], stage3_60[47], stage3_60[48]},
      {stage3_62[28], stage3_62[29], stage3_62[30], stage3_62[31], stage3_62[32], stage3_62[33]},
      {stage4_64[5],stage4_63[5],stage4_62[7],stage4_61[17],stage4_60[20]}
   );
   gpc606_5 gpc10036 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5], stage3_61[6]},
      {stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6]},
      {stage4_65[0],stage4_64[6],stage4_63[6],stage4_62[8],stage4_61[18]}
   );
   gpc606_5 gpc10037 (
      {stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11], stage3_61[12]},
      {stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11], stage3_63[12]},
      {stage4_65[1],stage4_64[7],stage4_63[7],stage4_62[9],stage4_61[19]}
   );
   gpc606_5 gpc10038 (
      {stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17], stage3_61[18]},
      {stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17], stage3_63[18]},
      {stage4_65[2],stage4_64[8],stage4_63[8],stage4_62[10],stage4_61[20]}
   );
   gpc606_5 gpc10039 (
      {stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23], stage3_61[24]},
      {stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23], stage3_63[24]},
      {stage4_65[3],stage4_64[9],stage4_63[9],stage4_62[11],stage4_61[21]}
   );
   gpc606_5 gpc10040 (
      {stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29], stage3_61[30]},
      {stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29], stage3_63[30]},
      {stage4_65[4],stage4_64[10],stage4_63[10],stage4_62[12],stage4_61[22]}
   );
   gpc606_5 gpc10041 (
      {stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35], stage3_61[36]},
      {stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35], stage3_63[36]},
      {stage4_65[5],stage4_64[11],stage4_63[11],stage4_62[13],stage4_61[23]}
   );
   gpc606_5 gpc10042 (
      {stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41], stage3_61[42]},
      {stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41], stage3_63[42]},
      {stage4_65[6],stage4_64[12],stage4_63[12],stage4_62[14],stage4_61[24]}
   );
   gpc606_5 gpc10043 (
      {stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47], stage3_61[48]},
      {stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47], stage3_63[48]},
      {stage4_65[7],stage4_64[13],stage4_63[13],stage4_62[15],stage4_61[25]}
   );
   gpc606_5 gpc10044 (
      {stage3_61[49], stage3_61[50], stage3_61[51], stage3_61[52], stage3_61[53], stage3_61[54]},
      {stage3_63[49], stage3_63[50], stage3_63[51], stage3_63[52], stage3_63[53], stage3_63[54]},
      {stage4_65[8],stage4_64[14],stage4_63[14],stage4_62[16],stage4_61[26]}
   );
   gpc606_5 gpc10045 (
      {stage3_63[55], stage3_63[56], stage3_63[57], stage3_63[58], stage3_63[59], stage3_63[60]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[9],stage4_64[15],stage4_63[15]}
   );
   gpc606_5 gpc10046 (
      {stage3_63[61], stage3_63[62], stage3_63[63], stage3_63[64], stage3_63[65], stage3_63[66]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[1],stage4_65[10],stage4_64[16],stage4_63[16]}
   );
   gpc606_5 gpc10047 (
      {stage3_63[67], stage3_63[68], stage3_63[69], stage3_63[70], stage3_63[71], 1'b0},
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage4_67[2],stage4_66[2],stage4_65[11],stage4_64[17],stage4_63[17]}
   );
   gpc1163_5 gpc10048 (
      {stage3_64[0], stage3_64[1], stage3_64[2]},
      {stage3_65[18], stage3_65[19], stage3_65[20], stage3_65[21], stage3_65[22], stage3_65[23]},
      {stage3_66[0]},
      {stage3_67[0]},
      {stage4_68[0],stage4_67[3],stage4_66[3],stage4_65[12],stage4_64[18]}
   );
   gpc606_5 gpc10049 (
      {stage3_64[3], stage3_64[4], stage3_64[5], stage3_64[6], stage3_64[7], stage3_64[8]},
      {stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5], stage3_66[6]},
      {stage4_68[1],stage4_67[4],stage4_66[4],stage4_65[13],stage4_64[19]}
   );
   gpc606_5 gpc10050 (
      {stage3_64[9], stage3_64[10], stage3_64[11], stage3_64[12], stage3_64[13], stage3_64[14]},
      {stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11], stage3_66[12]},
      {stage4_68[2],stage4_67[5],stage4_66[5],stage4_65[14],stage4_64[20]}
   );
   gpc606_5 gpc10051 (
      {stage3_64[15], stage3_64[16], stage3_64[17], stage3_64[18], stage3_64[19], stage3_64[20]},
      {stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17], stage3_66[18]},
      {stage4_68[3],stage4_67[6],stage4_66[6],stage4_65[15],stage4_64[21]}
   );
   gpc606_5 gpc10052 (
      {stage3_64[21], stage3_64[22], stage3_64[23], stage3_64[24], stage3_64[25], stage3_64[26]},
      {stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23], stage3_66[24]},
      {stage4_68[4],stage4_67[7],stage4_66[7],stage4_65[16],stage4_64[22]}
   );
   gpc606_5 gpc10053 (
      {stage3_64[27], stage3_64[28], stage3_64[29], stage3_64[30], stage3_64[31], stage3_64[32]},
      {stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29], stage3_66[30]},
      {stage4_68[5],stage4_67[8],stage4_66[8],stage4_65[17],stage4_64[23]}
   );
   gpc606_5 gpc10054 (
      {stage3_64[33], stage3_64[34], stage3_64[35], stage3_64[36], stage3_64[37], stage3_64[38]},
      {stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35], stage3_66[36]},
      {stage4_68[6],stage4_67[9],stage4_66[9],stage4_65[18],stage4_64[24]}
   );
   gpc606_5 gpc10055 (
      {stage3_64[39], stage3_64[40], stage3_64[41], stage3_64[42], stage3_64[43], stage3_64[44]},
      {stage3_66[37], stage3_66[38], stage3_66[39], stage3_66[40], stage3_66[41], stage3_66[42]},
      {stage4_68[7],stage4_67[10],stage4_66[10],stage4_65[19],stage4_64[25]}
   );
   gpc606_5 gpc10056 (
      {stage3_64[45], stage3_64[46], stage3_64[47], stage3_64[48], stage3_64[49], stage3_64[50]},
      {stage3_66[43], stage3_66[44], stage3_66[45], stage3_66[46], stage3_66[47], stage3_66[48]},
      {stage4_68[8],stage4_67[11],stage4_66[11],stage4_65[20],stage4_64[26]}
   );
   gpc606_5 gpc10057 (
      {stage3_65[24], stage3_65[25], stage3_65[26], stage3_65[27], stage3_65[28], stage3_65[29]},
      {stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5], stage3_67[6]},
      {stage4_69[0],stage4_68[9],stage4_67[12],stage4_66[12],stage4_65[21]}
   );
   gpc606_5 gpc10058 (
      {stage3_65[30], stage3_65[31], stage3_65[32], 1'b0, 1'b0, 1'b0},
      {stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11], stage3_67[12]},
      {stage4_69[1],stage4_68[10],stage4_67[13],stage4_66[13],stage4_65[22]}
   );
   gpc606_5 gpc10059 (
      {stage3_66[49], stage3_66[50], stage3_66[51], stage3_66[52], stage3_66[53], 1'b0},
      {stage3_68[0], stage3_68[1], stage3_68[2], stage3_68[3], stage3_68[4], 1'b0},
      {stage4_70[0],stage4_69[2],stage4_68[11],stage4_67[14],stage4_66[14]}
   );
   gpc1_1 gpc10060 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc10061 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc10062 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc10063 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc10064 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc10065 (
      {stage3_1[24]},
      {stage4_1[5]}
   );
   gpc1_1 gpc10066 (
      {stage3_1[25]},
      {stage4_1[6]}
   );
   gpc1_1 gpc10067 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc10068 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc10069 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc10070 (
      {stage3_3[39]},
      {stage4_3[9]}
   );
   gpc1_1 gpc10071 (
      {stage3_3[40]},
      {stage4_3[10]}
   );
   gpc1_1 gpc10072 (
      {stage3_3[41]},
      {stage4_3[11]}
   );
   gpc1_1 gpc10073 (
      {stage3_3[42]},
      {stage4_3[12]}
   );
   gpc1_1 gpc10074 (
      {stage3_3[43]},
      {stage4_3[13]}
   );
   gpc1_1 gpc10075 (
      {stage3_3[44]},
      {stage4_3[14]}
   );
   gpc1_1 gpc10076 (
      {stage3_3[45]},
      {stage4_3[15]}
   );
   gpc1_1 gpc10077 (
      {stage3_3[46]},
      {stage4_3[16]}
   );
   gpc1_1 gpc10078 (
      {stage3_3[47]},
      {stage4_3[17]}
   );
   gpc1_1 gpc10079 (
      {stage3_3[48]},
      {stage4_3[18]}
   );
   gpc1_1 gpc10080 (
      {stage3_3[49]},
      {stage4_3[19]}
   );
   gpc1_1 gpc10081 (
      {stage3_3[50]},
      {stage4_3[20]}
   );
   gpc1_1 gpc10082 (
      {stage3_3[51]},
      {stage4_3[21]}
   );
   gpc1_1 gpc10083 (
      {stage3_4[51]},
      {stage4_4[16]}
   );
   gpc1_1 gpc10084 (
      {stage3_4[52]},
      {stage4_4[17]}
   );
   gpc1_1 gpc10085 (
      {stage3_4[53]},
      {stage4_4[18]}
   );
   gpc1_1 gpc10086 (
      {stage3_4[54]},
      {stage4_4[19]}
   );
   gpc1_1 gpc10087 (
      {stage3_4[55]},
      {stage4_4[20]}
   );
   gpc1_1 gpc10088 (
      {stage3_4[56]},
      {stage4_4[21]}
   );
   gpc1_1 gpc10089 (
      {stage3_4[57]},
      {stage4_4[22]}
   );
   gpc1_1 gpc10090 (
      {stage3_4[58]},
      {stage4_4[23]}
   );
   gpc1_1 gpc10091 (
      {stage3_4[59]},
      {stage4_4[24]}
   );
   gpc1_1 gpc10092 (
      {stage3_5[24]},
      {stage4_5[16]}
   );
   gpc1_1 gpc10093 (
      {stage3_5[25]},
      {stage4_5[17]}
   );
   gpc1_1 gpc10094 (
      {stage3_5[26]},
      {stage4_5[18]}
   );
   gpc1_1 gpc10095 (
      {stage3_5[27]},
      {stage4_5[19]}
   );
   gpc1_1 gpc10096 (
      {stage3_5[28]},
      {stage4_5[20]}
   );
   gpc1_1 gpc10097 (
      {stage3_5[29]},
      {stage4_5[21]}
   );
   gpc1_1 gpc10098 (
      {stage3_5[30]},
      {stage4_5[22]}
   );
   gpc1_1 gpc10099 (
      {stage3_5[31]},
      {stage4_5[23]}
   );
   gpc1_1 gpc10100 (
      {stage3_5[32]},
      {stage4_5[24]}
   );
   gpc1_1 gpc10101 (
      {stage3_5[33]},
      {stage4_5[25]}
   );
   gpc1_1 gpc10102 (
      {stage3_5[34]},
      {stage4_5[26]}
   );
   gpc1_1 gpc10103 (
      {stage3_5[35]},
      {stage4_5[27]}
   );
   gpc1_1 gpc10104 (
      {stage3_5[36]},
      {stage4_5[28]}
   );
   gpc1_1 gpc10105 (
      {stage3_5[37]},
      {stage4_5[29]}
   );
   gpc1_1 gpc10106 (
      {stage3_5[38]},
      {stage4_5[30]}
   );
   gpc1_1 gpc10107 (
      {stage3_5[39]},
      {stage4_5[31]}
   );
   gpc1_1 gpc10108 (
      {stage3_5[40]},
      {stage4_5[32]}
   );
   gpc1_1 gpc10109 (
      {stage3_5[41]},
      {stage4_5[33]}
   );
   gpc1_1 gpc10110 (
      {stage3_5[42]},
      {stage4_5[34]}
   );
   gpc1_1 gpc10111 (
      {stage3_5[43]},
      {stage4_5[35]}
   );
   gpc1_1 gpc10112 (
      {stage3_5[44]},
      {stage4_5[36]}
   );
   gpc1_1 gpc10113 (
      {stage3_5[45]},
      {stage4_5[37]}
   );
   gpc1_1 gpc10114 (
      {stage3_5[46]},
      {stage4_5[38]}
   );
   gpc1_1 gpc10115 (
      {stage3_5[47]},
      {stage4_5[39]}
   );
   gpc1_1 gpc10116 (
      {stage3_5[48]},
      {stage4_5[40]}
   );
   gpc1_1 gpc10117 (
      {stage3_5[49]},
      {stage4_5[41]}
   );
   gpc1_1 gpc10118 (
      {stage3_5[50]},
      {stage4_5[42]}
   );
   gpc1_1 gpc10119 (
      {stage3_5[51]},
      {stage4_5[43]}
   );
   gpc1_1 gpc10120 (
      {stage3_5[52]},
      {stage4_5[44]}
   );
   gpc1_1 gpc10121 (
      {stage3_5[53]},
      {stage4_5[45]}
   );
   gpc1_1 gpc10122 (
      {stage3_5[54]},
      {stage4_5[46]}
   );
   gpc1_1 gpc10123 (
      {stage3_6[62]},
      {stage4_6[16]}
   );
   gpc1_1 gpc10124 (
      {stage3_6[63]},
      {stage4_6[17]}
   );
   gpc1_1 gpc10125 (
      {stage3_6[64]},
      {stage4_6[18]}
   );
   gpc1_1 gpc10126 (
      {stage3_6[65]},
      {stage4_6[19]}
   );
   gpc1_1 gpc10127 (
      {stage3_6[66]},
      {stage4_6[20]}
   );
   gpc1_1 gpc10128 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc10129 (
      {stage3_7[36]},
      {stage4_7[21]}
   );
   gpc1_1 gpc10130 (
      {stage3_7[37]},
      {stage4_7[22]}
   );
   gpc1_1 gpc10131 (
      {stage3_7[38]},
      {stage4_7[23]}
   );
   gpc1_1 gpc10132 (
      {stage3_7[39]},
      {stage4_7[24]}
   );
   gpc1_1 gpc10133 (
      {stage3_7[40]},
      {stage4_7[25]}
   );
   gpc1_1 gpc10134 (
      {stage3_7[41]},
      {stage4_7[26]}
   );
   gpc1_1 gpc10135 (
      {stage3_7[42]},
      {stage4_7[27]}
   );
   gpc1_1 gpc10136 (
      {stage3_7[43]},
      {stage4_7[28]}
   );
   gpc1_1 gpc10137 (
      {stage3_7[44]},
      {stage4_7[29]}
   );
   gpc1_1 gpc10138 (
      {stage3_7[45]},
      {stage4_7[30]}
   );
   gpc1_1 gpc10139 (
      {stage3_7[46]},
      {stage4_7[31]}
   );
   gpc1_1 gpc10140 (
      {stage3_7[47]},
      {stage4_7[32]}
   );
   gpc1_1 gpc10141 (
      {stage3_7[48]},
      {stage4_7[33]}
   );
   gpc1_1 gpc10142 (
      {stage3_7[49]},
      {stage4_7[34]}
   );
   gpc1_1 gpc10143 (
      {stage3_7[50]},
      {stage4_7[35]}
   );
   gpc1_1 gpc10144 (
      {stage3_7[51]},
      {stage4_7[36]}
   );
   gpc1_1 gpc10145 (
      {stage3_7[52]},
      {stage4_7[37]}
   );
   gpc1_1 gpc10146 (
      {stage3_7[53]},
      {stage4_7[38]}
   );
   gpc1_1 gpc10147 (
      {stage3_7[54]},
      {stage4_7[39]}
   );
   gpc1_1 gpc10148 (
      {stage3_8[29]},
      {stage4_8[17]}
   );
   gpc1_1 gpc10149 (
      {stage3_8[30]},
      {stage4_8[18]}
   );
   gpc1_1 gpc10150 (
      {stage3_8[31]},
      {stage4_8[19]}
   );
   gpc1_1 gpc10151 (
      {stage3_8[32]},
      {stage4_8[20]}
   );
   gpc1_1 gpc10152 (
      {stage3_8[33]},
      {stage4_8[21]}
   );
   gpc1_1 gpc10153 (
      {stage3_8[34]},
      {stage4_8[22]}
   );
   gpc1_1 gpc10154 (
      {stage3_8[35]},
      {stage4_8[23]}
   );
   gpc1_1 gpc10155 (
      {stage3_8[36]},
      {stage4_8[24]}
   );
   gpc1_1 gpc10156 (
      {stage3_8[37]},
      {stage4_8[25]}
   );
   gpc1_1 gpc10157 (
      {stage3_8[38]},
      {stage4_8[26]}
   );
   gpc1_1 gpc10158 (
      {stage3_8[39]},
      {stage4_8[27]}
   );
   gpc1_1 gpc10159 (
      {stage3_8[40]},
      {stage4_8[28]}
   );
   gpc1_1 gpc10160 (
      {stage3_8[41]},
      {stage4_8[29]}
   );
   gpc1_1 gpc10161 (
      {stage3_8[42]},
      {stage4_8[30]}
   );
   gpc1_1 gpc10162 (
      {stage3_8[43]},
      {stage4_8[31]}
   );
   gpc1_1 gpc10163 (
      {stage3_8[44]},
      {stage4_8[32]}
   );
   gpc1_1 gpc10164 (
      {stage3_8[45]},
      {stage4_8[33]}
   );
   gpc1_1 gpc10165 (
      {stage3_8[46]},
      {stage4_8[34]}
   );
   gpc1_1 gpc10166 (
      {stage3_10[65]},
      {stage4_10[26]}
   );
   gpc1_1 gpc10167 (
      {stage3_10[66]},
      {stage4_10[27]}
   );
   gpc1_1 gpc10168 (
      {stage3_10[67]},
      {stage4_10[28]}
   );
   gpc1_1 gpc10169 (
      {stage3_11[52]},
      {stage4_11[25]}
   );
   gpc1_1 gpc10170 (
      {stage3_11[53]},
      {stage4_11[26]}
   );
   gpc1_1 gpc10171 (
      {stage3_11[54]},
      {stage4_11[27]}
   );
   gpc1_1 gpc10172 (
      {stage3_11[55]},
      {stage4_11[28]}
   );
   gpc1_1 gpc10173 (
      {stage3_11[56]},
      {stage4_11[29]}
   );
   gpc1_1 gpc10174 (
      {stage3_11[57]},
      {stage4_11[30]}
   );
   gpc1_1 gpc10175 (
      {stage3_11[58]},
      {stage4_11[31]}
   );
   gpc1_1 gpc10176 (
      {stage3_11[59]},
      {stage4_11[32]}
   );
   gpc1_1 gpc10177 (
      {stage3_11[60]},
      {stage4_11[33]}
   );
   gpc1_1 gpc10178 (
      {stage3_13[43]},
      {stage4_13[24]}
   );
   gpc1_1 gpc10179 (
      {stage3_13[44]},
      {stage4_13[25]}
   );
   gpc1_1 gpc10180 (
      {stage3_13[45]},
      {stage4_13[26]}
   );
   gpc1_1 gpc10181 (
      {stage3_13[46]},
      {stage4_13[27]}
   );
   gpc1_1 gpc10182 (
      {stage3_14[31]},
      {stage4_14[26]}
   );
   gpc1_1 gpc10183 (
      {stage3_14[32]},
      {stage4_14[27]}
   );
   gpc1_1 gpc10184 (
      {stage3_14[33]},
      {stage4_14[28]}
   );
   gpc1_1 gpc10185 (
      {stage3_14[34]},
      {stage4_14[29]}
   );
   gpc1_1 gpc10186 (
      {stage3_15[45]},
      {stage4_15[17]}
   );
   gpc1_1 gpc10187 (
      {stage3_15[46]},
      {stage4_15[18]}
   );
   gpc1_1 gpc10188 (
      {stage3_15[47]},
      {stage4_15[19]}
   );
   gpc1_1 gpc10189 (
      {stage3_15[48]},
      {stage4_15[20]}
   );
   gpc1_1 gpc10190 (
      {stage3_15[49]},
      {stage4_15[21]}
   );
   gpc1_1 gpc10191 (
      {stage3_15[50]},
      {stage4_15[22]}
   );
   gpc1_1 gpc10192 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc10193 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc10194 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc10195 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc10196 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc10197 (
      {stage3_16[45]},
      {stage4_16[19]}
   );
   gpc1_1 gpc10198 (
      {stage3_16[46]},
      {stage4_16[20]}
   );
   gpc1_1 gpc10199 (
      {stage3_16[47]},
      {stage4_16[21]}
   );
   gpc1_1 gpc10200 (
      {stage3_16[48]},
      {stage4_16[22]}
   );
   gpc1_1 gpc10201 (
      {stage3_16[49]},
      {stage4_16[23]}
   );
   gpc1_1 gpc10202 (
      {stage3_16[50]},
      {stage4_16[24]}
   );
   gpc1_1 gpc10203 (
      {stage3_16[51]},
      {stage4_16[25]}
   );
   gpc1_1 gpc10204 (
      {stage3_16[52]},
      {stage4_16[26]}
   );
   gpc1_1 gpc10205 (
      {stage3_16[53]},
      {stage4_16[27]}
   );
   gpc1_1 gpc10206 (
      {stage3_16[54]},
      {stage4_16[28]}
   );
   gpc1_1 gpc10207 (
      {stage3_16[55]},
      {stage4_16[29]}
   );
   gpc1_1 gpc10208 (
      {stage3_16[56]},
      {stage4_16[30]}
   );
   gpc1_1 gpc10209 (
      {stage3_16[57]},
      {stage4_16[31]}
   );
   gpc1_1 gpc10210 (
      {stage3_16[58]},
      {stage4_16[32]}
   );
   gpc1_1 gpc10211 (
      {stage3_17[36]},
      {stage4_17[15]}
   );
   gpc1_1 gpc10212 (
      {stage3_17[37]},
      {stage4_17[16]}
   );
   gpc1_1 gpc10213 (
      {stage3_17[38]},
      {stage4_17[17]}
   );
   gpc1_1 gpc10214 (
      {stage3_17[39]},
      {stage4_17[18]}
   );
   gpc1_1 gpc10215 (
      {stage3_17[40]},
      {stage4_17[19]}
   );
   gpc1_1 gpc10216 (
      {stage3_17[41]},
      {stage4_17[20]}
   );
   gpc1_1 gpc10217 (
      {stage3_17[42]},
      {stage4_17[21]}
   );
   gpc1_1 gpc10218 (
      {stage3_17[43]},
      {stage4_17[22]}
   );
   gpc1_1 gpc10219 (
      {stage3_18[52]},
      {stage4_18[20]}
   );
   gpc1_1 gpc10220 (
      {stage3_18[53]},
      {stage4_18[21]}
   );
   gpc1_1 gpc10221 (
      {stage3_18[54]},
      {stage4_18[22]}
   );
   gpc1_1 gpc10222 (
      {stage3_18[55]},
      {stage4_18[23]}
   );
   gpc1_1 gpc10223 (
      {stage3_18[56]},
      {stage4_18[24]}
   );
   gpc1_1 gpc10224 (
      {stage3_18[57]},
      {stage4_18[25]}
   );
   gpc1_1 gpc10225 (
      {stage3_18[58]},
      {stage4_18[26]}
   );
   gpc1_1 gpc10226 (
      {stage3_18[59]},
      {stage4_18[27]}
   );
   gpc1_1 gpc10227 (
      {stage3_18[60]},
      {stage4_18[28]}
   );
   gpc1_1 gpc10228 (
      {stage3_18[61]},
      {stage4_18[29]}
   );
   gpc1_1 gpc10229 (
      {stage3_18[62]},
      {stage4_18[30]}
   );
   gpc1_1 gpc10230 (
      {stage3_18[63]},
      {stage4_18[31]}
   );
   gpc1_1 gpc10231 (
      {stage3_20[57]},
      {stage4_20[21]}
   );
   gpc1_1 gpc10232 (
      {stage3_21[61]},
      {stage4_21[25]}
   );
   gpc1_1 gpc10233 (
      {stage3_21[62]},
      {stage4_21[26]}
   );
   gpc1_1 gpc10234 (
      {stage3_24[29]},
      {stage4_24[18]}
   );
   gpc1_1 gpc10235 (
      {stage3_24[30]},
      {stage4_24[19]}
   );
   gpc1_1 gpc10236 (
      {stage3_24[31]},
      {stage4_24[20]}
   );
   gpc1_1 gpc10237 (
      {stage3_24[32]},
      {stage4_24[21]}
   );
   gpc1_1 gpc10238 (
      {stage3_24[33]},
      {stage4_24[22]}
   );
   gpc1_1 gpc10239 (
      {stage3_24[34]},
      {stage4_24[23]}
   );
   gpc1_1 gpc10240 (
      {stage3_25[48]},
      {stage4_25[16]}
   );
   gpc1_1 gpc10241 (
      {stage3_25[49]},
      {stage4_25[17]}
   );
   gpc1_1 gpc10242 (
      {stage3_25[50]},
      {stage4_25[18]}
   );
   gpc1_1 gpc10243 (
      {stage3_25[51]},
      {stage4_25[19]}
   );
   gpc1_1 gpc10244 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc10245 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc10246 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc10247 (
      {stage3_28[57]},
      {stage4_28[19]}
   );
   gpc1_1 gpc10248 (
      {stage3_28[58]},
      {stage4_28[20]}
   );
   gpc1_1 gpc10249 (
      {stage3_28[59]},
      {stage4_28[21]}
   );
   gpc1_1 gpc10250 (
      {stage3_28[60]},
      {stage4_28[22]}
   );
   gpc1_1 gpc10251 (
      {stage3_28[61]},
      {stage4_28[23]}
   );
   gpc1_1 gpc10252 (
      {stage3_28[62]},
      {stage4_28[24]}
   );
   gpc1_1 gpc10253 (
      {stage3_28[63]},
      {stage4_28[25]}
   );
   gpc1_1 gpc10254 (
      {stage3_28[64]},
      {stage4_28[26]}
   );
   gpc1_1 gpc10255 (
      {stage3_28[65]},
      {stage4_28[27]}
   );
   gpc1_1 gpc10256 (
      {stage3_28[66]},
      {stage4_28[28]}
   );
   gpc1_1 gpc10257 (
      {stage3_28[67]},
      {stage4_28[29]}
   );
   gpc1_1 gpc10258 (
      {stage3_28[68]},
      {stage4_28[30]}
   );
   gpc1_1 gpc10259 (
      {stage3_28[69]},
      {stage4_28[31]}
   );
   gpc1_1 gpc10260 (
      {stage3_30[36]},
      {stage4_30[23]}
   );
   gpc1_1 gpc10261 (
      {stage3_30[37]},
      {stage4_30[24]}
   );
   gpc1_1 gpc10262 (
      {stage3_30[38]},
      {stage4_30[25]}
   );
   gpc1_1 gpc10263 (
      {stage3_32[51]},
      {stage4_32[19]}
   );
   gpc1_1 gpc10264 (
      {stage3_32[52]},
      {stage4_32[20]}
   );
   gpc1_1 gpc10265 (
      {stage3_32[53]},
      {stage4_32[21]}
   );
   gpc1_1 gpc10266 (
      {stage3_32[54]},
      {stage4_32[22]}
   );
   gpc1_1 gpc10267 (
      {stage3_32[55]},
      {stage4_32[23]}
   );
   gpc1_1 gpc10268 (
      {stage3_33[53]},
      {stage4_33[24]}
   );
   gpc1_1 gpc10269 (
      {stage3_33[54]},
      {stage4_33[25]}
   );
   gpc1_1 gpc10270 (
      {stage3_33[55]},
      {stage4_33[26]}
   );
   gpc1_1 gpc10271 (
      {stage3_33[56]},
      {stage4_33[27]}
   );
   gpc1_1 gpc10272 (
      {stage3_33[57]},
      {stage4_33[28]}
   );
   gpc1_1 gpc10273 (
      {stage3_33[58]},
      {stage4_33[29]}
   );
   gpc1_1 gpc10274 (
      {stage3_33[59]},
      {stage4_33[30]}
   );
   gpc1_1 gpc10275 (
      {stage3_33[60]},
      {stage4_33[31]}
   );
   gpc1_1 gpc10276 (
      {stage3_33[61]},
      {stage4_33[32]}
   );
   gpc1_1 gpc10277 (
      {stage3_33[62]},
      {stage4_33[33]}
   );
   gpc1_1 gpc10278 (
      {stage3_34[32]},
      {stage4_34[17]}
   );
   gpc1_1 gpc10279 (
      {stage3_34[33]},
      {stage4_34[18]}
   );
   gpc1_1 gpc10280 (
      {stage3_34[34]},
      {stage4_34[19]}
   );
   gpc1_1 gpc10281 (
      {stage3_34[35]},
      {stage4_34[20]}
   );
   gpc1_1 gpc10282 (
      {stage3_34[36]},
      {stage4_34[21]}
   );
   gpc1_1 gpc10283 (
      {stage3_34[37]},
      {stage4_34[22]}
   );
   gpc1_1 gpc10284 (
      {stage3_34[38]},
      {stage4_34[23]}
   );
   gpc1_1 gpc10285 (
      {stage3_34[39]},
      {stage4_34[24]}
   );
   gpc1_1 gpc10286 (
      {stage3_34[40]},
      {stage4_34[25]}
   );
   gpc1_1 gpc10287 (
      {stage3_34[41]},
      {stage4_34[26]}
   );
   gpc1_1 gpc10288 (
      {stage3_34[42]},
      {stage4_34[27]}
   );
   gpc1_1 gpc10289 (
      {stage3_34[43]},
      {stage4_34[28]}
   );
   gpc1_1 gpc10290 (
      {stage3_34[44]},
      {stage4_34[29]}
   );
   gpc1_1 gpc10291 (
      {stage3_35[52]},
      {stage4_35[19]}
   );
   gpc1_1 gpc10292 (
      {stage3_35[53]},
      {stage4_35[20]}
   );
   gpc1_1 gpc10293 (
      {stage3_35[54]},
      {stage4_35[21]}
   );
   gpc1_1 gpc10294 (
      {stage3_35[55]},
      {stage4_35[22]}
   );
   gpc1_1 gpc10295 (
      {stage3_35[56]},
      {stage4_35[23]}
   );
   gpc1_1 gpc10296 (
      {stage3_36[39]},
      {stage4_36[21]}
   );
   gpc1_1 gpc10297 (
      {stage3_36[40]},
      {stage4_36[22]}
   );
   gpc1_1 gpc10298 (
      {stage3_36[41]},
      {stage4_36[23]}
   );
   gpc1_1 gpc10299 (
      {stage3_36[42]},
      {stage4_36[24]}
   );
   gpc1_1 gpc10300 (
      {stage3_36[43]},
      {stage4_36[25]}
   );
   gpc1_1 gpc10301 (
      {stage3_36[44]},
      {stage4_36[26]}
   );
   gpc1_1 gpc10302 (
      {stage3_36[45]},
      {stage4_36[27]}
   );
   gpc1_1 gpc10303 (
      {stage3_36[46]},
      {stage4_36[28]}
   );
   gpc1_1 gpc10304 (
      {stage3_36[47]},
      {stage4_36[29]}
   );
   gpc1_1 gpc10305 (
      {stage3_36[48]},
      {stage4_36[30]}
   );
   gpc1_1 gpc10306 (
      {stage3_36[49]},
      {stage4_36[31]}
   );
   gpc1_1 gpc10307 (
      {stage3_36[50]},
      {stage4_36[32]}
   );
   gpc1_1 gpc10308 (
      {stage3_36[51]},
      {stage4_36[33]}
   );
   gpc1_1 gpc10309 (
      {stage3_36[52]},
      {stage4_36[34]}
   );
   gpc1_1 gpc10310 (
      {stage3_36[53]},
      {stage4_36[35]}
   );
   gpc1_1 gpc10311 (
      {stage3_36[54]},
      {stage4_36[36]}
   );
   gpc1_1 gpc10312 (
      {stage3_36[55]},
      {stage4_36[37]}
   );
   gpc1_1 gpc10313 (
      {stage3_38[60]},
      {stage4_38[18]}
   );
   gpc1_1 gpc10314 (
      {stage3_38[61]},
      {stage4_38[19]}
   );
   gpc1_1 gpc10315 (
      {stage3_38[62]},
      {stage4_38[20]}
   );
   gpc1_1 gpc10316 (
      {stage3_38[63]},
      {stage4_38[21]}
   );
   gpc1_1 gpc10317 (
      {stage3_38[64]},
      {stage4_38[22]}
   );
   gpc1_1 gpc10318 (
      {stage3_38[65]},
      {stage4_38[23]}
   );
   gpc1_1 gpc10319 (
      {stage3_38[66]},
      {stage4_38[24]}
   );
   gpc1_1 gpc10320 (
      {stage3_38[67]},
      {stage4_38[25]}
   );
   gpc1_1 gpc10321 (
      {stage3_38[68]},
      {stage4_38[26]}
   );
   gpc1_1 gpc10322 (
      {stage3_40[36]},
      {stage4_40[19]}
   );
   gpc1_1 gpc10323 (
      {stage3_40[37]},
      {stage4_40[20]}
   );
   gpc1_1 gpc10324 (
      {stage3_40[38]},
      {stage4_40[21]}
   );
   gpc1_1 gpc10325 (
      {stage3_40[39]},
      {stage4_40[22]}
   );
   gpc1_1 gpc10326 (
      {stage3_40[40]},
      {stage4_40[23]}
   );
   gpc1_1 gpc10327 (
      {stage3_40[41]},
      {stage4_40[24]}
   );
   gpc1_1 gpc10328 (
      {stage3_40[42]},
      {stage4_40[25]}
   );
   gpc1_1 gpc10329 (
      {stage3_40[43]},
      {stage4_40[26]}
   );
   gpc1_1 gpc10330 (
      {stage3_40[44]},
      {stage4_40[27]}
   );
   gpc1_1 gpc10331 (
      {stage3_40[45]},
      {stage4_40[28]}
   );
   gpc1_1 gpc10332 (
      {stage3_41[54]},
      {stage4_41[21]}
   );
   gpc1_1 gpc10333 (
      {stage3_41[55]},
      {stage4_41[22]}
   );
   gpc1_1 gpc10334 (
      {stage3_41[56]},
      {stage4_41[23]}
   );
   gpc1_1 gpc10335 (
      {stage3_43[55]},
      {stage4_43[18]}
   );
   gpc1_1 gpc10336 (
      {stage3_43[56]},
      {stage4_43[19]}
   );
   gpc1_1 gpc10337 (
      {stage3_43[57]},
      {stage4_43[20]}
   );
   gpc1_1 gpc10338 (
      {stage3_43[58]},
      {stage4_43[21]}
   );
   gpc1_1 gpc10339 (
      {stage3_43[59]},
      {stage4_43[22]}
   );
   gpc1_1 gpc10340 (
      {stage3_44[68]},
      {stage4_44[23]}
   );
   gpc1_1 gpc10341 (
      {stage3_44[69]},
      {stage4_44[24]}
   );
   gpc1_1 gpc10342 (
      {stage3_44[70]},
      {stage4_44[25]}
   );
   gpc1_1 gpc10343 (
      {stage3_44[71]},
      {stage4_44[26]}
   );
   gpc1_1 gpc10344 (
      {stage3_44[72]},
      {stage4_44[27]}
   );
   gpc1_1 gpc10345 (
      {stage3_44[73]},
      {stage4_44[28]}
   );
   gpc1_1 gpc10346 (
      {stage3_44[74]},
      {stage4_44[29]}
   );
   gpc1_1 gpc10347 (
      {stage3_44[75]},
      {stage4_44[30]}
   );
   gpc1_1 gpc10348 (
      {stage3_44[76]},
      {stage4_44[31]}
   );
   gpc1_1 gpc10349 (
      {stage3_44[77]},
      {stage4_44[32]}
   );
   gpc1_1 gpc10350 (
      {stage3_44[78]},
      {stage4_44[33]}
   );
   gpc1_1 gpc10351 (
      {stage3_44[79]},
      {stage4_44[34]}
   );
   gpc1_1 gpc10352 (
      {stage3_44[80]},
      {stage4_44[35]}
   );
   gpc1_1 gpc10353 (
      {stage3_44[81]},
      {stage4_44[36]}
   );
   gpc1_1 gpc10354 (
      {stage3_44[82]},
      {stage4_44[37]}
   );
   gpc1_1 gpc10355 (
      {stage3_44[83]},
      {stage4_44[38]}
   );
   gpc1_1 gpc10356 (
      {stage3_44[84]},
      {stage4_44[39]}
   );
   gpc1_1 gpc10357 (
      {stage3_46[46]},
      {stage4_46[22]}
   );
   gpc1_1 gpc10358 (
      {stage3_46[47]},
      {stage4_46[23]}
   );
   gpc1_1 gpc10359 (
      {stage3_46[48]},
      {stage4_46[24]}
   );
   gpc1_1 gpc10360 (
      {stage3_47[71]},
      {stage4_47[23]}
   );
   gpc1_1 gpc10361 (
      {stage3_47[72]},
      {stage4_47[24]}
   );
   gpc1_1 gpc10362 (
      {stage3_47[73]},
      {stage4_47[25]}
   );
   gpc1_1 gpc10363 (
      {stage3_49[54]},
      {stage4_49[17]}
   );
   gpc1_1 gpc10364 (
      {stage3_49[55]},
      {stage4_49[18]}
   );
   gpc1_1 gpc10365 (
      {stage3_49[56]},
      {stage4_49[19]}
   );
   gpc1_1 gpc10366 (
      {stage3_49[57]},
      {stage4_49[20]}
   );
   gpc1_1 gpc10367 (
      {stage3_49[58]},
      {stage4_49[21]}
   );
   gpc1_1 gpc10368 (
      {stage3_49[59]},
      {stage4_49[22]}
   );
   gpc1_1 gpc10369 (
      {stage3_49[60]},
      {stage4_49[23]}
   );
   gpc1_1 gpc10370 (
      {stage3_49[61]},
      {stage4_49[24]}
   );
   gpc1_1 gpc10371 (
      {stage3_49[62]},
      {stage4_49[25]}
   );
   gpc1_1 gpc10372 (
      {stage3_49[63]},
      {stage4_49[26]}
   );
   gpc1_1 gpc10373 (
      {stage3_49[64]},
      {stage4_49[27]}
   );
   gpc1_1 gpc10374 (
      {stage3_50[63]},
      {stage4_50[23]}
   );
   gpc1_1 gpc10375 (
      {stage3_52[54]},
      {stage4_52[21]}
   );
   gpc1_1 gpc10376 (
      {stage3_52[55]},
      {stage4_52[22]}
   );
   gpc1_1 gpc10377 (
      {stage3_54[54]},
      {stage4_54[22]}
   );
   gpc1_1 gpc10378 (
      {stage3_54[55]},
      {stage4_54[23]}
   );
   gpc1_1 gpc10379 (
      {stage3_54[56]},
      {stage4_54[24]}
   );
   gpc1_1 gpc10380 (
      {stage3_54[57]},
      {stage4_54[25]}
   );
   gpc1_1 gpc10381 (
      {stage3_54[58]},
      {stage4_54[26]}
   );
   gpc1_1 gpc10382 (
      {stage3_54[59]},
      {stage4_54[27]}
   );
   gpc1_1 gpc10383 (
      {stage3_54[60]},
      {stage4_54[28]}
   );
   gpc1_1 gpc10384 (
      {stage3_54[61]},
      {stage4_54[29]}
   );
   gpc1_1 gpc10385 (
      {stage3_54[62]},
      {stage4_54[30]}
   );
   gpc1_1 gpc10386 (
      {stage3_55[40]},
      {stage4_55[22]}
   );
   gpc1_1 gpc10387 (
      {stage3_55[41]},
      {stage4_55[23]}
   );
   gpc1_1 gpc10388 (
      {stage3_55[42]},
      {stage4_55[24]}
   );
   gpc1_1 gpc10389 (
      {stage3_55[43]},
      {stage4_55[25]}
   );
   gpc1_1 gpc10390 (
      {stage3_55[44]},
      {stage4_55[26]}
   );
   gpc1_1 gpc10391 (
      {stage3_55[45]},
      {stage4_55[27]}
   );
   gpc1_1 gpc10392 (
      {stage3_55[46]},
      {stage4_55[28]}
   );
   gpc1_1 gpc10393 (
      {stage3_56[26]},
      {stage4_56[16]}
   );
   gpc1_1 gpc10394 (
      {stage3_56[27]},
      {stage4_56[17]}
   );
   gpc1_1 gpc10395 (
      {stage3_56[28]},
      {stage4_56[18]}
   );
   gpc1_1 gpc10396 (
      {stage3_56[29]},
      {stage4_56[19]}
   );
   gpc1_1 gpc10397 (
      {stage3_56[30]},
      {stage4_56[20]}
   );
   gpc1_1 gpc10398 (
      {stage3_56[31]},
      {stage4_56[21]}
   );
   gpc1_1 gpc10399 (
      {stage3_56[32]},
      {stage4_56[22]}
   );
   gpc1_1 gpc10400 (
      {stage3_56[33]},
      {stage4_56[23]}
   );
   gpc1_1 gpc10401 (
      {stage3_56[34]},
      {stage4_56[24]}
   );
   gpc1_1 gpc10402 (
      {stage3_56[35]},
      {stage4_56[25]}
   );
   gpc1_1 gpc10403 (
      {stage3_56[36]},
      {stage4_56[26]}
   );
   gpc1_1 gpc10404 (
      {stage3_56[37]},
      {stage4_56[27]}
   );
   gpc1_1 gpc10405 (
      {stage3_56[38]},
      {stage4_56[28]}
   );
   gpc1_1 gpc10406 (
      {stage3_57[51]},
      {stage4_57[23]}
   );
   gpc1_1 gpc10407 (
      {stage3_57[52]},
      {stage4_57[24]}
   );
   gpc1_1 gpc10408 (
      {stage3_58[48]},
      {stage4_58[15]}
   );
   gpc1_1 gpc10409 (
      {stage3_59[45]},
      {stage4_59[15]}
   );
   gpc1_1 gpc10410 (
      {stage3_60[49]},
      {stage4_60[21]}
   );
   gpc1_1 gpc10411 (
      {stage3_60[50]},
      {stage4_60[22]}
   );
   gpc1_1 gpc10412 (
      {stage3_60[51]},
      {stage4_60[23]}
   );
   gpc1_1 gpc10413 (
      {stage3_60[52]},
      {stage4_60[24]}
   );
   gpc1_1 gpc10414 (
      {stage3_61[55]},
      {stage4_61[27]}
   );
   gpc1_1 gpc10415 (
      {stage3_61[56]},
      {stage4_61[28]}
   );
   gpc1_1 gpc10416 (
      {stage3_62[34]},
      {stage4_62[17]}
   );
   gpc1_1 gpc10417 (
      {stage3_62[35]},
      {stage4_62[18]}
   );
   gpc1_1 gpc10418 (
      {stage3_62[36]},
      {stage4_62[19]}
   );
   gpc1_1 gpc10419 (
      {stage3_62[37]},
      {stage4_62[20]}
   );
   gpc1_1 gpc10420 (
      {stage3_62[38]},
      {stage4_62[21]}
   );
   gpc1_1 gpc10421 (
      {stage3_62[39]},
      {stage4_62[22]}
   );
   gpc1_1 gpc10422 (
      {stage3_62[40]},
      {stage4_62[23]}
   );
   gpc1_1 gpc10423 (
      {stage3_67[13]},
      {stage4_67[15]}
   );
   gpc1_1 gpc10424 (
      {stage3_67[14]},
      {stage4_67[16]}
   );
   gpc606_5 gpc10425 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1406_5 gpc10426 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc1163_5 gpc10427 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[4]},
      {stage4_5[1]},
      {stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc606_5 gpc10428 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16], stage4_3[17]},
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage5_7[0],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc606_5 gpc10429 (
      {stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[1],stage5_6[3],stage5_5[4],stage5_4[4]}
   );
   gpc606_5 gpc10430 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[2],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc10431 (
      {stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21], stage4_4[22]},
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17]},
      {stage5_8[2],stage5_7[3],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc606_5 gpc10432 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc10433 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc10434 (
      {stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24], stage4_5[25]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[5],stage5_7[6],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc10435 (
      {stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage4_7[18], stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23]},
      {stage5_9[3],stage5_8[6],stage5_7[7],stage5_6[9],stage5_5[10]}
   );
   gpc606_5 gpc10436 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37]},
      {stage4_7[24], stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29]},
      {stage5_9[4],stage5_8[7],stage5_7[8],stage5_6[10],stage5_5[11]}
   );
   gpc615_5 gpc10437 (
      {stage4_7[30], stage4_7[31], stage4_7[32], stage4_7[33], stage4_7[34]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[5],stage5_8[8],stage5_7[9]}
   );
   gpc615_5 gpc10438 (
      {stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38], stage4_7[39]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[6],stage5_8[9],stage5_7[10]}
   );
   gpc1406_5 gpc10439 (
      {stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[7],stage5_8[10]}
   );
   gpc215_4 gpc10440 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage5_11[3],stage5_10[3],stage5_9[8],stage5_8[11]}
   );
   gpc215_4 gpc10441 (
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[13]},
      {stage4_10[6], stage4_10[7]},
      {stage5_11[4],stage5_10[4],stage5_9[9],stage5_8[12]}
   );
   gpc207_4 gpc10442 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24]},
      {stage4_10[8], stage4_10[9]},
      {stage5_11[5],stage5_10[5],stage5_9[10],stage5_8[13]}
   );
   gpc606_5 gpc10443 (
      {stage4_8[25], stage4_8[26], stage4_8[27], stage4_8[28], stage4_8[29], stage4_8[30]},
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15]},
      {stage5_12[1],stage5_11[6],stage5_10[6],stage5_9[11],stage5_8[14]}
   );
   gpc606_5 gpc10444 (
      {stage4_8[31], stage4_8[32], stage4_8[33], stage4_8[34], 1'b0, 1'b0},
      {stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19], stage4_10[20], stage4_10[21]},
      {stage5_12[2],stage5_11[7],stage5_10[7],stage5_9[12],stage5_8[15]}
   );
   gpc1163_5 gpc10445 (
      {stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[0]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[3],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc10446 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], 1'b0},
      {stage4_11[7]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[1],stage5_12[4],stage5_11[9],stage5_10[9]}
   );
   gpc615_5 gpc10447 (
      {stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12]},
      {stage4_12[7]},
      {stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[5],stage5_11[10]}
   );
   gpc615_5 gpc10448 (
      {stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage4_12[8]},
      {stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[6],stage5_11[11]}
   );
   gpc615_5 gpc10449 (
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22]},
      {stage4_12[9]},
      {stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[7],stage5_11[12]}
   );
   gpc615_5 gpc10450 (
      {stage4_11[23], stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27]},
      {stage4_12[10]},
      {stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[8],stage5_11[13]}
   );
   gpc615_5 gpc10451 (
      {stage4_12[11], stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15]},
      {stage4_13[25]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[9]}
   );
   gpc615_5 gpc10452 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc10453 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc10454 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc10455 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[10]}
   );
   gpc615_5 gpc10456 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc10457 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc10458 (
      {stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc606_5 gpc10459 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7],stage5_17[7]}
   );
   gpc2116_5 gpc10460 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[6]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc2116_5 gpc10461 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[1]},
      {stage4_21[2], stage4_21[3]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc2116_5 gpc10462 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[8]},
      {stage4_20[2]},
      {stage4_21[4], stage4_21[5]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc10463 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[9]},
      {stage4_20[3], stage4_20[4], stage4_20[5], stage4_20[6], stage4_20[7], stage4_20[8]},
      {stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[7],stage5_18[11]}
   );
   gpc615_5 gpc10464 (
      {stage4_18[23], stage4_18[24], stage4_18[25], stage4_18[26], stage4_18[27]},
      {stage4_19[10]},
      {stage4_20[9], stage4_20[10], stage4_20[11], stage4_20[12], stage4_20[13], stage4_20[14]},
      {stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[8],stage5_18[12]}
   );
   gpc615_5 gpc10465 (
      {stage4_18[28], stage4_18[29], stage4_18[30], stage4_18[31], 1'b0},
      {stage4_19[11]},
      {stage4_20[15], stage4_20[16], stage4_20[17], stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[9],stage5_18[13]}
   );
   gpc615_5 gpc10466 (
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16]},
      {stage4_20[21]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[0],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc7_3 gpc10467 (
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[1],stage5_22[7],stage5_21[8]}
   );
   gpc7_3 gpc10468 (
      {stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23], stage4_21[24], stage4_21[25]},
      {stage5_23[2],stage5_22[8],stage5_21[9]}
   );
   gpc1163_5 gpc10469 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[3],stage5_22[9]}
   );
   gpc1163_5 gpc10470 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage4_24[1]},
      {stage4_25[1]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[4],stage5_22[10]}
   );
   gpc1163_5 gpc10471 (
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[2]},
      {stage4_25[2]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[5],stage5_22[11]}
   );
   gpc615_5 gpc10472 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[18]},
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[6],stage5_22[12]}
   );
   gpc615_5 gpc10473 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[19]},
      {stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12], stage4_24[13], stage4_24[14]},
      {stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[7],stage5_22[13]}
   );
   gpc615_5 gpc10474 (
      {stage4_22[19], stage4_22[20], 1'b0, 1'b0, 1'b0},
      {stage4_23[20]},
      {stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18], stage4_24[19], stage4_24[20]},
      {stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[8],stage5_22[14]}
   );
   gpc606_5 gpc10475 (
      {stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[6],stage5_25[6]}
   );
   gpc606_5 gpc10476 (
      {stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12], stage4_25[13], stage4_25[14]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[7],stage5_25[7]}
   );
   gpc207_4 gpc10477 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[8]}
   );
   gpc207_4 gpc10478 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {stage4_28[2], stage4_28[3]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[9]}
   );
   gpc615_5 gpc10479 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_28[4]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4]}
   );
   gpc606_5 gpc10480 (
      {stage4_28[5], stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[5],stage5_28[5]}
   );
   gpc606_5 gpc10481 (
      {stage4_28[11], stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[6],stage5_28[6]}
   );
   gpc606_5 gpc10482 (
      {stage4_28[17], stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[3],stage5_30[3],stage5_29[7],stage5_28[7]}
   );
   gpc606_5 gpc10483 (
      {stage4_28[23], stage4_28[24], stage4_28[25], stage4_28[26], stage4_28[27], stage4_28[28]},
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23]},
      {stage5_32[3],stage5_31[4],stage5_30[4],stage5_29[8],stage5_28[8]}
   );
   gpc207_4 gpc10484 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[4],stage5_31[5],stage5_30[5],stage5_29[9]}
   );
   gpc207_4 gpc10485 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17], stage4_29[18], stage4_29[19]},
      {stage4_31[2], stage4_31[3]},
      {stage5_32[5],stage5_31[6],stage5_30[6],stage5_29[10]}
   );
   gpc615_5 gpc10486 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[0]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[6],stage5_31[7]}
   );
   gpc615_5 gpc10487 (
      {stage4_31[9], stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13]},
      {stage4_32[1]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[1],stage5_33[1],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc10488 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[2],stage5_34[2],stage5_33[2],stage5_32[8]}
   );
   gpc606_5 gpc10489 (
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage5_36[1],stage5_35[3],stage5_34[3],stage5_33[3],stage5_32[9]}
   );
   gpc606_5 gpc10490 (
      {stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17], stage4_32[18], stage4_32[19]},
      {stage4_34[12], stage4_34[13], stage4_34[14], stage4_34[15], stage4_34[16], stage4_34[17]},
      {stage5_36[2],stage5_35[4],stage5_34[4],stage5_33[4],stage5_32[10]}
   );
   gpc606_5 gpc10491 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[3],stage5_35[5],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc10492 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[4],stage5_35[6],stage5_34[6],stage5_33[6]}
   );
   gpc606_5 gpc10493 (
      {stage4_33[24], stage4_33[25], stage4_33[26], stage4_33[27], stage4_33[28], stage4_33[29]},
      {stage4_35[12], stage4_35[13], stage4_35[14], stage4_35[15], stage4_35[16], stage4_35[17]},
      {stage5_37[2],stage5_36[5],stage5_35[7],stage5_34[7],stage5_33[7]}
   );
   gpc606_5 gpc10494 (
      {stage4_33[30], stage4_33[31], stage4_33[32], stage4_33[33], 1'b0, 1'b0},
      {stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21], stage4_35[22], stage4_35[23]},
      {stage5_37[3],stage5_36[6],stage5_35[8],stage5_34[8],stage5_33[8]}
   );
   gpc1163_5 gpc10495 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[4],stage5_36[7]}
   );
   gpc1163_5 gpc10496 (
      {stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage4_38[1]},
      {stage4_39[1]},
      {stage5_40[1],stage5_39[1],stage5_38[1],stage5_37[5],stage5_36[8]}
   );
   gpc1163_5 gpc10497 (
      {stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], 1'b0, 1'b0},
      {stage4_38[2]},
      {stage4_39[2]},
      {stage5_40[2],stage5_39[2],stage5_38[2],stage5_37[6],stage5_36[9]}
   );
   gpc606_5 gpc10498 (
      {stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12], stage4_36[13], stage4_36[14]},
      {stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6], stage4_38[7], stage4_38[8]},
      {stage5_40[3],stage5_39[3],stage5_38[3],stage5_37[7],stage5_36[10]}
   );
   gpc606_5 gpc10499 (
      {stage4_36[15], stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20]},
      {stage4_38[9], stage4_38[10], stage4_38[11], stage4_38[12], stage4_38[13], stage4_38[14]},
      {stage5_40[4],stage5_39[4],stage5_38[4],stage5_37[8],stage5_36[11]}
   );
   gpc606_5 gpc10500 (
      {stage4_36[21], stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26]},
      {stage4_38[15], stage4_38[16], stage4_38[17], stage4_38[18], stage4_38[19], stage4_38[20]},
      {stage5_40[5],stage5_39[5],stage5_38[5],stage5_37[9],stage5_36[12]}
   );
   gpc606_5 gpc10501 (
      {stage4_36[27], stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32]},
      {stage4_38[21], stage4_38[22], stage4_38[23], stage4_38[24], stage4_38[25], stage4_38[26]},
      {stage5_40[6],stage5_39[6],stage5_38[6],stage5_37[10],stage5_36[13]}
   );
   gpc135_4 gpc10502 (
      {stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6], stage4_39[7]},
      {stage4_40[0], stage4_40[1], stage4_40[2]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[7],stage5_39[7]}
   );
   gpc135_4 gpc10503 (
      {stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12]},
      {stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[8],stage5_39[8]}
   );
   gpc135_4 gpc10504 (
      {stage4_39[13], stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17]},
      {stage4_40[6], stage4_40[7], stage4_40[8]},
      {stage4_41[2]},
      {stage5_42[2],stage5_41[2],stage5_40[9],stage5_39[9]}
   );
   gpc615_5 gpc10505 (
      {stage4_39[18], stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22]},
      {stage4_40[9]},
      {stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7], stage4_41[8]},
      {stage5_43[0],stage5_42[3],stage5_41[3],stage5_40[10],stage5_39[10]}
   );
   gpc606_5 gpc10506 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[4],stage5_41[4],stage5_40[11]}
   );
   gpc606_5 gpc10507 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[2],stage5_42[5],stage5_41[5],stage5_40[12]}
   );
   gpc606_5 gpc10508 (
      {stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13], stage4_41[14]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[3],stage5_42[6],stage5_41[6]}
   );
   gpc606_5 gpc10509 (
      {stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19], stage4_41[20]},
      {stage4_43[6], stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage5_45[1],stage5_44[3],stage5_43[4],stage5_42[7],stage5_41[7]}
   );
   gpc606_5 gpc10510 (
      {stage4_41[21], stage4_41[22], stage4_41[23], 1'b0, 1'b0, 1'b0},
      {stage4_43[12], stage4_43[13], stage4_43[14], stage4_43[15], stage4_43[16], stage4_43[17]},
      {stage5_45[2],stage5_44[4],stage5_43[5],stage5_42[8],stage5_41[8]}
   );
   gpc7_3 gpc10511 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17], stage4_42[18]},
      {stage5_44[5],stage5_43[6],stage5_42[9]}
   );
   gpc615_5 gpc10512 (
      {stage4_43[18], stage4_43[19], stage4_43[20], stage4_43[21], stage4_43[22]},
      {stage4_44[0]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[3],stage5_44[6],stage5_43[7]}
   );
   gpc135_4 gpc10513 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[1],stage5_45[4],stage5_44[7]}
   );
   gpc135_4 gpc10514 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[2],stage5_45[5],stage5_44[8]}
   );
   gpc135_4 gpc10515 (
      {stage4_44[11], stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[3],stage5_45[6],stage5_44[9]}
   );
   gpc135_4 gpc10516 (
      {stage4_44[16], stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20]},
      {stage4_45[15], stage4_45[16], stage4_45[17]},
      {stage4_46[3]},
      {stage5_47[4],stage5_46[4],stage5_45[7],stage5_44[10]}
   );
   gpc135_4 gpc10517 (
      {stage4_44[21], stage4_44[22], stage4_44[23], stage4_44[24], stage4_44[25]},
      {stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_46[4]},
      {stage5_47[5],stage5_46[5],stage5_45[8],stage5_44[11]}
   );
   gpc606_5 gpc10518 (
      {stage4_45[21], stage4_45[22], stage4_45[23], stage4_45[24], stage4_45[25], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[6],stage5_46[6],stage5_45[9]}
   );
   gpc2135_5 gpc10519 (
      {stage4_46[5], stage4_46[6], stage4_46[7], stage4_46[8], stage4_46[9]},
      {stage4_47[6], stage4_47[7], stage4_47[8]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[7],stage5_46[7]}
   );
   gpc2135_5 gpc10520 (
      {stage4_46[10], stage4_46[11], stage4_46[12], stage4_46[13], stage4_46[14]},
      {stage4_47[9], stage4_47[10], stage4_47[11]},
      {stage4_48[1]},
      {stage4_49[2], stage4_49[3]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[8],stage5_46[8]}
   );
   gpc2135_5 gpc10521 (
      {stage4_46[15], stage4_46[16], stage4_46[17], stage4_46[18], stage4_46[19]},
      {stage4_47[12], stage4_47[13], stage4_47[14]},
      {stage4_48[2]},
      {stage4_49[4], stage4_49[5]},
      {stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[9],stage5_46[9]}
   );
   gpc615_5 gpc10522 (
      {stage4_46[20], stage4_46[21], stage4_46[22], stage4_46[23], stage4_46[24]},
      {stage4_47[15]},
      {stage4_48[3], stage4_48[4], stage4_48[5], stage4_48[6], stage4_48[7], stage4_48[8]},
      {stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[10],stage5_46[10]}
   );
   gpc615_5 gpc10523 (
      {stage4_47[16], stage4_47[17], stage4_47[18], stage4_47[19], stage4_47[20]},
      {stage4_48[9]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[0],stage5_50[4],stage5_49[5],stage5_48[5],stage5_47[11]}
   );
   gpc615_5 gpc10524 (
      {stage4_47[21], stage4_47[22], stage4_47[23], stage4_47[24], stage4_47[25]},
      {stage4_48[10]},
      {stage4_49[12], stage4_49[13], stage4_49[14], stage4_49[15], stage4_49[16], stage4_49[17]},
      {stage5_51[1],stage5_50[5],stage5_49[6],stage5_48[6],stage5_47[12]}
   );
   gpc7_3 gpc10525 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[6]}
   );
   gpc7_3 gpc10526 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11], stage4_50[12], stage4_50[13]},
      {stage5_52[1],stage5_51[3],stage5_50[7]}
   );
   gpc615_5 gpc10527 (
      {stage4_50[14], stage4_50[15], stage4_50[16], stage4_50[17], stage4_50[18]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[2],stage5_51[4],stage5_50[8]}
   );
   gpc615_5 gpc10528 (
      {stage4_50[19], stage4_50[20], stage4_50[21], stage4_50[22], stage4_50[23]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[3],stage5_51[5],stage5_50[9]}
   );
   gpc117_4 gpc10529 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6], stage4_51[7], stage4_51[8]},
      {stage4_52[12]},
      {stage4_53[0]},
      {stage5_54[2],stage5_53[2],stage5_52[4],stage5_51[6]}
   );
   gpc606_5 gpc10530 (
      {stage4_51[9], stage4_51[10], stage4_51[11], stage4_51[12], stage4_51[13], stage4_51[14]},
      {stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5], stage4_53[6]},
      {stage5_55[0],stage5_54[3],stage5_53[3],stage5_52[5],stage5_51[7]}
   );
   gpc606_5 gpc10531 (
      {stage4_51[15], stage4_51[16], stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20]},
      {stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11], stage4_53[12]},
      {stage5_55[1],stage5_54[4],stage5_53[4],stage5_52[6],stage5_51[8]}
   );
   gpc606_5 gpc10532 (
      {stage4_51[21], stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17], stage4_53[18]},
      {stage5_55[2],stage5_54[5],stage5_53[5],stage5_52[7],stage5_51[9]}
   );
   gpc606_5 gpc10533 (
      {stage4_52[13], stage4_52[14], stage4_52[15], stage4_52[16], stage4_52[17], stage4_52[18]},
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5]},
      {stage5_56[0],stage5_55[3],stage5_54[6],stage5_53[6],stage5_52[8]}
   );
   gpc606_5 gpc10534 (
      {stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23], stage4_53[24]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[1],stage5_55[4],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc10535 (
      {stage4_54[6], stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10]},
      {stage4_55[6]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[1],stage5_56[2],stage5_55[5],stage5_54[8]}
   );
   gpc615_5 gpc10536 (
      {stage4_54[11], stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15]},
      {stage4_55[7]},
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage5_58[1],stage5_57[2],stage5_56[3],stage5_55[6],stage5_54[9]}
   );
   gpc615_5 gpc10537 (
      {stage4_54[16], stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20]},
      {stage4_55[8]},
      {stage4_56[12], stage4_56[13], stage4_56[14], stage4_56[15], stage4_56[16], stage4_56[17]},
      {stage5_58[2],stage5_57[3],stage5_56[4],stage5_55[7],stage5_54[10]}
   );
   gpc615_5 gpc10538 (
      {stage4_54[21], stage4_54[22], stage4_54[23], stage4_54[24], stage4_54[25]},
      {stage4_55[9]},
      {stage4_56[18], stage4_56[19], stage4_56[20], stage4_56[21], stage4_56[22], stage4_56[23]},
      {stage5_58[3],stage5_57[4],stage5_56[5],stage5_55[8],stage5_54[11]}
   );
   gpc606_5 gpc10539 (
      {stage4_55[10], stage4_55[11], stage4_55[12], stage4_55[13], stage4_55[14], stage4_55[15]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage5_59[0],stage5_58[4],stage5_57[5],stage5_56[6],stage5_55[9]}
   );
   gpc606_5 gpc10540 (
      {stage4_55[16], stage4_55[17], stage4_55[18], stage4_55[19], stage4_55[20], stage4_55[21]},
      {stage4_57[6], stage4_57[7], stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11]},
      {stage5_59[1],stage5_58[5],stage5_57[6],stage5_56[7],stage5_55[10]}
   );
   gpc207_4 gpc10541 (
      {stage4_57[12], stage4_57[13], stage4_57[14], stage4_57[15], stage4_57[16], stage4_57[17], stage4_57[18]},
      {stage4_59[0], stage4_59[1]},
      {stage5_60[0],stage5_59[2],stage5_58[6],stage5_57[7]}
   );
   gpc207_4 gpc10542 (
      {stage4_57[19], stage4_57[20], stage4_57[21], stage4_57[22], stage4_57[23], stage4_57[24], 1'b0},
      {stage4_59[2], stage4_59[3]},
      {stage5_60[1],stage5_59[3],stage5_58[7],stage5_57[8]}
   );
   gpc606_5 gpc10543 (
      {stage4_59[4], stage4_59[5], stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[2],stage5_59[4]}
   );
   gpc606_5 gpc10544 (
      {stage4_59[10], stage4_59[11], stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[3],stage5_59[5]}
   );
   gpc606_5 gpc10545 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[2],stage5_61[2],stage5_60[4]}
   );
   gpc606_5 gpc10546 (
      {stage4_60[6], stage4_60[7], stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11]},
      {stage4_62[6], stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage5_64[1],stage5_63[3],stage5_62[3],stage5_61[3],stage5_60[5]}
   );
   gpc606_5 gpc10547 (
      {stage4_60[12], stage4_60[13], stage4_60[14], stage4_60[15], stage4_60[16], stage4_60[17]},
      {stage4_62[12], stage4_62[13], stage4_62[14], stage4_62[15], stage4_62[16], stage4_62[17]},
      {stage5_64[2],stage5_63[4],stage5_62[4],stage5_61[4],stage5_60[6]}
   );
   gpc7_3 gpc10548 (
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17], stage4_61[18]},
      {stage5_63[5],stage5_62[5],stage5_61[5]}
   );
   gpc7_3 gpc10549 (
      {stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22], stage4_61[23], stage4_61[24], stage4_61[25]},
      {stage5_63[6],stage5_62[6],stage5_61[6]}
   );
   gpc606_5 gpc10550 (
      {stage4_62[18], stage4_62[19], stage4_62[20], stage4_62[21], stage4_62[22], stage4_62[23]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[0],stage5_64[3],stage5_63[7],stage5_62[7]}
   );
   gpc606_5 gpc10551 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[4],stage5_63[8]}
   );
   gpc606_5 gpc10552 (
      {stage4_63[6], stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8], stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[5],stage5_63[9]}
   );
   gpc606_5 gpc10553 (
      {stage4_63[12], stage4_63[13], stage4_63[14], stage4_63[15], stage4_63[16], stage4_63[17]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage5_67[2],stage5_66[3],stage5_65[3],stage5_64[6],stage5_63[10]}
   );
   gpc135_4 gpc10554 (
      {stage4_64[6], stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10]},
      {stage4_65[18], stage4_65[19], stage4_65[20]},
      {stage4_66[0]},
      {stage5_67[3],stage5_66[4],stage5_65[4],stage5_64[7]}
   );
   gpc135_4 gpc10555 (
      {stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15]},
      {stage4_65[21], stage4_65[22], 1'b0},
      {stage4_66[1]},
      {stage5_67[4],stage5_66[5],stage5_65[5],stage5_64[8]}
   );
   gpc1163_5 gpc10556 (
      {stage4_66[2], stage4_66[3], stage4_66[4]},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage4_68[0]},
      {stage4_69[0]},
      {stage5_70[0],stage5_69[0],stage5_68[0],stage5_67[5],stage5_66[6]}
   );
   gpc1163_5 gpc10557 (
      {stage4_66[5], stage4_66[6], stage4_66[7]},
      {stage4_67[6], stage4_67[7], stage4_67[8], stage4_67[9], stage4_67[10], stage4_67[11]},
      {stage4_68[1]},
      {stage4_69[1]},
      {stage5_70[1],stage5_69[1],stage5_68[1],stage5_67[6],stage5_66[7]}
   );
   gpc1163_5 gpc10558 (
      {stage4_66[8], stage4_66[9], stage4_66[10]},
      {stage4_67[12], stage4_67[13], stage4_67[14], stage4_67[15], stage4_67[16], 1'b0},
      {stage4_68[2]},
      {stage4_69[2]},
      {stage5_70[2],stage5_69[2],stage5_68[2],stage5_67[7],stage5_66[8]}
   );
   gpc1_1 gpc10559 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc10560 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc10561 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc10562 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc10563 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc10564 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc10565 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc10566 (
      {stage4_3[18]},
      {stage5_3[4]}
   );
   gpc1_1 gpc10567 (
      {stage4_3[19]},
      {stage5_3[5]}
   );
   gpc1_1 gpc10568 (
      {stage4_3[20]},
      {stage5_3[6]}
   );
   gpc1_1 gpc10569 (
      {stage4_3[21]},
      {stage5_3[7]}
   );
   gpc1_1 gpc10570 (
      {stage4_4[23]},
      {stage5_4[7]}
   );
   gpc1_1 gpc10571 (
      {stage4_4[24]},
      {stage5_4[8]}
   );
   gpc1_1 gpc10572 (
      {stage4_5[38]},
      {stage5_5[12]}
   );
   gpc1_1 gpc10573 (
      {stage4_5[39]},
      {stage5_5[13]}
   );
   gpc1_1 gpc10574 (
      {stage4_5[40]},
      {stage5_5[14]}
   );
   gpc1_1 gpc10575 (
      {stage4_5[41]},
      {stage5_5[15]}
   );
   gpc1_1 gpc10576 (
      {stage4_5[42]},
      {stage5_5[16]}
   );
   gpc1_1 gpc10577 (
      {stage4_5[43]},
      {stage5_5[17]}
   );
   gpc1_1 gpc10578 (
      {stage4_5[44]},
      {stage5_5[18]}
   );
   gpc1_1 gpc10579 (
      {stage4_5[45]},
      {stage5_5[19]}
   );
   gpc1_1 gpc10580 (
      {stage4_5[46]},
      {stage5_5[20]}
   );
   gpc1_1 gpc10581 (
      {stage4_6[18]},
      {stage5_6[11]}
   );
   gpc1_1 gpc10582 (
      {stage4_6[19]},
      {stage5_6[12]}
   );
   gpc1_1 gpc10583 (
      {stage4_6[20]},
      {stage5_6[13]}
   );
   gpc1_1 gpc10584 (
      {stage4_11[28]},
      {stage5_11[14]}
   );
   gpc1_1 gpc10585 (
      {stage4_11[29]},
      {stage5_11[15]}
   );
   gpc1_1 gpc10586 (
      {stage4_11[30]},
      {stage5_11[16]}
   );
   gpc1_1 gpc10587 (
      {stage4_11[31]},
      {stage5_11[17]}
   );
   gpc1_1 gpc10588 (
      {stage4_11[32]},
      {stage5_11[18]}
   );
   gpc1_1 gpc10589 (
      {stage4_11[33]},
      {stage5_11[19]}
   );
   gpc1_1 gpc10590 (
      {stage4_12[16]},
      {stage5_12[10]}
   );
   gpc1_1 gpc10591 (
      {stage4_12[17]},
      {stage5_12[11]}
   );
   gpc1_1 gpc10592 (
      {stage4_12[18]},
      {stage5_12[12]}
   );
   gpc1_1 gpc10593 (
      {stage4_12[19]},
      {stage5_12[13]}
   );
   gpc1_1 gpc10594 (
      {stage4_13[26]},
      {stage5_13[7]}
   );
   gpc1_1 gpc10595 (
      {stage4_13[27]},
      {stage5_13[8]}
   );
   gpc1_1 gpc10596 (
      {stage4_14[26]},
      {stage5_14[11]}
   );
   gpc1_1 gpc10597 (
      {stage4_14[27]},
      {stage5_14[12]}
   );
   gpc1_1 gpc10598 (
      {stage4_14[28]},
      {stage5_14[13]}
   );
   gpc1_1 gpc10599 (
      {stage4_14[29]},
      {stage5_14[14]}
   );
   gpc1_1 gpc10600 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc10601 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc10602 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc10603 (
      {stage4_15[22]},
      {stage5_15[15]}
   );
   gpc1_1 gpc10604 (
      {stage4_16[27]},
      {stage5_16[8]}
   );
   gpc1_1 gpc10605 (
      {stage4_16[28]},
      {stage5_16[9]}
   );
   gpc1_1 gpc10606 (
      {stage4_16[29]},
      {stage5_16[10]}
   );
   gpc1_1 gpc10607 (
      {stage4_16[30]},
      {stage5_16[11]}
   );
   gpc1_1 gpc10608 (
      {stage4_16[31]},
      {stage5_16[12]}
   );
   gpc1_1 gpc10609 (
      {stage4_16[32]},
      {stage5_16[13]}
   );
   gpc1_1 gpc10610 (
      {stage4_19[17]},
      {stage5_19[11]}
   );
   gpc1_1 gpc10611 (
      {stage4_19[18]},
      {stage5_19[12]}
   );
   gpc1_1 gpc10612 (
      {stage4_19[19]},
      {stage5_19[13]}
   );
   gpc1_1 gpc10613 (
      {stage4_21[26]},
      {stage5_21[10]}
   );
   gpc1_1 gpc10614 (
      {stage4_23[21]},
      {stage5_23[9]}
   );
   gpc1_1 gpc10615 (
      {stage4_23[22]},
      {stage5_23[10]}
   );
   gpc1_1 gpc10616 (
      {stage4_23[23]},
      {stage5_23[11]}
   );
   gpc1_1 gpc10617 (
      {stage4_24[21]},
      {stage5_24[6]}
   );
   gpc1_1 gpc10618 (
      {stage4_24[22]},
      {stage5_24[7]}
   );
   gpc1_1 gpc10619 (
      {stage4_24[23]},
      {stage5_24[8]}
   );
   gpc1_1 gpc10620 (
      {stage4_25[15]},
      {stage5_25[8]}
   );
   gpc1_1 gpc10621 (
      {stage4_25[16]},
      {stage5_25[9]}
   );
   gpc1_1 gpc10622 (
      {stage4_25[17]},
      {stage5_25[10]}
   );
   gpc1_1 gpc10623 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc10624 (
      {stage4_25[19]},
      {stage5_25[12]}
   );
   gpc1_1 gpc10625 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc10626 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc10627 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc10628 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc10629 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc10630 (
      {stage4_26[19]},
      {stage5_26[15]}
   );
   gpc1_1 gpc10631 (
      {stage4_26[20]},
      {stage5_26[16]}
   );
   gpc1_1 gpc10632 (
      {stage4_27[17]},
      {stage5_27[5]}
   );
   gpc1_1 gpc10633 (
      {stage4_27[18]},
      {stage5_27[6]}
   );
   gpc1_1 gpc10634 (
      {stage4_27[19]},
      {stage5_27[7]}
   );
   gpc1_1 gpc10635 (
      {stage4_27[20]},
      {stage5_27[8]}
   );
   gpc1_1 gpc10636 (
      {stage4_28[29]},
      {stage5_28[9]}
   );
   gpc1_1 gpc10637 (
      {stage4_28[30]},
      {stage5_28[10]}
   );
   gpc1_1 gpc10638 (
      {stage4_28[31]},
      {stage5_28[11]}
   );
   gpc1_1 gpc10639 (
      {stage4_29[20]},
      {stage5_29[11]}
   );
   gpc1_1 gpc10640 (
      {stage4_29[21]},
      {stage5_29[12]}
   );
   gpc1_1 gpc10641 (
      {stage4_29[22]},
      {stage5_29[13]}
   );
   gpc1_1 gpc10642 (
      {stage4_29[23]},
      {stage5_29[14]}
   );
   gpc1_1 gpc10643 (
      {stage4_30[24]},
      {stage5_30[7]}
   );
   gpc1_1 gpc10644 (
      {stage4_30[25]},
      {stage5_30[8]}
   );
   gpc1_1 gpc10645 (
      {stage4_31[14]},
      {stage5_31[9]}
   );
   gpc1_1 gpc10646 (
      {stage4_31[15]},
      {stage5_31[10]}
   );
   gpc1_1 gpc10647 (
      {stage4_31[16]},
      {stage5_31[11]}
   );
   gpc1_1 gpc10648 (
      {stage4_32[20]},
      {stage5_32[11]}
   );
   gpc1_1 gpc10649 (
      {stage4_32[21]},
      {stage5_32[12]}
   );
   gpc1_1 gpc10650 (
      {stage4_32[22]},
      {stage5_32[13]}
   );
   gpc1_1 gpc10651 (
      {stage4_32[23]},
      {stage5_32[14]}
   );
   gpc1_1 gpc10652 (
      {stage4_34[18]},
      {stage5_34[9]}
   );
   gpc1_1 gpc10653 (
      {stage4_34[19]},
      {stage5_34[10]}
   );
   gpc1_1 gpc10654 (
      {stage4_34[20]},
      {stage5_34[11]}
   );
   gpc1_1 gpc10655 (
      {stage4_34[21]},
      {stage5_34[12]}
   );
   gpc1_1 gpc10656 (
      {stage4_34[22]},
      {stage5_34[13]}
   );
   gpc1_1 gpc10657 (
      {stage4_34[23]},
      {stage5_34[14]}
   );
   gpc1_1 gpc10658 (
      {stage4_34[24]},
      {stage5_34[15]}
   );
   gpc1_1 gpc10659 (
      {stage4_34[25]},
      {stage5_34[16]}
   );
   gpc1_1 gpc10660 (
      {stage4_34[26]},
      {stage5_34[17]}
   );
   gpc1_1 gpc10661 (
      {stage4_34[27]},
      {stage5_34[18]}
   );
   gpc1_1 gpc10662 (
      {stage4_34[28]},
      {stage5_34[19]}
   );
   gpc1_1 gpc10663 (
      {stage4_34[29]},
      {stage5_34[20]}
   );
   gpc1_1 gpc10664 (
      {stage4_36[33]},
      {stage5_36[14]}
   );
   gpc1_1 gpc10665 (
      {stage4_36[34]},
      {stage5_36[15]}
   );
   gpc1_1 gpc10666 (
      {stage4_36[35]},
      {stage5_36[16]}
   );
   gpc1_1 gpc10667 (
      {stage4_36[36]},
      {stage5_36[17]}
   );
   gpc1_1 gpc10668 (
      {stage4_36[37]},
      {stage5_36[18]}
   );
   gpc1_1 gpc10669 (
      {stage4_40[22]},
      {stage5_40[13]}
   );
   gpc1_1 gpc10670 (
      {stage4_40[23]},
      {stage5_40[14]}
   );
   gpc1_1 gpc10671 (
      {stage4_40[24]},
      {stage5_40[15]}
   );
   gpc1_1 gpc10672 (
      {stage4_40[25]},
      {stage5_40[16]}
   );
   gpc1_1 gpc10673 (
      {stage4_40[26]},
      {stage5_40[17]}
   );
   gpc1_1 gpc10674 (
      {stage4_40[27]},
      {stage5_40[18]}
   );
   gpc1_1 gpc10675 (
      {stage4_40[28]},
      {stage5_40[19]}
   );
   gpc1_1 gpc10676 (
      {stage4_42[19]},
      {stage5_42[10]}
   );
   gpc1_1 gpc10677 (
      {stage4_42[20]},
      {stage5_42[11]}
   );
   gpc1_1 gpc10678 (
      {stage4_42[21]},
      {stage5_42[12]}
   );
   gpc1_1 gpc10679 (
      {stage4_42[22]},
      {stage5_42[13]}
   );
   gpc1_1 gpc10680 (
      {stage4_42[23]},
      {stage5_42[14]}
   );
   gpc1_1 gpc10681 (
      {stage4_42[24]},
      {stage5_42[15]}
   );
   gpc1_1 gpc10682 (
      {stage4_42[25]},
      {stage5_42[16]}
   );
   gpc1_1 gpc10683 (
      {stage4_42[26]},
      {stage5_42[17]}
   );
   gpc1_1 gpc10684 (
      {stage4_42[27]},
      {stage5_42[18]}
   );
   gpc1_1 gpc10685 (
      {stage4_42[28]},
      {stage5_42[19]}
   );
   gpc1_1 gpc10686 (
      {stage4_44[26]},
      {stage5_44[12]}
   );
   gpc1_1 gpc10687 (
      {stage4_44[27]},
      {stage5_44[13]}
   );
   gpc1_1 gpc10688 (
      {stage4_44[28]},
      {stage5_44[14]}
   );
   gpc1_1 gpc10689 (
      {stage4_44[29]},
      {stage5_44[15]}
   );
   gpc1_1 gpc10690 (
      {stage4_44[30]},
      {stage5_44[16]}
   );
   gpc1_1 gpc10691 (
      {stage4_44[31]},
      {stage5_44[17]}
   );
   gpc1_1 gpc10692 (
      {stage4_44[32]},
      {stage5_44[18]}
   );
   gpc1_1 gpc10693 (
      {stage4_44[33]},
      {stage5_44[19]}
   );
   gpc1_1 gpc10694 (
      {stage4_44[34]},
      {stage5_44[20]}
   );
   gpc1_1 gpc10695 (
      {stage4_44[35]},
      {stage5_44[21]}
   );
   gpc1_1 gpc10696 (
      {stage4_44[36]},
      {stage5_44[22]}
   );
   gpc1_1 gpc10697 (
      {stage4_44[37]},
      {stage5_44[23]}
   );
   gpc1_1 gpc10698 (
      {stage4_44[38]},
      {stage5_44[24]}
   );
   gpc1_1 gpc10699 (
      {stage4_44[39]},
      {stage5_44[25]}
   );
   gpc1_1 gpc10700 (
      {stage4_48[11]},
      {stage5_48[7]}
   );
   gpc1_1 gpc10701 (
      {stage4_48[12]},
      {stage5_48[8]}
   );
   gpc1_1 gpc10702 (
      {stage4_48[13]},
      {stage5_48[9]}
   );
   gpc1_1 gpc10703 (
      {stage4_48[14]},
      {stage5_48[10]}
   );
   gpc1_1 gpc10704 (
      {stage4_48[15]},
      {stage5_48[11]}
   );
   gpc1_1 gpc10705 (
      {stage4_48[16]},
      {stage5_48[12]}
   );
   gpc1_1 gpc10706 (
      {stage4_48[17]},
      {stage5_48[13]}
   );
   gpc1_1 gpc10707 (
      {stage4_48[18]},
      {stage5_48[14]}
   );
   gpc1_1 gpc10708 (
      {stage4_48[19]},
      {stage5_48[15]}
   );
   gpc1_1 gpc10709 (
      {stage4_48[20]},
      {stage5_48[16]}
   );
   gpc1_1 gpc10710 (
      {stage4_48[21]},
      {stage5_48[17]}
   );
   gpc1_1 gpc10711 (
      {stage4_49[18]},
      {stage5_49[7]}
   );
   gpc1_1 gpc10712 (
      {stage4_49[19]},
      {stage5_49[8]}
   );
   gpc1_1 gpc10713 (
      {stage4_49[20]},
      {stage5_49[9]}
   );
   gpc1_1 gpc10714 (
      {stage4_49[21]},
      {stage5_49[10]}
   );
   gpc1_1 gpc10715 (
      {stage4_49[22]},
      {stage5_49[11]}
   );
   gpc1_1 gpc10716 (
      {stage4_49[23]},
      {stage5_49[12]}
   );
   gpc1_1 gpc10717 (
      {stage4_49[24]},
      {stage5_49[13]}
   );
   gpc1_1 gpc10718 (
      {stage4_49[25]},
      {stage5_49[14]}
   );
   gpc1_1 gpc10719 (
      {stage4_49[26]},
      {stage5_49[15]}
   );
   gpc1_1 gpc10720 (
      {stage4_49[27]},
      {stage5_49[16]}
   );
   gpc1_1 gpc10721 (
      {stage4_52[19]},
      {stage5_52[9]}
   );
   gpc1_1 gpc10722 (
      {stage4_52[20]},
      {stage5_52[10]}
   );
   gpc1_1 gpc10723 (
      {stage4_52[21]},
      {stage5_52[11]}
   );
   gpc1_1 gpc10724 (
      {stage4_52[22]},
      {stage5_52[12]}
   );
   gpc1_1 gpc10725 (
      {stage4_53[25]},
      {stage5_53[8]}
   );
   gpc1_1 gpc10726 (
      {stage4_53[26]},
      {stage5_53[9]}
   );
   gpc1_1 gpc10727 (
      {stage4_53[27]},
      {stage5_53[10]}
   );
   gpc1_1 gpc10728 (
      {stage4_53[28]},
      {stage5_53[11]}
   );
   gpc1_1 gpc10729 (
      {stage4_54[26]},
      {stage5_54[12]}
   );
   gpc1_1 gpc10730 (
      {stage4_54[27]},
      {stage5_54[13]}
   );
   gpc1_1 gpc10731 (
      {stage4_54[28]},
      {stage5_54[14]}
   );
   gpc1_1 gpc10732 (
      {stage4_54[29]},
      {stage5_54[15]}
   );
   gpc1_1 gpc10733 (
      {stage4_54[30]},
      {stage5_54[16]}
   );
   gpc1_1 gpc10734 (
      {stage4_55[22]},
      {stage5_55[11]}
   );
   gpc1_1 gpc10735 (
      {stage4_55[23]},
      {stage5_55[12]}
   );
   gpc1_1 gpc10736 (
      {stage4_55[24]},
      {stage5_55[13]}
   );
   gpc1_1 gpc10737 (
      {stage4_55[25]},
      {stage5_55[14]}
   );
   gpc1_1 gpc10738 (
      {stage4_55[26]},
      {stage5_55[15]}
   );
   gpc1_1 gpc10739 (
      {stage4_55[27]},
      {stage5_55[16]}
   );
   gpc1_1 gpc10740 (
      {stage4_55[28]},
      {stage5_55[17]}
   );
   gpc1_1 gpc10741 (
      {stage4_56[24]},
      {stage5_56[8]}
   );
   gpc1_1 gpc10742 (
      {stage4_56[25]},
      {stage5_56[9]}
   );
   gpc1_1 gpc10743 (
      {stage4_56[26]},
      {stage5_56[10]}
   );
   gpc1_1 gpc10744 (
      {stage4_56[27]},
      {stage5_56[11]}
   );
   gpc1_1 gpc10745 (
      {stage4_56[28]},
      {stage5_56[12]}
   );
   gpc1_1 gpc10746 (
      {stage4_58[0]},
      {stage5_58[8]}
   );
   gpc1_1 gpc10747 (
      {stage4_58[1]},
      {stage5_58[9]}
   );
   gpc1_1 gpc10748 (
      {stage4_58[2]},
      {stage5_58[10]}
   );
   gpc1_1 gpc10749 (
      {stage4_58[3]},
      {stage5_58[11]}
   );
   gpc1_1 gpc10750 (
      {stage4_58[4]},
      {stage5_58[12]}
   );
   gpc1_1 gpc10751 (
      {stage4_58[5]},
      {stage5_58[13]}
   );
   gpc1_1 gpc10752 (
      {stage4_58[6]},
      {stage5_58[14]}
   );
   gpc1_1 gpc10753 (
      {stage4_58[7]},
      {stage5_58[15]}
   );
   gpc1_1 gpc10754 (
      {stage4_58[8]},
      {stage5_58[16]}
   );
   gpc1_1 gpc10755 (
      {stage4_58[9]},
      {stage5_58[17]}
   );
   gpc1_1 gpc10756 (
      {stage4_58[10]},
      {stage5_58[18]}
   );
   gpc1_1 gpc10757 (
      {stage4_58[11]},
      {stage5_58[19]}
   );
   gpc1_1 gpc10758 (
      {stage4_58[12]},
      {stage5_58[20]}
   );
   gpc1_1 gpc10759 (
      {stage4_58[13]},
      {stage5_58[21]}
   );
   gpc1_1 gpc10760 (
      {stage4_58[14]},
      {stage5_58[22]}
   );
   gpc1_1 gpc10761 (
      {stage4_58[15]},
      {stage5_58[23]}
   );
   gpc1_1 gpc10762 (
      {stage4_60[18]},
      {stage5_60[7]}
   );
   gpc1_1 gpc10763 (
      {stage4_60[19]},
      {stage5_60[8]}
   );
   gpc1_1 gpc10764 (
      {stage4_60[20]},
      {stage5_60[9]}
   );
   gpc1_1 gpc10765 (
      {stage4_60[21]},
      {stage5_60[10]}
   );
   gpc1_1 gpc10766 (
      {stage4_60[22]},
      {stage5_60[11]}
   );
   gpc1_1 gpc10767 (
      {stage4_60[23]},
      {stage5_60[12]}
   );
   gpc1_1 gpc10768 (
      {stage4_60[24]},
      {stage5_60[13]}
   );
   gpc1_1 gpc10769 (
      {stage4_61[26]},
      {stage5_61[7]}
   );
   gpc1_1 gpc10770 (
      {stage4_61[27]},
      {stage5_61[8]}
   );
   gpc1_1 gpc10771 (
      {stage4_61[28]},
      {stage5_61[9]}
   );
   gpc1_1 gpc10772 (
      {stage4_64[16]},
      {stage5_64[9]}
   );
   gpc1_1 gpc10773 (
      {stage4_64[17]},
      {stage5_64[10]}
   );
   gpc1_1 gpc10774 (
      {stage4_64[18]},
      {stage5_64[11]}
   );
   gpc1_1 gpc10775 (
      {stage4_64[19]},
      {stage5_64[12]}
   );
   gpc1_1 gpc10776 (
      {stage4_64[20]},
      {stage5_64[13]}
   );
   gpc1_1 gpc10777 (
      {stage4_64[21]},
      {stage5_64[14]}
   );
   gpc1_1 gpc10778 (
      {stage4_64[22]},
      {stage5_64[15]}
   );
   gpc1_1 gpc10779 (
      {stage4_64[23]},
      {stage5_64[16]}
   );
   gpc1_1 gpc10780 (
      {stage4_64[24]},
      {stage5_64[17]}
   );
   gpc1_1 gpc10781 (
      {stage4_64[25]},
      {stage5_64[18]}
   );
   gpc1_1 gpc10782 (
      {stage4_64[26]},
      {stage5_64[19]}
   );
   gpc1_1 gpc10783 (
      {stage4_66[11]},
      {stage5_66[9]}
   );
   gpc1_1 gpc10784 (
      {stage4_66[12]},
      {stage5_66[10]}
   );
   gpc1_1 gpc10785 (
      {stage4_66[13]},
      {stage5_66[11]}
   );
   gpc1_1 gpc10786 (
      {stage4_66[14]},
      {stage5_66[12]}
   );
   gpc1_1 gpc10787 (
      {stage4_68[3]},
      {stage5_68[3]}
   );
   gpc1_1 gpc10788 (
      {stage4_68[4]},
      {stage5_68[4]}
   );
   gpc1_1 gpc10789 (
      {stage4_68[5]},
      {stage5_68[5]}
   );
   gpc1_1 gpc10790 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc10791 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc10792 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc10793 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc10794 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc10795 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc10796 (
      {stage4_70[0]},
      {stage5_70[3]}
   );
   gpc615_5 gpc10797 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc207_4 gpc10798 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc10799 (
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc606_5 gpc10800 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], stage5_5[16], stage5_5[17]},
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10], 1'b0},
      {stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc117_4 gpc10801 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {1'b0},
      {stage5_8[0]},
      {stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[4]}
   );
   gpc615_5 gpc10802 (
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12], stage5_6[13]},
      {1'b0},
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[5],stage6_6[5]}
   );
   gpc606_5 gpc10803 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[4],stage6_8[4]}
   );
   gpc606_5 gpc10804 (
      {stage5_8[13], stage5_8[14], stage5_8[15], 1'b0, 1'b0, 1'b0},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], 1'b0, 1'b0},
      {stage6_12[1],stage6_11[1],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc207_4 gpc10805 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5], stage5_9[6]},
      {stage5_11[0], stage5_11[1]},
      {stage6_12[2],stage6_11[2],stage6_10[3],stage6_9[6]}
   );
   gpc606_5 gpc10806 (
      {stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11], stage5_9[12]},
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7]},
      {stage6_13[0],stage6_12[3],stage6_11[3],stage6_10[4],stage6_9[7]}
   );
   gpc1406_5 gpc10807 (
      {stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[4],stage6_11[4]}
   );
   gpc1406_5 gpc10808 (
      {stage5_11[14], stage5_11[15], stage5_11[16], stage5_11[17], stage5_11[18], stage5_11[19]},
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7]},
      {stage5_14[1]},
      {stage6_15[1],stage6_14[1],stage6_13[2],stage6_12[5],stage6_11[5]}
   );
   gpc117_4 gpc10809 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage5_13[8]},
      {stage5_14[2]},
      {stage6_15[2],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc117_4 gpc10810 (
      {stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {1'b0},
      {stage5_14[3]},
      {stage6_15[3],stage6_14[3],stage6_13[4],stage6_12[7]}
   );
   gpc1343_5 gpc10811 (
      {stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[4],stage6_14[4]}
   );
   gpc1343_5 gpc10812 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[5],stage6_14[5]}
   );
   gpc1343_5 gpc10813 (
      {stage5_14[10], stage5_14[11], stage5_14[12]},
      {stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage5_16[6], stage5_16[7], stage5_16[8]},
      {stage5_17[2]},
      {stage6_18[2],stage6_17[2],stage6_16[2],stage6_15[6],stage6_14[6]}
   );
   gpc1343_5 gpc10814 (
      {stage5_14[13], stage5_14[14], 1'b0},
      {stage5_15[12], stage5_15[13], stage5_15[14], stage5_15[15]},
      {stage5_16[9], stage5_16[10], stage5_16[11]},
      {stage5_17[3]},
      {stage6_18[3],stage6_17[3],stage6_16[3],stage6_15[7],stage6_14[7]}
   );
   gpc207_4 gpc10815 (
      {stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7], 1'b0, 1'b0, 1'b0},
      {stage5_19[0], stage5_19[1]},
      {stage6_20[0],stage6_19[0],stage6_18[4],stage6_17[4]}
   );
   gpc7_3 gpc10816 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage6_20[1],stage6_19[1],stage6_18[5]}
   );
   gpc7_3 gpc10817 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13]},
      {stage6_20[2],stage6_19[2],stage6_18[6]}
   );
   gpc2135_5 gpc10818 (
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[3],stage6_19[3]}
   );
   gpc7_3 gpc10819 (
      {stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13]},
      {stage6_21[1],stage6_20[4],stage6_19[4]}
   );
   gpc1415_5 gpc10820 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_21[1]},
      {stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[2],stage6_20[5]}
   );
   gpc207_4 gpc10821 (
      {stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5], stage5_21[6], stage5_21[7], stage5_21[8]},
      {stage5_23[1], stage5_23[2]},
      {stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[3]}
   );
   gpc606_5 gpc10822 (
      {stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[3]}
   );
   gpc606_5 gpc10823 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3]}
   );
   gpc1343_5 gpc10824 (
      {stage5_26[6], stage5_26[7], stage5_26[8]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[2],stage6_26[2]}
   );
   gpc1343_5 gpc10825 (
      {stage5_26[9], stage5_26[10], stage5_26[11]},
      {stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage5_29[1]},
      {stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc10826 (
      {stage5_26[12], stage5_26[13], stage5_26[14], stage5_26[15], stage5_26[16]},
      {stage5_27[8]},
      {stage5_28[6], stage5_28[7], stage5_28[8], stage5_28[9], stage5_28[10], stage5_28[11]},
      {stage6_30[2],stage6_29[2],stage6_28[3],stage6_27[4],stage6_26[4]}
   );
   gpc606_5 gpc10827 (
      {stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6], stage5_29[7]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[3],stage6_29[3]}
   );
   gpc606_5 gpc10828 (
      {stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11], stage5_29[12], stage5_29[13]},
      {stage5_31[6], stage5_31[7], stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11]},
      {stage6_33[1],stage6_32[1],stage6_31[1],stage6_30[4],stage6_29[4]}
   );
   gpc7_3 gpc10829 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage6_32[2],stage6_31[2],stage6_30[5]}
   );
   gpc1415_5 gpc10830 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4]},
      {stage5_33[0]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3]},
      {stage5_35[0]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[2],stage6_32[3]}
   );
   gpc1415_5 gpc10831 (
      {stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage5_33[1]},
      {stage5_34[4], stage5_34[5], stage5_34[6], stage5_34[7]},
      {stage5_35[1]},
      {stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[3],stage6_32[4]}
   );
   gpc606_5 gpc10832 (
      {stage5_32[10], stage5_32[11], stage5_32[12], stage5_32[13], stage5_32[14], 1'b0},
      {stage5_34[8], stage5_34[9], stage5_34[10], stage5_34[11], stage5_34[12], stage5_34[13]},
      {stage6_36[2],stage6_35[2],stage6_34[2],stage6_33[4],stage6_32[5]}
   );
   gpc615_5 gpc10833 (
      {stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_34[14]},
      {stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5], stage5_35[6], stage5_35[7]},
      {stage6_37[0],stage6_36[3],stage6_35[3],stage6_34[3],stage6_33[5]}
   );
   gpc615_5 gpc10834 (
      {stage5_34[15], stage5_34[16], stage5_34[17], stage5_34[18], stage5_34[19]},
      {stage5_35[8]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[4],stage6_35[4],stage6_34[4]}
   );
   gpc2135_5 gpc10835 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10]},
      {stage5_37[0], stage5_37[1], stage5_37[2]},
      {stage5_38[0]},
      {stage5_39[0], stage5_39[1]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[2],stage6_36[5]}
   );
   gpc2135_5 gpc10836 (
      {stage5_36[11], stage5_36[12], stage5_36[13], stage5_36[14], stage5_36[15]},
      {stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage5_38[1]},
      {stage5_39[2], stage5_39[3]},
      {stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[3],stage6_36[6]}
   );
   gpc606_5 gpc10837 (
      {stage5_36[16], stage5_36[17], stage5_36[18], 1'b0, 1'b0, 1'b0},
      {stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5], stage5_38[6], 1'b0},
      {stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[4],stage6_36[7]}
   );
   gpc606_5 gpc10838 (
      {stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10], 1'b0},
      {stage5_39[4], stage5_39[5], stage5_39[6], stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage6_41[0],stage6_40[3],stage6_39[3],stage6_38[4],stage6_37[5]}
   );
   gpc606_5 gpc10839 (
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[1],stage6_40[4]}
   );
   gpc606_5 gpc10840 (
      {stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9], stage5_40[10], stage5_40[11]},
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10], stage5_42[11]},
      {stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[2],stage6_40[5]}
   );
   gpc1325_5 gpc10841 (
      {stage5_40[12], stage5_40[13], stage5_40[14], stage5_40[15], stage5_40[16]},
      {stage5_41[0], stage5_41[1]},
      {stage5_42[12], stage5_42[13], stage5_42[14]},
      {stage5_43[0]},
      {stage6_44[2],stage6_43[2],stage6_42[2],stage6_41[3],stage6_40[6]}
   );
   gpc615_5 gpc10842 (
      {stage5_42[15], stage5_42[16], stage5_42[17], stage5_42[18], stage5_42[19]},
      {stage5_43[1]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[0],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc7_3 gpc10843 (
      {stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5], stage5_43[6], stage5_43[7], 1'b0},
      {stage6_45[1],stage6_44[4],stage6_43[4]}
   );
   gpc7_3 gpc10844 (
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11], stage5_44[12]},
      {stage6_46[1],stage6_45[2],stage6_44[5]}
   );
   gpc7_3 gpc10845 (
      {stage5_44[13], stage5_44[14], stage5_44[15], stage5_44[16], stage5_44[17], stage5_44[18], stage5_44[19]},
      {stage6_46[2],stage6_45[3],stage6_44[6]}
   );
   gpc606_5 gpc10846 (
      {stage5_44[20], stage5_44[21], stage5_44[22], stage5_44[23], stage5_44[24], stage5_44[25]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[3],stage6_45[4],stage6_44[7]}
   );
   gpc606_5 gpc10847 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc10848 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], 1'b0, 1'b0},
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10], stage5_47[11]},
      {stage6_49[1],stage6_48[2],stage6_47[2],stage6_46[5],stage6_45[6]}
   );
   gpc615_5 gpc10849 (
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10]},
      {stage5_47[12]},
      {stage5_48[0], stage5_48[1], stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5]},
      {stage6_50[0],stage6_49[2],stage6_48[3],stage6_47[3],stage6_46[6]}
   );
   gpc606_5 gpc10850 (
      {stage5_48[6], stage5_48[7], stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[1],stage6_49[3],stage6_48[4]}
   );
   gpc606_5 gpc10851 (
      {stage5_48[12], stage5_48[13], stage5_48[14], stage5_48[15], stage5_48[16], stage5_48[17]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], 1'b0, 1'b0},
      {stage6_52[1],stage6_51[1],stage6_50[2],stage6_49[4],stage6_48[5]}
   );
   gpc207_4 gpc10852 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5], stage5_49[6]},
      {stage5_51[0], stage5_51[1]},
      {stage6_52[2],stage6_51[2],stage6_50[3],stage6_49[5]}
   );
   gpc207_4 gpc10853 (
      {stage5_49[7], stage5_49[8], stage5_49[9], stage5_49[10], stage5_49[11], stage5_49[12], stage5_49[13]},
      {stage5_51[2], stage5_51[3]},
      {stage6_52[3],stage6_51[3],stage6_50[4],stage6_49[6]}
   );
   gpc606_5 gpc10854 (
      {stage5_51[4], stage5_51[5], stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[0],stage6_52[4],stage6_51[4]}
   );
   gpc606_5 gpc10855 (
      {stage5_52[0], stage5_52[1], stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5]},
      {stage5_54[0], stage5_54[1], stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5]},
      {stage6_56[0],stage6_55[1],stage6_54[1],stage6_53[1],stage6_52[5]}
   );
   gpc606_5 gpc10856 (
      {stage5_52[6], stage5_52[7], stage5_52[8], stage5_52[9], stage5_52[10], stage5_52[11]},
      {stage5_54[6], stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage6_56[1],stage6_55[2],stage6_54[2],stage6_53[2],stage6_52[6]}
   );
   gpc606_5 gpc10857 (
      {stage5_53[6], stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11]},
      {stage5_55[0], stage5_55[1], stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5]},
      {stage6_57[0],stage6_56[2],stage6_55[3],stage6_54[3],stage6_53[3]}
   );
   gpc1163_5 gpc10858 (
      {stage5_54[12], stage5_54[13], stage5_54[14]},
      {stage5_55[6], stage5_55[7], stage5_55[8], stage5_55[9], stage5_55[10], stage5_55[11]},
      {stage5_56[0]},
      {stage5_57[0]},
      {stage6_58[0],stage6_57[1],stage6_56[3],stage6_55[4],stage6_54[4]}
   );
   gpc1163_5 gpc10859 (
      {stage5_54[15], stage5_54[16], 1'b0},
      {stage5_55[12], stage5_55[13], stage5_55[14], stage5_55[15], stage5_55[16], stage5_55[17]},
      {stage5_56[1]},
      {stage5_57[1]},
      {stage6_58[1],stage6_57[2],stage6_56[4],stage6_55[5],stage6_54[5]}
   );
   gpc606_5 gpc10860 (
      {stage5_56[2], stage5_56[3], stage5_56[4], stage5_56[5], stage5_56[6], stage5_56[7]},
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage6_60[0],stage6_59[0],stage6_58[2],stage6_57[3],stage6_56[5]}
   );
   gpc606_5 gpc10861 (
      {stage5_56[8], stage5_56[9], stage5_56[10], stage5_56[11], stage5_56[12], 1'b0},
      {stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9], stage5_58[10], stage5_58[11]},
      {stage6_60[1],stage6_59[1],stage6_58[3],stage6_57[4],stage6_56[6]}
   );
   gpc606_5 gpc10862 (
      {stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5], stage5_57[6], stage5_57[7]},
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage6_61[0],stage6_60[2],stage6_59[2],stage6_58[4],stage6_57[5]}
   );
   gpc606_5 gpc10863 (
      {stage5_58[12], stage5_58[13], stage5_58[14], stage5_58[15], stage5_58[16], stage5_58[17]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[1],stage6_60[3],stage6_59[3],stage6_58[5]}
   );
   gpc606_5 gpc10864 (
      {stage5_58[18], stage5_58[19], stage5_58[20], stage5_58[21], stage5_58[22], stage5_58[23]},
      {stage5_60[6], stage5_60[7], stage5_60[8], stage5_60[9], stage5_60[10], stage5_60[11]},
      {stage6_62[1],stage6_61[2],stage6_60[4],stage6_59[4],stage6_58[6]}
   );
   gpc1343_5 gpc10865 (
      {stage5_61[0], stage5_61[1], stage5_61[2]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3]},
      {stage5_63[0], stage5_63[1], stage5_63[2]},
      {stage5_64[0]},
      {stage6_65[0],stage6_64[0],stage6_63[0],stage6_62[2],stage6_61[3]}
   );
   gpc1343_5 gpc10866 (
      {stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage5_62[4], stage5_62[5], stage5_62[6], stage5_62[7]},
      {stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage5_64[1]},
      {stage6_65[1],stage6_64[1],stage6_63[1],stage6_62[3],stage6_61[4]}
   );
   gpc606_5 gpc10867 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], 1'b0, 1'b0},
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], 1'b0},
      {stage6_65[2],stage6_64[2],stage6_63[2],stage6_62[4],stage6_61[5]}
   );
   gpc117_4 gpc10868 (
      {stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5], stage5_64[6], stage5_64[7], stage5_64[8]},
      {stage5_65[0]},
      {stage5_66[0]},
      {stage6_67[0],stage6_66[0],stage6_65[3],stage6_64[3]}
   );
   gpc606_5 gpc10869 (
      {stage5_64[9], stage5_64[10], stage5_64[11], stage5_64[12], stage5_64[13], stage5_64[14]},
      {stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], stage5_66[5], stage5_66[6]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[4],stage6_64[4]}
   );
   gpc615_5 gpc10870 (
      {stage5_64[15], stage5_64[16], stage5_64[17], stage5_64[18], stage5_64[19]},
      {stage5_65[1]},
      {stage5_66[7], stage5_66[8], stage5_66[9], stage5_66[10], stage5_66[11], stage5_66[12]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[5],stage6_64[5]}
   );
   gpc2135_5 gpc10871 (
      {stage5_67[0], stage5_67[1], stage5_67[2], stage5_67[3], stage5_67[4]},
      {stage5_68[0], stage5_68[1], stage5_68[2]},
      {stage5_69[0]},
      {stage5_70[0], stage5_70[1]},
      {stage6_71[0],stage6_70[0],stage6_69[0],stage6_68[2],stage6_67[3]}
   );
   gpc2135_5 gpc10872 (
      {stage5_67[5], stage5_67[6], stage5_67[7], 1'b0, 1'b0},
      {stage5_68[3], stage5_68[4], stage5_68[5]},
      {stage5_69[1]},
      {stage5_70[2], stage5_70[3]},
      {stage6_71[1],stage6_70[1],stage6_69[1],stage6_68[3],stage6_67[4]}
   );
   gpc1_1 gpc10873 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc10874 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc10875 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc10876 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc10877 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc10878 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc10879 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc10880 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc10881 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc10882 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc10883 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc10884 (
      {stage5_3[5]},
      {stage6_3[1]}
   );
   gpc1_1 gpc10885 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc10886 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc10887 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc10888 (
      {stage5_5[18]},
      {stage6_5[4]}
   );
   gpc1_1 gpc10889 (
      {stage5_5[19]},
      {stage6_5[5]}
   );
   gpc1_1 gpc10890 (
      {stage5_5[20]},
      {stage6_5[6]}
   );
   gpc1_1 gpc10891 (
      {stage5_16[12]},
      {stage6_16[4]}
   );
   gpc1_1 gpc10892 (
      {stage5_16[13]},
      {stage6_16[5]}
   );
   gpc1_1 gpc10893 (
      {stage5_21[9]},
      {stage6_21[4]}
   );
   gpc1_1 gpc10894 (
      {stage5_21[10]},
      {stage6_21[5]}
   );
   gpc1_1 gpc10895 (
      {stage5_22[6]},
      {stage6_22[3]}
   );
   gpc1_1 gpc10896 (
      {stage5_22[7]},
      {stage6_22[4]}
   );
   gpc1_1 gpc10897 (
      {stage5_22[8]},
      {stage6_22[5]}
   );
   gpc1_1 gpc10898 (
      {stage5_22[9]},
      {stage6_22[6]}
   );
   gpc1_1 gpc10899 (
      {stage5_22[10]},
      {stage6_22[7]}
   );
   gpc1_1 gpc10900 (
      {stage5_22[11]},
      {stage6_22[8]}
   );
   gpc1_1 gpc10901 (
      {stage5_22[12]},
      {stage6_22[9]}
   );
   gpc1_1 gpc10902 (
      {stage5_22[13]},
      {stage6_22[10]}
   );
   gpc1_1 gpc10903 (
      {stage5_22[14]},
      {stage6_22[11]}
   );
   gpc1_1 gpc10904 (
      {stage5_23[9]},
      {stage6_23[4]}
   );
   gpc1_1 gpc10905 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc10906 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc10907 (
      {stage5_24[6]},
      {stage6_24[4]}
   );
   gpc1_1 gpc10908 (
      {stage5_24[7]},
      {stage6_24[5]}
   );
   gpc1_1 gpc10909 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc10910 (
      {stage5_25[6]},
      {stage6_25[2]}
   );
   gpc1_1 gpc10911 (
      {stage5_25[7]},
      {stage6_25[3]}
   );
   gpc1_1 gpc10912 (
      {stage5_25[8]},
      {stage6_25[4]}
   );
   gpc1_1 gpc10913 (
      {stage5_25[9]},
      {stage6_25[5]}
   );
   gpc1_1 gpc10914 (
      {stage5_25[10]},
      {stage6_25[6]}
   );
   gpc1_1 gpc10915 (
      {stage5_25[11]},
      {stage6_25[7]}
   );
   gpc1_1 gpc10916 (
      {stage5_25[12]},
      {stage6_25[8]}
   );
   gpc1_1 gpc10917 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc10918 (
      {stage5_30[7]},
      {stage6_30[6]}
   );
   gpc1_1 gpc10919 (
      {stage5_30[8]},
      {stage6_30[7]}
   );
   gpc1_1 gpc10920 (
      {stage5_33[7]},
      {stage6_33[6]}
   );
   gpc1_1 gpc10921 (
      {stage5_33[8]},
      {stage6_33[7]}
   );
   gpc1_1 gpc10922 (
      {stage5_34[20]},
      {stage6_34[5]}
   );
   gpc1_1 gpc10923 (
      {stage5_39[10]},
      {stage6_39[4]}
   );
   gpc1_1 gpc10924 (
      {stage5_40[17]},
      {stage6_40[7]}
   );
   gpc1_1 gpc10925 (
      {stage5_40[18]},
      {stage6_40[8]}
   );
   gpc1_1 gpc10926 (
      {stage5_40[19]},
      {stage6_40[9]}
   );
   gpc1_1 gpc10927 (
      {stage5_41[2]},
      {stage6_41[4]}
   );
   gpc1_1 gpc10928 (
      {stage5_41[3]},
      {stage6_41[5]}
   );
   gpc1_1 gpc10929 (
      {stage5_41[4]},
      {stage6_41[6]}
   );
   gpc1_1 gpc10930 (
      {stage5_41[5]},
      {stage6_41[7]}
   );
   gpc1_1 gpc10931 (
      {stage5_41[6]},
      {stage6_41[8]}
   );
   gpc1_1 gpc10932 (
      {stage5_41[7]},
      {stage6_41[9]}
   );
   gpc1_1 gpc10933 (
      {stage5_41[8]},
      {stage6_41[10]}
   );
   gpc1_1 gpc10934 (
      {stage5_49[14]},
      {stage6_49[7]}
   );
   gpc1_1 gpc10935 (
      {stage5_49[15]},
      {stage6_49[8]}
   );
   gpc1_1 gpc10936 (
      {stage5_49[16]},
      {stage6_49[9]}
   );
   gpc1_1 gpc10937 (
      {stage5_52[12]},
      {stage6_52[7]}
   );
   gpc1_1 gpc10938 (
      {stage5_57[8]},
      {stage6_57[6]}
   );
   gpc1_1 gpc10939 (
      {stage5_60[12]},
      {stage6_60[5]}
   );
   gpc1_1 gpc10940 (
      {stage5_60[13]},
      {stage6_60[6]}
   );
   gpc1_1 gpc10941 (
      {stage5_65[2]},
      {stage6_65[6]}
   );
   gpc1_1 gpc10942 (
      {stage5_65[3]},
      {stage6_65[7]}
   );
   gpc1_1 gpc10943 (
      {stage5_65[4]},
      {stage6_65[8]}
   );
   gpc1_1 gpc10944 (
      {stage5_65[5]},
      {stage6_65[9]}
   );
   gpc1_1 gpc10945 (
      {stage5_68[6]},
      {stage6_68[4]}
   );
   gpc1_1 gpc10946 (
      {stage5_68[7]},
      {stage6_68[5]}
   );
   gpc1_1 gpc10947 (
      {stage5_68[8]},
      {stage6_68[6]}
   );
   gpc1_1 gpc10948 (
      {stage5_68[9]},
      {stage6_68[7]}
   );
   gpc1_1 gpc10949 (
      {stage5_68[10]},
      {stage6_68[8]}
   );
   gpc1_1 gpc10950 (
      {stage5_68[11]},
      {stage6_68[9]}
   );
   gpc1_1 gpc10951 (
      {stage5_69[2]},
      {stage6_69[2]}
   );
   gpc135_4 gpc10952 (
      {stage6_4[0], stage6_4[1], stage6_4[2], 1'b0, 1'b0},
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc615_5 gpc10953 (
      {stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_7[0]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1],stage7_6[1]}
   );
   gpc15_3 gpc10954 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc623_5 gpc10955 (
      {stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[2]}
   );
   gpc23_3 gpc10956 (
      {stage6_11[2], stage6_11[3], stage6_11[4]},
      {stage6_12[6], stage6_12[7]},
      {stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc117_4 gpc10957 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage6_15[0]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1]}
   );
   gpc7_3 gpc10958 (
      {stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5], stage6_15[6], stage6_15[7]},
      {stage7_17[1],stage7_16[1],stage7_15[1]}
   );
   gpc15_3 gpc10959 (
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4]},
      {stage6_18[0]},
      {stage7_19[0],stage7_18[0],stage7_17[2]}
   );
   gpc606_5 gpc10960 (
      {stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5], stage6_18[6]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[1],stage7_18[1]}
   );
   gpc1163_5 gpc10961 (
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_23[0]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1]}
   );
   gpc1163_5 gpc10962 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[6], stage6_22[7], stage6_22[8], stage6_22[9], stage6_22[10], stage6_22[11]},
      {stage6_23[1]},
      {stage6_24[1]},
      {stage7_25[1],stage7_24[1],stage7_23[1],stage7_22[2],stage7_21[2]}
   );
   gpc15_3 gpc10963 (
      {stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5], stage6_24[6]},
      {stage6_25[0]},
      {stage7_26[0],stage7_25[2],stage7_24[2]}
   );
   gpc606_5 gpc10964 (
      {stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5], stage6_25[6]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], 1'b0},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[3]}
   );
   gpc606_5 gpc10965 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], 1'b0, 1'b0},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[1]}
   );
   gpc1406_5 gpc10966 (
      {stage6_29[0], stage6_29[1], stage6_29[2], stage6_29[3], stage6_29[4], stage6_29[5]},
      {stage6_31[0], stage6_31[1], stage6_31[2], 1'b0},
      {stage6_32[0]},
      {stage7_33[0],stage7_32[1],stage7_31[1],stage7_30[1],stage7_29[2]}
   );
   gpc135_4 gpc10967 (
      {stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage6_33[0], stage6_33[1], stage6_33[2]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[1],stage7_32[2]}
   );
   gpc15_3 gpc10968 (
      {stage6_33[3], stage6_33[4], stage6_33[5], stage6_33[6], stage6_33[7]},
      {stage6_34[1]},
      {stage7_35[1],stage7_34[1],stage7_33[2]}
   );
   gpc117_4 gpc10969 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage6_37[0]},
      {stage6_38[0]},
      {stage7_39[0],stage7_38[0],stage7_37[0],stage7_36[0]}
   );
   gpc15_3 gpc10970 (
      {stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_38[1]},
      {stage7_39[1],stage7_38[1],stage7_37[1]}
   );
   gpc3_2 gpc10971 (
      {stage6_38[2], stage6_38[3], stage6_38[4]},
      {stage7_39[2],stage7_38[2]}
   );
   gpc2135_5 gpc10972 (
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], stage6_39[4]},
      {stage6_40[0], stage6_40[1], stage6_40[2]},
      {stage6_41[0]},
      {stage6_42[0], stage6_42[1]},
      {stage7_43[0],stage7_42[0],stage7_41[0],stage7_40[0],stage7_39[3]}
   );
   gpc207_4 gpc10973 (
      {stage6_40[3], stage6_40[4], stage6_40[5], stage6_40[6], stage6_40[7], stage6_40[8], stage6_40[9]},
      {stage6_42[2], stage6_42[3]},
      {stage7_43[1],stage7_42[1],stage7_41[1],stage7_40[1]}
   );
   gpc7_3 gpc10974 (
      {stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4], stage6_41[5], stage6_41[6], stage6_41[7]},
      {stage7_43[2],stage7_42[2],stage7_41[2]}
   );
   gpc215_4 gpc10975 (
      {stage6_43[0], stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4]},
      {stage6_44[0]},
      {stage6_45[0], stage6_45[1]},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[3]}
   );
   gpc207_4 gpc10976 (
      {stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], stage6_44[5], stage6_44[6], stage6_44[7]},
      {stage6_46[0], stage6_46[1]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1]}
   );
   gpc615_5 gpc10977 (
      {stage6_47[0], stage6_47[1], stage6_47[2], stage6_47[3], 1'b0},
      {stage6_48[0]},
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage7_51[0],stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1]}
   );
   gpc7_3 gpc10978 (
      {stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5], 1'b0, 1'b0},
      {stage7_50[1],stage7_49[1],stage7_48[1]}
   );
   gpc615_5 gpc10979 (
      {stage6_50[0], stage6_50[1], stage6_50[2], stage6_50[3], stage6_50[4]},
      {stage6_51[0]},
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4], stage6_52[5]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[2]}
   );
   gpc1343_5 gpc10980 (
      {stage6_52[6], stage6_52[7], 1'b0},
      {stage6_53[0], stage6_53[1], stage6_53[2], stage6_53[3]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc15_3 gpc10981 (
      {stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4], stage6_55[5]},
      {stage6_56[0]},
      {stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1423_5 gpc10982 (
      {stage6_56[1], stage6_56[2], stage6_56[3]},
      {stage6_57[0], stage6_57[1]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3]},
      {stage6_59[0]},
      {stage7_60[0],stage7_59[0],stage7_58[0],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc10983 (
      {stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5], stage6_57[6]},
      {stage6_58[4], stage6_58[5], stage6_58[6]},
      {stage6_59[1]},
      {stage7_60[1],stage7_59[1],stage7_58[1],stage7_57[2]}
   );
   gpc606_5 gpc10984 (
      {stage6_59[2], stage6_59[3], stage6_59[4], 1'b0, 1'b0, 1'b0},
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4], stage6_61[5]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[2],stage7_59[2]}
   );
   gpc606_5 gpc10985 (
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3], stage6_60[4], stage6_60[5]},
      {stage6_62[0], stage6_62[1], stage6_62[2], stage6_62[3], stage6_62[4], 1'b0},
      {stage7_64[0],stage7_63[1],stage7_62[1],stage7_61[1],stage7_60[3]}
   );
   gpc3_2 gpc10986 (
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage7_65[0],stage7_64[1]}
   );
   gpc3_2 gpc10987 (
      {stage6_64[3], stage6_64[4], stage6_64[5]},
      {stage7_65[1],stage7_64[2]}
   );
   gpc1163_5 gpc10988 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[0]}
   );
   gpc117_4 gpc10989 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc1_1 gpc10990 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc10991 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc10992 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc10993 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc10994 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc10995 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc10996 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc10997 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc10998 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc10999 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc11000 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc11001 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc11002 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc11003 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc11004 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc11005 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc11006 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc11007 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc11008 (
      {stage6_5[6]},
      {stage7_5[4]}
   );
   gpc1_1 gpc11009 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc11010 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc11011 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc11012 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc11013 (
      {stage6_7[5]},
      {stage7_7[6]}
   );
   gpc1_1 gpc11014 (
      {stage6_9[5]},
      {stage7_9[2]}
   );
   gpc1_1 gpc11015 (
      {stage6_9[6]},
      {stage7_9[3]}
   );
   gpc1_1 gpc11016 (
      {stage6_9[7]},
      {stage7_9[4]}
   );
   gpc1_1 gpc11017 (
      {stage6_10[4]},
      {stage7_10[3]}
   );
   gpc1_1 gpc11018 (
      {stage6_11[5]},
      {stage7_11[3]}
   );
   gpc1_1 gpc11019 (
      {stage6_13[0]},
      {stage7_13[2]}
   );
   gpc1_1 gpc11020 (
      {stage6_13[1]},
      {stage7_13[3]}
   );
   gpc1_1 gpc11021 (
      {stage6_13[2]},
      {stage7_13[4]}
   );
   gpc1_1 gpc11022 (
      {stage6_13[3]},
      {stage7_13[5]}
   );
   gpc1_1 gpc11023 (
      {stage6_13[4]},
      {stage7_13[6]}
   );
   gpc1_1 gpc11024 (
      {stage6_14[7]},
      {stage7_14[2]}
   );
   gpc1_1 gpc11025 (
      {stage6_16[1]},
      {stage7_16[2]}
   );
   gpc1_1 gpc11026 (
      {stage6_16[2]},
      {stage7_16[3]}
   );
   gpc1_1 gpc11027 (
      {stage6_16[3]},
      {stage7_16[4]}
   );
   gpc1_1 gpc11028 (
      {stage6_16[4]},
      {stage7_16[5]}
   );
   gpc1_1 gpc11029 (
      {stage6_16[5]},
      {stage7_16[6]}
   );
   gpc1_1 gpc11030 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc11031 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc11032 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc11033 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc11034 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc11035 (
      {stage6_23[2]},
      {stage7_23[2]}
   );
   gpc1_1 gpc11036 (
      {stage6_23[3]},
      {stage7_23[3]}
   );
   gpc1_1 gpc11037 (
      {stage6_23[4]},
      {stage7_23[4]}
   );
   gpc1_1 gpc11038 (
      {stage6_23[5]},
      {stage7_23[5]}
   );
   gpc1_1 gpc11039 (
      {stage6_23[6]},
      {stage7_23[6]}
   );
   gpc1_1 gpc11040 (
      {stage6_25[7]},
      {stage7_25[4]}
   );
   gpc1_1 gpc11041 (
      {stage6_25[8]},
      {stage7_25[5]}
   );
   gpc1_1 gpc11042 (
      {stage6_26[0]},
      {stage7_26[2]}
   );
   gpc1_1 gpc11043 (
      {stage6_26[1]},
      {stage7_26[3]}
   );
   gpc1_1 gpc11044 (
      {stage6_26[2]},
      {stage7_26[4]}
   );
   gpc1_1 gpc11045 (
      {stage6_26[3]},
      {stage7_26[5]}
   );
   gpc1_1 gpc11046 (
      {stage6_26[4]},
      {stage7_26[6]}
   );
   gpc1_1 gpc11047 (
      {stage6_30[6]},
      {stage7_30[2]}
   );
   gpc1_1 gpc11048 (
      {stage6_30[7]},
      {stage7_30[3]}
   );
   gpc1_1 gpc11049 (
      {stage6_34[2]},
      {stage7_34[2]}
   );
   gpc1_1 gpc11050 (
      {stage6_34[3]},
      {stage7_34[3]}
   );
   gpc1_1 gpc11051 (
      {stage6_34[4]},
      {stage7_34[4]}
   );
   gpc1_1 gpc11052 (
      {stage6_34[5]},
      {stage7_34[5]}
   );
   gpc1_1 gpc11053 (
      {stage6_35[0]},
      {stage7_35[2]}
   );
   gpc1_1 gpc11054 (
      {stage6_35[1]},
      {stage7_35[3]}
   );
   gpc1_1 gpc11055 (
      {stage6_35[2]},
      {stage7_35[4]}
   );
   gpc1_1 gpc11056 (
      {stage6_35[3]},
      {stage7_35[5]}
   );
   gpc1_1 gpc11057 (
      {stage6_35[4]},
      {stage7_35[6]}
   );
   gpc1_1 gpc11058 (
      {stage6_36[7]},
      {stage7_36[1]}
   );
   gpc1_1 gpc11059 (
      {stage6_41[8]},
      {stage7_41[3]}
   );
   gpc1_1 gpc11060 (
      {stage6_41[9]},
      {stage7_41[4]}
   );
   gpc1_1 gpc11061 (
      {stage6_41[10]},
      {stage7_41[5]}
   );
   gpc1_1 gpc11062 (
      {stage6_45[2]},
      {stage7_45[2]}
   );
   gpc1_1 gpc11063 (
      {stage6_45[3]},
      {stage7_45[3]}
   );
   gpc1_1 gpc11064 (
      {stage6_45[4]},
      {stage7_45[4]}
   );
   gpc1_1 gpc11065 (
      {stage6_45[5]},
      {stage7_45[5]}
   );
   gpc1_1 gpc11066 (
      {stage6_45[6]},
      {stage7_45[6]}
   );
   gpc1_1 gpc11067 (
      {stage6_46[2]},
      {stage7_46[2]}
   );
   gpc1_1 gpc11068 (
      {stage6_46[3]},
      {stage7_46[3]}
   );
   gpc1_1 gpc11069 (
      {stage6_46[4]},
      {stage7_46[4]}
   );
   gpc1_1 gpc11070 (
      {stage6_46[5]},
      {stage7_46[5]}
   );
   gpc1_1 gpc11071 (
      {stage6_46[6]},
      {stage7_46[6]}
   );
   gpc1_1 gpc11072 (
      {stage6_49[6]},
      {stage7_49[2]}
   );
   gpc1_1 gpc11073 (
      {stage6_49[7]},
      {stage7_49[3]}
   );
   gpc1_1 gpc11074 (
      {stage6_49[8]},
      {stage7_49[4]}
   );
   gpc1_1 gpc11075 (
      {stage6_49[9]},
      {stage7_49[5]}
   );
   gpc1_1 gpc11076 (
      {stage6_51[1]},
      {stage7_51[2]}
   );
   gpc1_1 gpc11077 (
      {stage6_51[2]},
      {stage7_51[3]}
   );
   gpc1_1 gpc11078 (
      {stage6_51[3]},
      {stage7_51[4]}
   );
   gpc1_1 gpc11079 (
      {stage6_51[4]},
      {stage7_51[5]}
   );
   gpc1_1 gpc11080 (
      {stage6_54[3]},
      {stage7_54[2]}
   );
   gpc1_1 gpc11081 (
      {stage6_54[4]},
      {stage7_54[3]}
   );
   gpc1_1 gpc11082 (
      {stage6_54[5]},
      {stage7_54[4]}
   );
   gpc1_1 gpc11083 (
      {stage6_56[4]},
      {stage7_56[3]}
   );
   gpc1_1 gpc11084 (
      {stage6_56[5]},
      {stage7_56[4]}
   );
   gpc1_1 gpc11085 (
      {stage6_56[6]},
      {stage7_56[5]}
   );
   gpc1_1 gpc11086 (
      {stage6_60[6]},
      {stage7_60[4]}
   );
   gpc1_1 gpc11087 (
      {stage6_63[0]},
      {stage7_63[2]}
   );
   gpc1_1 gpc11088 (
      {stage6_63[1]},
      {stage7_63[3]}
   );
   gpc1_1 gpc11089 (
      {stage6_63[2]},
      {stage7_63[4]}
   );
   gpc1_1 gpc11090 (
      {stage6_65[0]},
      {stage7_65[2]}
   );
   gpc1_1 gpc11091 (
      {stage6_65[1]},
      {stage7_65[3]}
   );
   gpc1_1 gpc11092 (
      {stage6_65[2]},
      {stage7_65[4]}
   );
   gpc1_1 gpc11093 (
      {stage6_65[3]},
      {stage7_65[5]}
   );
   gpc1_1 gpc11094 (
      {stage6_65[4]},
      {stage7_65[6]}
   );
   gpc1_1 gpc11095 (
      {stage6_65[5]},
      {stage7_65[7]}
   );
   gpc1_1 gpc11096 (
      {stage6_65[6]},
      {stage7_65[8]}
   );
   gpc1_1 gpc11097 (
      {stage6_65[7]},
      {stage7_65[9]}
   );
   gpc1_1 gpc11098 (
      {stage6_65[8]},
      {stage7_65[10]}
   );
   gpc1_1 gpc11099 (
      {stage6_65[9]},
      {stage7_65[11]}
   );
   gpc1_1 gpc11100 (
      {stage6_68[8]},
      {stage7_68[2]}
   );
   gpc1_1 gpc11101 (
      {stage6_68[9]},
      {stage7_68[3]}
   );
   gpc1_1 gpc11102 (
      {stage6_69[2]},
      {stage7_69[2]}
   );
   gpc1_1 gpc11103 (
      {stage6_70[1]},
      {stage7_70[2]}
   );
   gpc1_1 gpc11104 (
      {stage6_71[0]},
      {stage7_71[1]}
   );
   gpc1_1 gpc11105 (
      {stage6_71[1]},
      {stage7_71[2]}
   );
   gpc615_5 gpc11106 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], 1'b0, 1'b0, 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1415_5 gpc11107 (
      {stage7_3[0], stage7_3[1], stage7_3[2], stage7_3[3], 1'b0},
      {stage7_4[0]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc7_3 gpc11108 (
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5], stage7_7[6]},
      {stage8_9[0],stage8_8[0],stage8_7[1]}
   );
   gpc1415_5 gpc11109 (
      {stage7_9[0], stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4]},
      {stage7_10[0]},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc3_2 gpc11110 (
      {stage7_10[1], stage7_10[2], stage7_10[3]},
      {stage8_11[1],stage8_10[1]}
   );
   gpc7_3 gpc11111 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], stage7_13[6]},
      {stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc623_5 gpc11112 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[0], stage7_15[1]},
      {stage7_16[0], stage7_16[1], stage7_16[2], stage7_16[3], stage7_16[4], stage7_16[5]},
      {stage8_18[0],stage8_17[0],stage8_16[0],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc11113 (
      {stage7_17[0], stage7_17[1], stage7_17[2]},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc2223_5 gpc11114 (
      {stage7_21[0], stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1]},
      {stage7_23[0], stage7_23[1]},
      {stage7_24[0], stage7_24[1]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1]}
   );
   gpc615_5 gpc11115 (
      {stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[2]},
      {stage7_25[0], stage7_25[1], stage7_25[2], stage7_25[3], stage7_25[4], stage7_25[5]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc117_4 gpc11116 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], stage7_26[6]},
      {stage7_27[0]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[0],stage8_27[1],stage8_26[1]}
   );
   gpc15_3 gpc11117 (
      {stage7_29[0], stage7_29[1], stage7_29[2], 1'b0, 1'b0},
      {stage7_30[0]},
      {stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc2223_5 gpc11118 (
      {stage7_30[1], stage7_30[2], stage7_30[3]},
      {stage7_31[0], stage7_31[1]},
      {stage7_32[0], stage7_32[1]},
      {stage7_33[0], stage7_33[1]},
      {stage8_34[0],stage8_33[0],stage8_32[0],stage8_31[1],stage8_30[1]}
   );
   gpc207_4 gpc11119 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc207_4 gpc11120 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], stage7_35[6]},
      {stage7_37[0], stage7_37[1]},
      {stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc3_2 gpc11121 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage8_39[0],stage8_38[1]}
   );
   gpc2116_5 gpc11122 (
      {stage7_39[0], stage7_39[1], stage7_39[2], stage7_39[3], 1'b0, 1'b0},
      {stage7_40[0]},
      {stage7_41[0]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[0],stage8_39[1]}
   );
   gpc1415_5 gpc11123 (
      {stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4], stage7_41[5]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc207_4 gpc11124 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4], stage7_45[5], stage7_45[6]},
      {stage7_47[0], stage7_47[1]},
      {stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc11125 (
      {stage7_46[0], stage7_46[1], stage7_46[2], stage7_46[3], stage7_46[4], stage7_46[5], stage7_46[6]},
      {stage7_48[0], stage7_48[1]},
      {stage8_49[0],stage8_48[1],stage8_47[1],stage8_46[1]}
   );
   gpc207_4 gpc11126 (
      {stage7_49[0], stage7_49[1], stage7_49[2], stage7_49[3], stage7_49[4], stage7_49[5], 1'b0},
      {stage7_51[0], stage7_51[1]},
      {stage8_52[0],stage8_51[0],stage8_50[0],stage8_49[1]}
   );
   gpc1343_5 gpc11127 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage7_51[2], stage7_51[3], stage7_51[4], stage7_51[5]},
      {stage7_52[0], stage7_52[1], 1'b0},
      {stage7_53[0]},
      {stage8_54[0],stage8_53[0],stage8_52[1],stage8_51[1],stage8_50[1]}
   );
   gpc1415_5 gpc11128 (
      {stage7_54[0], stage7_54[1], stage7_54[2], stage7_54[3], stage7_54[4]},
      {stage7_55[0]},
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3]},
      {stage7_57[0]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[0],stage8_54[1]}
   );
   gpc2223_5 gpc11129 (
      {stage7_56[4], stage7_56[5], 1'b0},
      {stage7_57[1], stage7_57[2]},
      {stage7_58[0], stage7_58[1]},
      {stage7_59[0], stage7_59[1]},
      {stage8_60[0],stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc215_4 gpc11130 (
      {stage7_60[0], stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4]},
      {stage7_61[0]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[0],stage8_61[0],stage8_60[1]}
   );
   gpc606_5 gpc11131 (
      {stage7_63[0], stage7_63[1], stage7_63[2], stage7_63[3], stage7_63[4], 1'b0},
      {stage7_65[0], stage7_65[1], stage7_65[2], stage7_65[3], stage7_65[4], stage7_65[5]},
      {stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[0],stage8_63[1]}
   );
   gpc1163_5 gpc11132 (
      {stage7_64[0], stage7_64[1], stage7_64[2]},
      {stage7_65[6], stage7_65[7], stage7_65[8], stage7_65[9], stage7_65[10], stage7_65[11]},
      {stage7_66[0]},
      {stage7_67[0]},
      {stage8_68[0],stage8_67[1],stage8_66[1],stage8_65[1],stage8_64[1]}
   );
   gpc606_5 gpc11133 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], 1'b0, 1'b0},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc11134 (
      {stage7_69[0], stage7_69[1], stage7_69[2], 1'b0, 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], stage7_71[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc11135 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc11136 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc11137 (
      {stage7_5[4]},
      {stage8_5[1]}
   );
   gpc1_1 gpc11138 (
      {stage7_6[1]},
      {stage8_6[1]}
   );
   gpc1_1 gpc11139 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc11140 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc11141 (
      {stage7_16[6]},
      {stage8_16[1]}
   );
   gpc1_1 gpc11142 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc11143 (
      {stage7_20[0]},
      {stage8_20[1]}
   );
   gpc1_1 gpc11144 (
      {stage7_22[2]},
      {stage8_22[1]}
   );
   gpc1_1 gpc11145 (
      {stage7_28[1]},
      {stage8_28[1]}
   );
   gpc1_1 gpc11146 (
      {stage7_32[2]},
      {stage8_32[1]}
   );
   gpc1_1 gpc11147 (
      {stage7_33[2]},
      {stage8_33[1]}
   );
   gpc1_1 gpc11148 (
      {stage7_40[1]},
      {stage8_40[1]}
   );
   gpc1_1 gpc11149 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc11150 (
      {stage7_53[1]},
      {stage8_53[1]}
   );
   gpc1_1 gpc11151 (
      {stage7_55[1]},
      {stage8_55[1]}
   );
   gpc1_1 gpc11152 (
      {stage7_59[2]},
      {stage8_59[1]}
   );
   gpc1_1 gpc11153 (
      {stage7_61[1]},
      {stage8_61[1]}
   );
endmodule
module rowadder2_1_73(input [72:0] src0, input [72:0] src1, output [73:0] dst0);
    wire [72:0] gene;
    wire [72:0] prop;
    wire [75:0] out;
    wire [75:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_41_gene (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(gene[41])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_41_prop (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(prop[41])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_42_gene (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(gene[42])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_42_prop (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(prop[42])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_43_gene (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(gene[43])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_43_prop (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(prop[43])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_44_gene (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(gene[44])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_44_prop (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(prop[44])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_45_gene (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(gene[45])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_45_prop (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(prop[45])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_46_gene (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(gene[46])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_46_prop (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(prop[46])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_47_gene (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(gene[47])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_47_prop (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(prop[47])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_48_gene (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(gene[48])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_48_prop (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(prop[48])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_49_gene (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(gene[49])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_49_prop (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(prop[49])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_50_gene (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(gene[50])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_50_prop (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(prop[50])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_51_gene (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(gene[51])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_51_prop (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(prop[51])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_52_gene (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(gene[52])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_52_prop (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(prop[52])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_53_gene (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(gene[53])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_53_prop (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(prop[53])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_54_gene (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(gene[54])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_54_prop (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(prop[54])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_55_gene (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(gene[55])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_55_prop (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(prop[55])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_56_gene (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(gene[56])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_56_prop (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(prop[56])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_57_gene (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(gene[57])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_57_prop (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(prop[57])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_58_gene (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(gene[58])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_58_prop (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(prop[58])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_59_gene (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(gene[59])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_59_prop (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(prop[59])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_60_gene (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(gene[60])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_60_prop (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(prop[60])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_61_gene (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(gene[61])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_61_prop (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(prop[61])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_62_gene (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(gene[62])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_62_prop (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(prop[62])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_63_gene (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(gene[63])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_63_prop (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(prop[63])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_64_gene (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(gene[64])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_64_prop (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(prop[64])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_65_gene (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(gene[65])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_65_prop (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(prop[65])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_66_gene (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(gene[66])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_66_prop (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(prop[66])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_67_gene (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(gene[67])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_67_prop (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(prop[67])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_68_gene (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(gene[68])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_68_prop (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(prop[68])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_69_gene (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(gene[69])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_69_prop (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(prop[69])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_70_gene (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(gene[70])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_70_prop (
        .I0(src0[70]),
        .I1(src1[70]),
        .O(prop[70])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_71_gene (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(gene[71])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_71_prop (
        .I0(src0[71]),
        .I1(src1[71]),
        .O(prop[71])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_72_gene (
        .I0(src0[72]),
        .I1(src1[72]),
        .O(gene[72])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_72_prop (
        .I0(src0[72]),
        .I1(src1[72]),
        .O(prop[72])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_47_44 (
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CI(carryout[43]),
        .CYINIT(1'h0),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_51_48 (
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CI(carryout[47]),
        .CYINIT(1'h0),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_55_52 (
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CI(carryout[51]),
        .CYINIT(1'h0),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_59_56 (
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CI(carryout[55]),
        .CYINIT(1'h0),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    CARRY4 carry4_63_60 (
        .CO(carryout[63:60]),
        .O(out[63:60]),
        .CI(carryout[59]),
        .CYINIT(1'h0),
        .DI(gene[63:60]),
        .S(prop[63:60])
    );
    CARRY4 carry4_67_64 (
        .CO(carryout[67:64]),
        .O(out[67:64]),
        .CI(carryout[63]),
        .CYINIT(1'h0),
        .DI(gene[67:64]),
        .S(prop[67:64])
    );
    CARRY4 carry4_71_68 (
        .CO(carryout[71:68]),
        .O(out[71:68]),
        .CI(carryout[67]),
        .CYINIT(1'h0),
        .DI(gene[71:68]),
        .S(prop[71:68])
    );
    CARRY4 carry4_75_72 (
        .CO(carryout[75:72]),
        .O(out[75:72]),
        .CI(carryout[71]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[72:72]}),
        .S({3'h0, prop[72:72]})
    );
    assign dst0 = {carryout[72], out[72:0]};
endmodule


module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    reg [511:0] src32;
    reg [511:0] src33;
    reg [511:0] src34;
    reg [511:0] src35;
    reg [511:0] src36;
    reg [511:0] src37;
    reg [511:0] src38;
    reg [511:0] src39;
    reg [511:0] src40;
    reg [511:0] src41;
    reg [511:0] src42;
    reg [511:0] src43;
    reg [511:0] src44;
    reg [511:0] src45;
    reg [511:0] src46;
    reg [511:0] src47;
    reg [511:0] src48;
    reg [511:0] src49;
    reg [511:0] src50;
    reg [511:0] src51;
    reg [511:0] src52;
    reg [511:0] src53;
    reg [511:0] src54;
    reg [511:0] src55;
    reg [511:0] src56;
    reg [511:0] src57;
    reg [511:0] src58;
    reg [511:0] src59;
    reg [511:0] src60;
    reg [511:0] src61;
    reg [511:0] src62;
    reg [511:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor2_1_512_64 compressor2_1_512_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485] + src32[486] + src32[487] + src32[488] + src32[489] + src32[490] + src32[491] + src32[492] + src32[493] + src32[494] + src32[495] + src32[496] + src32[497] + src32[498] + src32[499] + src32[500] + src32[501] + src32[502] + src32[503] + src32[504] + src32[505] + src32[506] + src32[507] + src32[508] + src32[509] + src32[510] + src32[511])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485] + src33[486] + src33[487] + src33[488] + src33[489] + src33[490] + src33[491] + src33[492] + src33[493] + src33[494] + src33[495] + src33[496] + src33[497] + src33[498] + src33[499] + src33[500] + src33[501] + src33[502] + src33[503] + src33[504] + src33[505] + src33[506] + src33[507] + src33[508] + src33[509] + src33[510] + src33[511])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485] + src34[486] + src34[487] + src34[488] + src34[489] + src34[490] + src34[491] + src34[492] + src34[493] + src34[494] + src34[495] + src34[496] + src34[497] + src34[498] + src34[499] + src34[500] + src34[501] + src34[502] + src34[503] + src34[504] + src34[505] + src34[506] + src34[507] + src34[508] + src34[509] + src34[510] + src34[511])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485] + src35[486] + src35[487] + src35[488] + src35[489] + src35[490] + src35[491] + src35[492] + src35[493] + src35[494] + src35[495] + src35[496] + src35[497] + src35[498] + src35[499] + src35[500] + src35[501] + src35[502] + src35[503] + src35[504] + src35[505] + src35[506] + src35[507] + src35[508] + src35[509] + src35[510] + src35[511])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485] + src36[486] + src36[487] + src36[488] + src36[489] + src36[490] + src36[491] + src36[492] + src36[493] + src36[494] + src36[495] + src36[496] + src36[497] + src36[498] + src36[499] + src36[500] + src36[501] + src36[502] + src36[503] + src36[504] + src36[505] + src36[506] + src36[507] + src36[508] + src36[509] + src36[510] + src36[511])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485] + src37[486] + src37[487] + src37[488] + src37[489] + src37[490] + src37[491] + src37[492] + src37[493] + src37[494] + src37[495] + src37[496] + src37[497] + src37[498] + src37[499] + src37[500] + src37[501] + src37[502] + src37[503] + src37[504] + src37[505] + src37[506] + src37[507] + src37[508] + src37[509] + src37[510] + src37[511])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485] + src38[486] + src38[487] + src38[488] + src38[489] + src38[490] + src38[491] + src38[492] + src38[493] + src38[494] + src38[495] + src38[496] + src38[497] + src38[498] + src38[499] + src38[500] + src38[501] + src38[502] + src38[503] + src38[504] + src38[505] + src38[506] + src38[507] + src38[508] + src38[509] + src38[510] + src38[511])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485] + src39[486] + src39[487] + src39[488] + src39[489] + src39[490] + src39[491] + src39[492] + src39[493] + src39[494] + src39[495] + src39[496] + src39[497] + src39[498] + src39[499] + src39[500] + src39[501] + src39[502] + src39[503] + src39[504] + src39[505] + src39[506] + src39[507] + src39[508] + src39[509] + src39[510] + src39[511])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485] + src40[486] + src40[487] + src40[488] + src40[489] + src40[490] + src40[491] + src40[492] + src40[493] + src40[494] + src40[495] + src40[496] + src40[497] + src40[498] + src40[499] + src40[500] + src40[501] + src40[502] + src40[503] + src40[504] + src40[505] + src40[506] + src40[507] + src40[508] + src40[509] + src40[510] + src40[511])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485] + src41[486] + src41[487] + src41[488] + src41[489] + src41[490] + src41[491] + src41[492] + src41[493] + src41[494] + src41[495] + src41[496] + src41[497] + src41[498] + src41[499] + src41[500] + src41[501] + src41[502] + src41[503] + src41[504] + src41[505] + src41[506] + src41[507] + src41[508] + src41[509] + src41[510] + src41[511])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485] + src42[486] + src42[487] + src42[488] + src42[489] + src42[490] + src42[491] + src42[492] + src42[493] + src42[494] + src42[495] + src42[496] + src42[497] + src42[498] + src42[499] + src42[500] + src42[501] + src42[502] + src42[503] + src42[504] + src42[505] + src42[506] + src42[507] + src42[508] + src42[509] + src42[510] + src42[511])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485] + src43[486] + src43[487] + src43[488] + src43[489] + src43[490] + src43[491] + src43[492] + src43[493] + src43[494] + src43[495] + src43[496] + src43[497] + src43[498] + src43[499] + src43[500] + src43[501] + src43[502] + src43[503] + src43[504] + src43[505] + src43[506] + src43[507] + src43[508] + src43[509] + src43[510] + src43[511])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485] + src44[486] + src44[487] + src44[488] + src44[489] + src44[490] + src44[491] + src44[492] + src44[493] + src44[494] + src44[495] + src44[496] + src44[497] + src44[498] + src44[499] + src44[500] + src44[501] + src44[502] + src44[503] + src44[504] + src44[505] + src44[506] + src44[507] + src44[508] + src44[509] + src44[510] + src44[511])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485] + src45[486] + src45[487] + src45[488] + src45[489] + src45[490] + src45[491] + src45[492] + src45[493] + src45[494] + src45[495] + src45[496] + src45[497] + src45[498] + src45[499] + src45[500] + src45[501] + src45[502] + src45[503] + src45[504] + src45[505] + src45[506] + src45[507] + src45[508] + src45[509] + src45[510] + src45[511])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485] + src46[486] + src46[487] + src46[488] + src46[489] + src46[490] + src46[491] + src46[492] + src46[493] + src46[494] + src46[495] + src46[496] + src46[497] + src46[498] + src46[499] + src46[500] + src46[501] + src46[502] + src46[503] + src46[504] + src46[505] + src46[506] + src46[507] + src46[508] + src46[509] + src46[510] + src46[511])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485] + src47[486] + src47[487] + src47[488] + src47[489] + src47[490] + src47[491] + src47[492] + src47[493] + src47[494] + src47[495] + src47[496] + src47[497] + src47[498] + src47[499] + src47[500] + src47[501] + src47[502] + src47[503] + src47[504] + src47[505] + src47[506] + src47[507] + src47[508] + src47[509] + src47[510] + src47[511])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485] + src48[486] + src48[487] + src48[488] + src48[489] + src48[490] + src48[491] + src48[492] + src48[493] + src48[494] + src48[495] + src48[496] + src48[497] + src48[498] + src48[499] + src48[500] + src48[501] + src48[502] + src48[503] + src48[504] + src48[505] + src48[506] + src48[507] + src48[508] + src48[509] + src48[510] + src48[511])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485] + src49[486] + src49[487] + src49[488] + src49[489] + src49[490] + src49[491] + src49[492] + src49[493] + src49[494] + src49[495] + src49[496] + src49[497] + src49[498] + src49[499] + src49[500] + src49[501] + src49[502] + src49[503] + src49[504] + src49[505] + src49[506] + src49[507] + src49[508] + src49[509] + src49[510] + src49[511])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485] + src50[486] + src50[487] + src50[488] + src50[489] + src50[490] + src50[491] + src50[492] + src50[493] + src50[494] + src50[495] + src50[496] + src50[497] + src50[498] + src50[499] + src50[500] + src50[501] + src50[502] + src50[503] + src50[504] + src50[505] + src50[506] + src50[507] + src50[508] + src50[509] + src50[510] + src50[511])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485] + src51[486] + src51[487] + src51[488] + src51[489] + src51[490] + src51[491] + src51[492] + src51[493] + src51[494] + src51[495] + src51[496] + src51[497] + src51[498] + src51[499] + src51[500] + src51[501] + src51[502] + src51[503] + src51[504] + src51[505] + src51[506] + src51[507] + src51[508] + src51[509] + src51[510] + src51[511])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485] + src52[486] + src52[487] + src52[488] + src52[489] + src52[490] + src52[491] + src52[492] + src52[493] + src52[494] + src52[495] + src52[496] + src52[497] + src52[498] + src52[499] + src52[500] + src52[501] + src52[502] + src52[503] + src52[504] + src52[505] + src52[506] + src52[507] + src52[508] + src52[509] + src52[510] + src52[511])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485] + src53[486] + src53[487] + src53[488] + src53[489] + src53[490] + src53[491] + src53[492] + src53[493] + src53[494] + src53[495] + src53[496] + src53[497] + src53[498] + src53[499] + src53[500] + src53[501] + src53[502] + src53[503] + src53[504] + src53[505] + src53[506] + src53[507] + src53[508] + src53[509] + src53[510] + src53[511])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485] + src54[486] + src54[487] + src54[488] + src54[489] + src54[490] + src54[491] + src54[492] + src54[493] + src54[494] + src54[495] + src54[496] + src54[497] + src54[498] + src54[499] + src54[500] + src54[501] + src54[502] + src54[503] + src54[504] + src54[505] + src54[506] + src54[507] + src54[508] + src54[509] + src54[510] + src54[511])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485] + src55[486] + src55[487] + src55[488] + src55[489] + src55[490] + src55[491] + src55[492] + src55[493] + src55[494] + src55[495] + src55[496] + src55[497] + src55[498] + src55[499] + src55[500] + src55[501] + src55[502] + src55[503] + src55[504] + src55[505] + src55[506] + src55[507] + src55[508] + src55[509] + src55[510] + src55[511])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485] + src56[486] + src56[487] + src56[488] + src56[489] + src56[490] + src56[491] + src56[492] + src56[493] + src56[494] + src56[495] + src56[496] + src56[497] + src56[498] + src56[499] + src56[500] + src56[501] + src56[502] + src56[503] + src56[504] + src56[505] + src56[506] + src56[507] + src56[508] + src56[509] + src56[510] + src56[511])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485] + src57[486] + src57[487] + src57[488] + src57[489] + src57[490] + src57[491] + src57[492] + src57[493] + src57[494] + src57[495] + src57[496] + src57[497] + src57[498] + src57[499] + src57[500] + src57[501] + src57[502] + src57[503] + src57[504] + src57[505] + src57[506] + src57[507] + src57[508] + src57[509] + src57[510] + src57[511])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485] + src58[486] + src58[487] + src58[488] + src58[489] + src58[490] + src58[491] + src58[492] + src58[493] + src58[494] + src58[495] + src58[496] + src58[497] + src58[498] + src58[499] + src58[500] + src58[501] + src58[502] + src58[503] + src58[504] + src58[505] + src58[506] + src58[507] + src58[508] + src58[509] + src58[510] + src58[511])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485] + src59[486] + src59[487] + src59[488] + src59[489] + src59[490] + src59[491] + src59[492] + src59[493] + src59[494] + src59[495] + src59[496] + src59[497] + src59[498] + src59[499] + src59[500] + src59[501] + src59[502] + src59[503] + src59[504] + src59[505] + src59[506] + src59[507] + src59[508] + src59[509] + src59[510] + src59[511])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485] + src60[486] + src60[487] + src60[488] + src60[489] + src60[490] + src60[491] + src60[492] + src60[493] + src60[494] + src60[495] + src60[496] + src60[497] + src60[498] + src60[499] + src60[500] + src60[501] + src60[502] + src60[503] + src60[504] + src60[505] + src60[506] + src60[507] + src60[508] + src60[509] + src60[510] + src60[511])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485] + src61[486] + src61[487] + src61[488] + src61[489] + src61[490] + src61[491] + src61[492] + src61[493] + src61[494] + src61[495] + src61[496] + src61[497] + src61[498] + src61[499] + src61[500] + src61[501] + src61[502] + src61[503] + src61[504] + src61[505] + src61[506] + src61[507] + src61[508] + src61[509] + src61[510] + src61[511])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485] + src62[486] + src62[487] + src62[488] + src62[489] + src62[490] + src62[491] + src62[492] + src62[493] + src62[494] + src62[495] + src62[496] + src62[497] + src62[498] + src62[499] + src62[500] + src62[501] + src62[502] + src62[503] + src62[504] + src62[505] + src62[506] + src62[507] + src62[508] + src62[509] + src62[510] + src62[511])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485] + src63[486] + src63[487] + src63[488] + src63[489] + src63[490] + src63[491] + src63[492] + src63[493] + src63[494] + src63[495] + src63[496] + src63[497] + src63[498] + src63[499] + src63[500] + src63[501] + src63[502] + src63[503] + src63[504] + src63[505] + src63[506] + src63[507] + src63[508] + src63[509] + src63[510] + src63[511])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8be5c93c326905165b5d0a105d34f49c28f9cd3aebea62f8bd08cc0cc09f9f1467b539dca4c9a61a7acfbef79cf98f35c1ead39509a8cd8560ca3fce7734cae4189371c02d2d6e5d6126a513f5d6b7fd76ef1e2ac59ff31e0678d81fd9bef797364064fc7ad2b56c559caa32555fb51411e7050e988769d709766a243682064c34fce55759f631bb5a8a58c538b7cfed76e7d07c5b8409d562dbdd55d7cd65a56f04bf6f02d9faa7e8fcdd38fef807a514201c19220a22c75c5e5d0d08601cac456acd0cae30e0f3cf993e7958525a9caedd4955ff2f7a97d3d8de0922f66c5428401acd5ac7bfd7f606b1e5010642faf2d4ea2d0554bf35ca0ce435db68ccd36a2992dc570c870e5f16214681eec753a8e9831e7c8dd0c3d31d699e34ba2c5ca1d9ab990714b371843b1f78ae7f4c8ff5b70c8fb8fe0ccfa775e89d23cfca1aafb61ae25fe220946c114d3fe27cfa427cdd8595facedfb06d39222c915df75fbf3d08aeea2a5e4a9a55038928e4ebd82b2fc97135d272008001865d8ca146949d6495e6c92ba26b2e3ee2cbcacc4f95c0fab0544047cbe88b30f521b86d9d687ce9c27085d7f7c1d071d357602fc2be1aa4626f077a075cefc1a80029b31f88f88c787b83b7da81923110d7f20003571001d3d48156854947e747cd25e97599d69645fbe1a4ddb793f2ba377b3e48922f1c372a6ea1e922b5adff108e42a68513a8b77c3b3326ee7e07d574cb2b8749cb6b6c2f31b3e822b346dd32130956b0fef33a831d5991b1e4d86140cbfafe6fe60f625400939f6b5ea1b64e9e6b7f7531dc0d0421d77c2c0bbf09dc061049adf0f50f50cfb0ecbf04a1fdf85d03ee9b439776357457e4bbf2bfaf761bdb2b6b5c98212e8fb39d4be50cfef772976cee3f6e905cb3f7728778bf9ba4f9bd4591aabffed23c08014b058869503cdb106eac0b9dea187357bae270a1a1174004e02310484ac2dfdc2389433a4dd93d4aa255c665f5af92b71fe64e062634814e3e16d09f4904e8265a99eaaa60f56f17e694e48e38a4095fc9592865c365fa4de5760ae362964252019adcc02509a8990b6646964c59b3bf37b714fad765d1a1311fefc05bc62853288477ab98d82814c3bb543256fe099c30386a4458250382af82fdf47a9cf629b3eb083dbdf9803e66fee28aefda1451e29e81b39b0141b601052a2f92b2be0194a9b827ed47e261805a5597191c67ee17936be8be5b4b4c2a482b274b9df734f230b7dc634a919afe50a83328b30d6d1f39d2b0db648ee89121de757ac9c2c239eb83dc4fa15432b2fbea8e8b09ae0ee43136b30acec92a1c083d15a748017daff47777f27d24f9c301a034e75b49b21c694ba525354bb1e176027e8a65e773037854236afbc6b9e589134528b27d7a16201965669d2a09db3c51e475718f08843dbf76c8ae21fc2ec0123cd209d76f777cecd9455409f8c0ab4a9ecfa3a4ead815e3eeeadcfd4941107c775a5aa851ce2ce03a1d8ac5d129f11415b3bbbb2af43c26c6e34fb91afaada1eefe7783fee763e9b0a9726fa640453d7784770e9c7bd00ed4669d34f2121fd3c9afed5a8c68cb189a3a8bcb32b7cfea339721947a5130b090c7ce47749d317a8027eb760e83ce125835c1d67208fc4eb4bf6355bc8320f856f3344ccc5e94d5d79cdd31f88dc735eff7b2ae798f429fad9074ee0e00e7d66c216352dba412ce18fea519b8e9c4f73bf3919e910b4d596d975d92a7b9289abd94bc0955115afc3c4433d029c0378e834bb5717a58fde24d09fe4e33c8d7dc0b744d97791b045b82717542dd120ecea8ea652d54df6d2ec4fe1e55329fdebd0541527d3202b28a115fcadbbdbf54b28a6a7c63936d79c1c3641376b7649380466952f0f4ffb3725d68264b889f8245af739761fdae4dbc1eee36171bc1f1eb3472edc855debb8c9a98eafb99113cece51752ba580bac222ea75390def512059362963dcf4dd41ad0a4f68b2e46a7423dd69603eb94aed4d340ae7eca47c7400fbd4a8e70c547321daeae46c9ad572896b6b6597900f15327bf1ddbdca8c3a89142e4571e3f0b0ce5930ebc5fa5840d3e2d1738f9bf7d426e865e06bca72725e445bf35d89a3d0d99e46cd2c86b3497c24bc6e06085d4b6fcda485b62c433f7aea49e352b5e02788eb0a5dadfa2944a5af0400b5c99a2431216cb01fe9f528f85ab7f7eae658013e2b66ca630ef57c1e33968a8a887502647bd15316851e8f26ad6c838a45f072b462f3a24494ca91778bc328c14697b93da0aeb632500712268614e09f89e06c87122c0d4a6ae66d88faa370fc91692d440d08678472af6871d948001fe49b57a53063aed7141ec09baa268abfa211cf1f73c2edd6ec7b2b66c62c7f0eb0b1682edaa7e660495318a695871c88f187aa0f058392f49a5cd7250137b88410e8f00e9f40b92bb198022bb4f922e18e3fd4837b4bd0d0a8b1e5bf754acef795c0998548a5c04e7f5eedfd1e0f15118f9a63923ab5ed3df731e9f4452d957c8ccb05a876325749cd5ae78f5da5181ac85bb7e389a237566016568ad3adb4b589e317737b300c8d0458f5f6044c6b95b10e2752c54a5bb65b0234d0e0765cef81a2876425fb6a4ba44d09b075d171d3b7cbfe0e9769c7c04fd3d895f755532b4bf7f055e0e5edb4d9e51008a2388607a1b0cf5ef5ea5246f96c9bff9e96cf56249379c6d01672bbbefcfda8f47732b6fa0678c3f97e3ccc33d87e082d3612c945de87b93a25e727694cb427d0e1feb628481a2de718cfe53f1d8e2baf5f8d27602e6a1eba94d147454bf494258c3da95db447e96a545532c01632651b78f3da5c05b9702ed9b2a124d2aacfb7f84e316aaac3eacc7f20489024662b83981e0b1ae93b7d86dc7fdee2a9f48fce5e9c5d281f6fb53fc04de963837d2d72d4240ce14d44d4d4c416ffbddd55c904cdc74016d7587162dcc9abcde7110b1bd6aa417a419890552fde11df661d09e44ca44344e4ea2c4bea1feb2a1d45764c40be319e30cb1cd7560a95dd908f774bbea1dd268d7182220c6eee6346ebadaa89f444a022abac0a32e28ddf3fec6f09faab1f91ace27c7ff22b0941824f5853303c9e70d64f2a99355fcfd212613c8f85659ac94d5d8c9685e835bb5c73400ea373500ce65ebccd3df663a1fb145e20850698d73d020d2258114a841b8b97a45c771de8ea5d811bf1556c45f6deeaa30c9b794810a8eb56fdd5db29df6e298bc4de85c2b0a8a724243b87838f2c2e34c7aaadc5a14179221286977504ca1993dd8ea6ac2899c3ae3812e380dd8d75e6ef347a0248bbd81c42f2b119783948405c75f008fbda76a26f9a9b8d30a1a7a00d5b6449631d5bef148eaccbc94011f560ab61590c1824b540b185cca7c21f7bbd154c216ff1b21bfe58e1cb0bb86911881834c299f78258faa38294cc48c2960294f2193b9079d53a5b9107027d7382a6195878bb751e8e4c9490dc77da11f2b8bfb486cb01cbdcc6d592bc68de2dcb4ecc68ee8b8d8fe15f4b42c3e4b72190803b5933adf675f23ea832d34797f06a46c3ff8256d20e2577a03507a8acffe5c4bf9b83ba47b3fd3425bd7cf0dca3afae2b0be0d9813fa24dca6396f61e9079d95a15d53125316abc773dee21fcfc6c7083a75f8d7ef8c83aaf6bce3816bfb84fc723b93b4494b56182c3ce6d16e06510c3d516079f121ca162fb40ba5ee2dd05b9d418977a60c2e8061a5128200eb4e3b9c21b5123a4344acc7fd1ea911f1bee33290dcbbe4d0616788a2ef4a852e586bccdfe989fa810bf2424cc3db223629993bb132b4b1333e76f89709d7ad44e925ade16a0855d013516338fbb82b42a40adf08b6e821ff160157e591ef69d9813496f96e8bda810fd30ec9748bf14004ad23d3950eca0013b3d4d1c86f655c7d5859c2ba48d80d3410e6d6ab149628b142462dadbec02ac2d5383c942e1ab3d0ab318207849a5a777b970a0c28dff9d8c800436221b29eb8dfa0266f0c0ed841e4fab1eb98094243150826f53f5f511f34cb279d4227818c258b5d53fa407263888d0d5869bda47ccdac32c47c6e0887f19430b721df0c62953d348d7ee80ef05e7c85fed3f4b28d1395ec347749e49f6e5bebbdf17ca23c878985380dd48641a9b0f621eaf2b57a0e756e90a26cee13ec8600ee50939ef582f59382fabd221ed2b87d4ee56641afce4bc221f8df454a832724953965f12903b36aebdb09ccf8e898c124a3421971a8a825434b7ded016b0cb3e3d4183c6dbeb8e9342a44289f4883e051db59ecd567e2f6aaf2b16fe16b529337604c8905ece511c4300f8b9640f75b05c5dd4351ba08078d64c83a642a9e8be600a992f3e56cae409e877acac80b7dc6a3bde1637bbca9d2509703bd4bdc3752762045a4a4c9ebf7a760efb83ff388e581f1a0b1fdbdf4dd75f789a40c03488ff9a56eafe5c477bde4868b374a005214cfe7afc7bea5afffe0eecb9adede8a108688c743af4fc47a60666d19c5af98cb274661e0244ed8eaf568eb2c3d21f5a959aec19487b39cf9a8f082410f57046ec52a0d2fdbbc55aa6b6e6ab2fbb6d7b090fc37b96f7df827ce8b462bd31b33736383fa4445f5ddaca33260e4610d83d5d6bec0eee4e01a3661da16a19de5619be16c53ed7a16dcef770e2c8751c7e237a734e98856ba60bd1b394962ec8a287fb6448bb3fef32c54a4bb3403a01a105411bf52fee11872a61a22a3fbac58b06bddaa280092e4b4dddde4cd69120a7a0c698d62a3c84371894bebdfe4d3bfab2ec35a3ec6c01299c2a53283d4076daf453ab548da512950c7a5736bb0a258243a4d8f1acce1934f4fa529efbd20519cba2f3bdd2d389fcd017ea7757e425cb4fc0a56461452afbd8c052e701d20bc4cfb6011864ece62d41a80db93e285caf7abe3ce9c00a49dce475a11358888401630b212f5bd65e3ee7c528363b8e2e5c6ed76d7fb51a8d3906c747b20db37873de180343f150ce5c61c64ede352d34728b68a32e8740ead91520379575b597facf4e53a0d79aec7065ad82d6f23582996568a155be67e70bd831b42b0a4b5c3ecfcbba984b706efc8753db00e7ce5adc2ff7017bcd5185bccfccdbde0a92f8fe1aab791b9ad35f4fb12fa7d36f8ae8a5b8e5c2e021eca7973ee3aa497fac54f8a2b564cdca6736c765ab96976f11dce56c923abc1eb11dde7f374cf05b9d02a1d4013ba1dc3c0563f8dcc7740bb15a2596cfddb0218475aa1f1fc483f597acabc36afbdefc06e55c632957ea468a4f88c2c0c29c79f16aa57eff2d550b6d9d4180b5d96faffbd0f0ea11bed9446935f957049a3ca03372bbb22714fb65e99c3dee7c7eadab9235374927f7af8008a38aa5b597c914aa31faf55219a9be9e0e04003b37130fbb4b482971518b85fd681053eddf7d1278a377c7c2dc13a72d42251966151455b55417e74fad398581cb9ba188388a82b2ebe8d492169023cd700a90175a7a1a60e5ec5e3e5d6a315412e86f4598da6c973283f7e53001cc83349fdfcaff0f869fefa13fae9929610926615b3dccc542da469fb5f78c6bfe3f1b89901f83fd328147e6a0608741d561cd5826cf06ad831011a5a226655bdca29086f9a1c36061d438c0ec8cff4151216245d6a598b1509c1e724201070e0be6eb5d1fee6f06d8ad067d6058abbd39e79f84c972309727da80bd7ec1180cfd74bbe010f9ecc557d547b2906ad5178bbcb8ab393a20ca5a0e7481442febe8d7d2ce527f9e3b6ba9f4224e367292b48632c64e24;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h374b1859a76db860d05a0aeb3a8430f3862403864104bf24570caf47076a40deb971022bc5a7728e4efcf434627dc43203c792687b6ba2fd0448fd4301e15d1dd56e6069cd15e642752900cafb97665da43c656360d13a0848c41bbf77a9da4440df8b8595892d373e7735a0a3e8385e186334e10df6fe542ecdbc119bfede62ecc75a443fa7a690bc7f3e8238cba851d85d1b1b489540c59f03aef64746239576c0194febcbc355f3cab71c32b45361e5bcbcb2da1800585b2cdfeb45e09769a8fe4501693fa03982c1beaba337d9d46db22e552a08374002ab0288878f7f17db917dfa21d2da7b06ccbd4ed529a674599c5e13bb5b1eeedb00f5fbb70310fedbfbe45fe0e6fc385e45dbd78573feb74e9a71eaad9aaa69ad447bd249e3270f9dfd3cac4acdfbc4f6c838df48f5775dcfc92feda0360dfd713bfc0d5a4c6a23ccc947d8f672a5f2a249ad4c4d87e732366f0de22d98e86bfe08019a637728b49f745b3c341121509bcdf3ec5cadf051b005dac632050afde15766556e1c9a9294dbffd0301ec789f907703685a336a5432d4789faa0ae4d4219d8374bb15be569d9606784870537c2e42665225be109a51d2706104e06109464395f8885adcb094be794b71e797bbe0f6c8eedace31169ea9d01abc3aec722cff2e65a679a00653b2395c4290825cf5639b5612d0e139e8abc79772bb04cf9f3ce764fb2fdce238b8f2cce93b25eb5a59ca1b916b98027395329bdf3ba47c0dd93f31a1c26b47fe617de82f8df9d6c5c49bb71d5cd0af9530a9429487fce27b4f9d5e1b189d64a58a7daee6e543bc77d7879b21992ee67f98e2ba1d186e487b23dac54e73719d0cc9a5a39701bd30f2dce9c9be158c2edc04a3c52f5ceffe1cb851cffa11aebefa1dae6b4c400974ae9648b1cd41d19c73645902d2b8a44e0f1e03c76288195fde905bdf835c960776742445a9d249bc336ccb7a000d6cec8828c92de4ecd55441282c597b716537a643e5dcb0b81bdcee09435d6f8d13f1c209a7f730933668c08da7ddaf8d7434954ad86027c7f6a8ad05ae5219b4d7bca7b5122222710b711dbd56a37cd4c7d32e54d95afeb1991eceb641d66f189b4a970cc7e475b091ddb68a0db38e15c9c2d3dab2c1587da06fa2b5c0f1a7c1a6b786d729a1beb5a6a431c5b06b416f60b083750918b13db0913edaff21476135093925b98ca9a2306f623d127ae1f911f7c1807a302dae9beb29694b459ee558af23d1597c407d54036df61399ccbced89803dd95ef33abbec04cb131100916bd086938d96befdde1056d23dd155ce407dd6c612394f11391be3cd8a9c10b26f9fc8d9b7ca17883ed1bf76146d269e522185436bff546807c35a2dae4839bbebbcf73acee275167e7ba4f9c4cc60c2dc5f1c1ffc4d61d82b46ce4b24fc99db65c989513ebf6894e381dc697097a69dc19048f2264419e6a73ac287b5cb8dea189d3fb5292889d489def90bb5927e2ff794a151ee71975a99812937c322941040ac6405764fe128c8054adc95ebcac319c381a1ff94e1986ee624ed0ccd97ae4c858a3d12cb590cda837c853bce4af5d1978b1fd4e2d9f4084fbcc6e9bb408177bd4caf38df6af65e3c7fde6258865acc328ba9781bf0249285c3761487bbffe25290c415d52f550323a19237cbf74cd675731d4b09c0ac0c6c8f45b0b06f01d7aa6dbb269304772244298ead02750fe6ee3be73f7bafe9c8f081557b4912a816a992e0948f87f3118faab6ff0bb6420394964ce0e2098da0e13ea187923a578c622e5df48119090833956d34b9404638939cc343d7d6bf6d7a8966392dec7603177e7f990cfbc2f2b1c267fd3936a937741755dd044a3afd6baedb63f60fd7a817f3352ab9645346d64ef7882cba61b56477b3102bf7e376f7ab16472d97b28ae56ad74a17571668c8a5dae1f8154f4fdce8cbebcc68dbb6b50c32d1f3813dad229b4aa716a2a3ecdae0a019c382632d157237114a994d4da874b5c4ffbdbf10e0368707e13c833176ba1ea6db7e5531c71a7fe6710d46c0d35712ab67d4a21cb7a5530d3b2d28dc3cc6816a1fb5b36131c00ba167676749b83585a5f84fadbb2fd29a78afa5ed3b14da4482292f5ea1a1923c6c814a1cace80a985fbbddc05a4769c06fae7814cdf936be64df605e935c774a13771bd789d4886326c5eed3f398c3502f56bfaa6f16c70d1cc4f7e59c99fd46f68268ea4ebb5b068078bbe77170772cea68f393e64f1dea72ae6130a92331869308ddcd48a95d75f2796cd31b4b5e9e06b67a85f5c012861174ca01061a0179b976a80549d0fbf43c06c9ff671b4c6f65d3abe19d61b7f4945290d7bf580f66e0026e027767749eab29b103ec51d475412c28dd3250ef9dc35972b36eef2ae8a6b2adb3255d4d942cf365a1a115a1049c177649b22eee16f9f97e90e0d0487c644f5b077c5de6d450f15ecd2df90c45b7ef5c3702a1fad442d76e581bf1ded84f08fe17fb4fdb90fe95b197c4e083409d64c0e59a36cde565f8bf84c41c4dcf2b5a1cd5245565dd4d3d192b606d2faf57bbba9a210410aabbe0dfd9e1c76c25b7c169534deb735e4afed1cda53343aa0b86ffd502f4aa56b493e55613d9ba2d30ace23061b85b3bff64400b73beb45fb14890eabc2fd62bdef649619abe10f01f59571e8103ead6cf79e92306271c2450274d05e5039ec69d7bc3f207fa0f833d4b292e5710cfe8e4e62792eae1fe49edf8611e752e9be72e52adeb1236f4b2b6a996a0083c4f55611b7c275446fed19c8084a3f3b923b05f053fd39fea8305c282fcaf1e8b634680af344b50ea47fa9118dbc5fda6c8e603c12487bbd3e8be3f3c99f2e240a39ac83e7465c136ab9233b0045b7d60d237d896ac59e72e7b4832cadffbf69e2af873578ac995d5578d117fcb4f95fb871fa46b4f59a6a09a7ea9d8d8d7eabf9c8683cce6dad26f964b3960ad4c8b97827a6ccebcaddbc54794e937be23419cb73f42f4e505cf07eed047454bdc27f24ad04d8cac6753ebc080b902a3efda95300d10da7e6b9c6325669dee53b35e4d8ec18086bee58437896a1fb9b395425ce52748103c5800d3295bdb6d1dec603bba823f091330e686cb5866e08bf67ea26c6a85fc41155b7fca75dece37766004c30fec71e1f08628c7201cca691f993a86ce8a82d21c35b4ec46b99c3dd20c100114625fe36b758cae9448c0363117dbb4b0a221bd538f7e1ac90e9385700fee398cad856d9f0b287bf5017726cd951984b392a98c0480450f9d7f84ad8d9f70f4cc6b073eeaea898e10d74dd45ac3abf741fe52c79fdeed512df20d0e0034f1932e06962fbc4f01fe6669106fc83eab00224ae46df60cfa015a4e2db412a125b5496a66c988117a4e60331c8627abd8f668401c3110de77ca6efeca233eeb5373b0a80885ffb930e44b01d25ce90450cc37997ed47035548d1c090b8b38c6a6dcfe6b55d467ba1f01fed0c236dbbcec7f910a5a9f3686de206161e3ace1fd37fce27c10c377a1bcaf9498f38c4368986b23a79f2e05b10084454e90e0eec37ee34709da89ff847c26550efdde70c3e9b65096081ea12293367ff540d582b7b57e01bee6db945d40e24650f4a93ee8802ff4279c77fb1ddaf2d5a6d8b607a5b9c9ea572f054210ad2c014e5165664d244941a8775fc563de2bd551b0762d69b55562f99ddc5a8b6b74845df62c6255cbb2030e0c774fd32a47714c35de2181f1a21b56bdc438c78f36315bb8b4375f0bf72b2187cc7a31f8affe763df4af26dcdf91d3fbaaebeb12990ffdf0a26bbf1d35b185c487cce3f8f5bca7bc2272be179fff930816ace4112f5cd2deddd401c9e3b0a4a8f0ed9803c243cb91aecc43a62c33c38ad3b9945cd2b6ba01c9f6ab2a014637dd67a8b7e44a8112fdb595df865f3d8fedf494c976da7dd17f072d2483c5b321a35f9381e899ce53728d23e125445d5af2eb8b0d31ef4820e31dd0b987ec5a81fd413cf66d2aab54455c662717f542dfafa4227e3cd6e59cc4e0af74308f5d678174ddfd05a0fbb358029ce4ed9cd8b01f8527efa981e025c5f2002c4ae44237d978ec3dbf16bd64179c89fbf8954aae3fc04b5c5785eccf4728f79ca296c772fa56c3ba9946c2a64f4aad654b39f71307460dfe261d47986af9df930c8457bfdcace164969949b69ba38bebb038400603e7a636088b06d361d8e83487b0b89f2e11a1070fd9ab389cd7953af44170a4a2ec8c75318be4afe4f63a84e473903a118527e45b45c737e956d1d767038878f487f18e7e3b97f9c8f625824bb254e15a823a273b42a9c52c1f0a1fb0ca4807b397142897608f8d2a34bcd274451a1a23ceaaa66f7a958aa2cd3a0b8e98d005e26c746b93c0c26cd5eb38f59b3fc4c55eca2321d66e47878f261cfe15f5e67011369e9af7ef2b814d27c95a9e40f172dc30d06efaeff00bb0215241a2d396d42b672d8d723b9b0e3577f067f244ad1343a77b5d5c8f93cdf97b4d514c03b28c5e1b412ebe259cd59bb6f572ce74e89f93e0b09febf7b2533dc271b0c44ed801e70b1dbb46f8d4b50c003a543d60a230d79e2306c97d3696018112ba0fe73b8c120661343cbd3bb364cce2862ff61c0cd667692828b01f5d627b6d5bb9ac8b508691cf61d1b9a47b13442dc7e61f8da59d01ec8eb2eee2ec36ba3132b3ad9c70332085de1d1e9bb7ea11c54f2af9be862ce26ecef72d6f07160671adf6ec3940f3dee42a0126f923ded81ef8346a815195d4cbb1d01b76f79542c80fa56f58df22777eaa143b7e31116d2c6044642e384c74dde935eeea5043f9b320f48a070cd5ad910ef3f49a2e4d5b5be817cf61a0a80d4a5498b204feb1d43e8130255dfc2a6da76066b6e0b0b013756c50b5fb2108634c5e63868a010e76db66fcf9fb4c0c60688768ebc5dbf93bc81d8c211e4aa3ecda35da375eb2eeec3c2f9859f2f11b02af5659f97d3818d778edc2a72d766a1f4081ff4ae8bae4f265c12d9545f9d051f197980a0ead71f28b735787703468a5da76ea4e6e0ebb0d3e8f92b97ef170e0a70d1432d3b140e68e35de35562c7eb69e10d9109476bbbc540799ce308c7fa5cf045936eb237f70eba0f190e37b2fbb5a106a9cbe660bebf03a5c5e413f19ab04a9fd4a232f811b5d782d35faee444fc433f514fb724f20aee67d9aacc10289b97b78bd51ef0856f5d2f3b49c5d40fc6ebd3acb3bb4fe190e959810de8435fd4678c04992959b3762b8d69fd18d961fc4167010e46e8a6431d68b8e27271d34cc482523b99481c6e8e49433dd765436890da1a578af4679c541e386014a32831cde9ec55733aef730f5a38d021002dc63df84c81132edfb896511439891a0b4109bf2b246aac5b5a207710a888d3a71a2e432952440cfb74b453c3f9eee6f11ba6d82bff30dc10035ac38ee3a0097d9997d83a81947f4aa581f34b03aa7073e880d3e49b54a12f0ca44bded9f1f473928ed4e5a0a997d8b939860f5dc7047a3d80cda1c5c890ea4f8faaebf0344b6e788ee2a92d598b84017fcf145da23f6451a97a25263663d8ee0e80b45a477d0f71ef4dbf5057f9f0f4fa735e3cfc5937429c9ea584e03178c819a4ac05c66d22e27cdbbe2b8bd6d4359bc27798349903c3d837004fbe468f180c971c2645b2760bc1307f5da1b1f63dc8deb4dc810212bedce1c7186c79a642c514d4b6bc3725ae9b7b9cfefdb62f6ddac3520568892d4296c928643da4e39178600f6d71dd01e304a0022ad63d106241c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'heaeb9b161db7b502906bb60f306a7402c3d5d6d2fa5c27553c1ca302dc7631a77afaeb5a84c367c33ae858bc7b76f029a2143a55f17951e745a2153794e6996ecdc50f2e0137cb6245ee64cb167bc9dc59451c1b32ef023237cd2aac851f4ac3fa8f2cc38948a4de1d9371477bdccc885bb1127fd7e8cfa6fa49c89cebe07c96faa25aac0d2a7a9fc70cc31e935c3d846923fccb9f35bd878fdfc24b241bb1132703e9bd077d204d50ec497281b7d7b79c418556b619566f68d1939fea5d703083a5327a1cb8d6a4c7972fd3943cf506edfc89b20f194b1bb727b95a4d461c0b98bdaf7c2215fdddb09c5e126f7475b81c3514b3840521cf5d681bf2b8a78e8bc9bc816d8936b8edb0cfd6420ef17836601c5fd00bd107d8d7dbb328d99bb95b28e50aaab5bdbc41ada4c9846419a729b6acb94d7db081d5c56ac377ee5fc0de172e0905a78e6b69f80a3a9b058b6db3c9ec744478fafd28d4568a1b0315feb3ad255ec553746706911072e0720d07d28bb8fac75536ac8793ee0b51250bc8baa656f666f6434f0741e2bcb69e40f291a5cd298c6801bbe4879d240197d2bfa1aead92417d773bbf209b020fae1fc6d662759cf2b2b71c39a45051405b105e2b0f00099b9b09bd5f1e8011fe9201434939b86b912885cc1e6979295fe591a044c9c59793c2113dc0d06e67f5d852a287054f9e2ac02fa1ede41f06ba4c0547b2b7f9959650078f3890bedc0bb854d7f56b8b15d93b1aaa072f1950a8c3be6724c6f73c8b39ab9aac26c33534e97a041028e54c2eb29b7929655e18939e61b882dc40686b1fe599905721ecd6b09a29a2081a177be2db9cc5143154c6808f73e41ad6ea2e2d1cf0d2c82db0d0cf79fda008494e22f0f0e24a156654d2e6c13acb96bca057cbeed8d46b0050e13068cc8e78d9f55f3b0df141ff950154ebb6c7c1c891b3a87c7ff8b0ca97c4fa0dce2820e76250f54f9961617acd1d31c271e3e4ef1e568fa040e1926144809a74600112fd5e1812e3dc33567894fca946c6e82ed3158df4d18e2b8bd2f8c4435172cb6d917feb2ad570759e1010e79d4dcc1ba54a67da0ed1cd7c0b3e78d4aa574f951075d31e4456951009b7ac536b1dae37a0db2cb5312b192a44ce26825e4102b0a2aebbefd1835c2552a074bd2aad42476cfd7d790982f8ba5bd6a58c1a77bafb465bf8c04d0519b12b0f9a4ba4dd6059b87422857ad4bceda16ef3a3b5b1e0844c2f9a9a50b11959a02c90fd316b0ad32ce808aaca902230b674993958509b1934589e544d927b2c2e4a6171f9507d591c558042dc31beeffd3794809b02bdf34864c5ed9b89fe41b5c8d612e542557e1087bc38294c750aaac4fad8cc448700e723e4520c902436688a44c6c6a644293aea93957fbec4ad220703c31e07dd6486162793f655a42c8e65124b0aae65fe94756bdf492041682552b5ab039f334adceee88a4facb39ae1d5c18e55a457785ab0a172351d4909894962ba34fa18c8385b3608561bf8f77ea5d34819bbbf7d11db0f8b112e4ef1be8d366eaeab9ec89cf638f70faefcb990d39c6891d674d030ae0552dfe3a998e3fd952d0a9fe032899cc0532ef2e51e85255c89e42ceb7f01e43f4a7e8029f2f98fa5de7484e5e58c9c9fd48aa32f761be79a0b77898fefe599ac896243d9f974717b6dcf46565246a7533e26965a0d241c460dea7d31995d49d6b228a74fe71586e37ed4808fa437571d36f0a6ff48075b74aa340ee43fc361f934c24f221f2b2aa20139c85e4a4299384b9c846b9e2e14d695ef08adf8abd026daedf8e8313b79305daaec95aefb7adfe1feb88f806a78a2eead02c363d1e46dff541dec5e35108e96724218cf88c8e5c32d660734de21e24646f056d629da17b00d48301c67103720a63518a6231fc5d72fc75d530ba3d99cdac679e3016cb024f6852ff9060ff8cf9e2ca75862640df9130a6ce1d5c7558fce3a37a20bd5056a566bead8fec75e0347367eb52f384ffac1dffcbfa68f2287eb21e10ec4479e81c68dcba5aff51a292d61a90656edd65ae0cd51daa9d7068b0fe1174ce69ffcf508f9b7ba0538d5b7dd66d9ef5547ca6f542e13358168f3644bedeb047da80ce970f7fae77983e3671a987328b78dda3c4c0b6c86cb94e264f5b98edbc56012cfd9610b9f2698f21eb699c0cb42c0ecc900106350a683c20c981f06607f43a23d1d604e16c12b267827318280f505a8493f0ea86b719216c9033fd07fa48e9c4bbf730b051f52108767341fe8c87c65f1321f8d07a227884f752ffc99c4661c2ffd68dbbd03f531f3bc1d7116365932d121718402c33ec089574557f2e56857f1f6cc18428b8c97136cacdc1e1bcbf6a39ed221e6b36ca8aedd0a489935c9ded8d7d5b2d1ecf3bddf0862aff95234ae090734f7ffbd612cde1ed428a36834ef19f2aedf0996737dec6add5b46d9c41224d7ed044430c74b95d52caa517d012807689da5ae67798eb1994f1b8b4e4cb2f3c256aff65bd563c0d7603d0057042f3612474e169d8b29c8735a95883d3d642b1846fe7ba5980bcf9613516519ae720f1470153193eb4968226e3931244e2d8cdba5a0957ee99cdd45c6e679da3833702804c2f22c8d8e9103b4dd59bdd78867d27d091edc0eef6c2344873f94d01afc33e823232992df8cda88f4f4d703d7d325d127f1ca79cd68a435db2e36401a30243b82fca53501816fa053f5ec77b88ba169b0b45f6e8b876c9ea49da2ac438986d80112a96262547fbff967a137c9bf668a594c9641fc9f40b2501a3093ecb555158e11b6aa933acfb9cb592e564aa2a1af5ba81ddec0f0fcb6ebb2c4de35057adaeb86c704f079d11aac0929bcbf0aaf0db0e7e59df7988b60319c9532ce1d51e4d3148b8eed3e4048232a1e6724c814ff3210902534f7f1387e3cd462f67a73e8937758f658c013bea0d62bb123e8c8cd5f7b3f838396ec15644a1df49800650b9821feaee0c4f0efb5160b0fbf52d7f70f1ec785227053d9a4113422441e08ed1aa4a7a3831031d88f4b5e5448de7464916557ed09e7864556a96eaa7a7076e96ef65c20990953215e0b0547de9e9eeb39a97f81262d3c50981ec00fd64a22812e5444172d1a3bc427ca3786c8ca5e89b2a7d9a7ddd0b42c6dd7c36927d75180ca505583fd12bf0ea97434fcc62bda8aac83c89e5d232a48514fb9705d587feb001ca3b9954d78dae0fbb0ba85d6211e56964b03986f1569a09b27a15f28e05701acdc178faeb07cfdbbf76793d0a2715edd6b1dbdc79f873284bbabdb0107d7b75f6e12cd52f75819e75d75deb53bb3f06770ca3215a0b92d66a4f935c0bd1fe485b68ffa6f398a530e98deef2f71db397467785158a031828cd180bdb34c57d280daf0f52b514159c384178d0e689c54fe19020e9c1654f25dd0860a0d59fcb2a6a0f41857f691bc4594681db8757bf976d12ed8c6daaf36915cb2c86218206f20ee035e133e02da0f47d921c92168fd34c4106780181b9be59adb0434599ab132e6a12d84aa21217e815cf2f14116c2891f3972bac794efc92ebc16f1a49254878c6945a69815814f5833601f264241a0d2145bec4fbe8b0e8397a9dc5e8130beeed98ef74953c260321f7c74e9796b9d4307a06ace00507fb7a84c7874d93a69c659bac49eb650773ab1b897f0cd9ba491a17c78cc4e95729e6332cb1e502e822b01ee55844cd1b4ac38bf5500649b2469a33ef1bc02170d91e599ade694665698ff5f21b911d15f04971071a1711c794bc5251cd2231b0116a0de95219fb8c5cf60dbfbc86714d705f78a5de474818d869472ae7696ed3f7ed15e17c87fd955f773271365efef96e27b7da1334e49742439396c238844fe7f6e59239fa5d222253c5806201e40a1a0cf1bc68c0c7c8526850e178974d1b8a74362a673be3360328f2cf9702b5f3f2a3a0ff0d9f6474cd5356a8782c1aa984ce8dac04c72e914ebaae3b24950f021b6f41d085380052edb478999adcfc912d2e4008c936f203b7ac9de4df323d66426b92aaa9779e274af18691826d84a0bc95273d5a15eaf72372757a14fa1d516dbbd22cb1e41aa01bb860f5298b60e004b12235de5820e1ceed3b2faa0c2b03f0a4b396677818d148f972abdc355f80e90e04a6d94456b19ccfbc69ba966b717ec1bcb9438788180b8ed96d164703dd85d6e0d912b6e35da4c7d62c2484fa96c0706268ef9acb48a4c76e7116dcc02eab077cdcab74c9f694f552aed4db9063ece0d2c8a8b7a6396fe0bbf463dd9e21aed540d2ca5275a3937b0a9ad2ae1338e37d5d74304f03cfc44080ebd66b04fe723b616c489931852622ed7ec40679c3713187dab0c0a0bdd18505c9ddcaa9cbdd44e80926ca6486f0431f1209b391a8cf88e4a1bc454e6b0f4416175287d3167cb8e1415adc8bb77828b6d03a2ef2971e52ddd5c18cd54b012c427ec8d95bea6dc11c5a10453dcca6d3d25d3e3471fb9af126349344202ff3e284c90a4b0813e2e3f150a050b6adadd3bebc1529ec854dc167a25288f0691323344890f5f90ffc00bb9b2e42d530c6b08c1000e8eb43b2713089093a0a67f12bcef2697f13a9f2b42f93988b4cbd73fe2fa62d663a53ac733afda725e3d238fe7dcd4bc1b1322d1db14d599177050726f4d862fa4ea14817c9d16ac8d715f708d0070c0fef4098e2a7445e2b5a201ff6b6cb404200692dad87ef0928133ea5546d38901963cdefa227c185f6283b5417f9c9f107701e49dcd05ae2d88031b370a43f42dce991c9447220bb7459aed2f7247571cb18b2b3f578d16805f3ef9a0651936b3c3f3bb422bb752fb92a34d6b4d867bebf9486d52b9c0ff2de482352a80849bf86b5deb5cbf8fd8fef43ce6458bea84465705ded3bacaa909d61edef98ff2d3e21f2e442800e461bf4067a4b00f2286053813df7a394b1f4a7ccfd425a78ab9a63d5d3813357ef8b86361417012b85e01a396c5197a9980826f3ecf455d228418a7b647e8a05cf81b2f7fef074738e3cc3362e7279f46cd8d9d927414262ffcb206c71e2c59a5f5c74583a530adfdb10213dbb79a0a18f82552a2242c97ba3cfc926a11a338a50c3b962d2a47ac9d7d2949b693705a8fc88da090192f866c321b315d1a8a4ae35d7674589a06965ed885697699823d886d5e21ea9e212bbb8a7a931203d06ac242b4c2035961b5519d6b1c2c04e6fda70619a45e19d1e8a9520a68aa59cea45c8ff8f947cd92f7367f411578670b5ad259f6604735127c143dd24ecb92233e41811be4b757faeffc004f8645e3431f5b146ecf5fb07ecac9b4582f6001a77a961566d47625a06f4e6296c282936c0e2e35a49e03a4159168ccf93487e5d0418cb4344c2cdc422ec5edb9af78b8c77de31c771c4fc1b25a1bdeff1eb89491310bda5174d8bd34bfe3a8c9e418b3f32474f475c99abeeb001c8210bdc318d4dd1f5cced0a156c6afa1898bff03456ddf3ceaafc5c9df6fdb030b79c41f9d3814e0513d9cca0bf8e251eb86e93ab80485c4adb3707f21deb0a316cb9b87fd06db69196a32a5b3f5e0165a250f982b123600aa9a8f605bda6efa0bf7b1f5aa8bb140d407b5ce7963c444e12d1b7769727e8c447c19186ae7d1928fb2c58d5232dde39de1cdc287bf0af51cc1690667edb39455602c617a9aa23b44a3fccc126c35fd36c1f531de9467b960c09e4d6955faa17912e8922a9fe9b1625082370717cc71ebeb5a623f338a2dc0b0d97caa9fc04d4407ea84622aa47fa1fc4ebe7f0d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf8adc22d1aca811536bf6dcb26d269683187775719d9bc8fd995f00fe82b6112fc2c233481ae996ebf71a5f94f351373df4b75302fb439a6fdda0621250edf7cc34acd3eb2f2e721c59ef260664e7bf09555729a42281e775c55b8354b5d4d24bb81cd840344652e1925f2b86ac4c2dccf5c4b93b542b474136ecc6ce19a621e51d2100e9629e3a88b65200df14ee41d6d56a0e1e91d5bf8c1dee316ae03398c8075386a76eb0d4eb87ef096deb05989212b7dabf11a43f614a349b26b90f2f5ad6ce1077c0f1b40dc52f5554b12ca4ee59805525581115fa9ad99a676c976996a515e0e98bd14bb55eef23256ff7af056ce57625996d09ed29baf4be1aa154d2de2dba6d69edd019d176cc58ba7fdf54b7871edf52a152e04b42703516b9bb3eccaa95cc38a4bec5fb19a030ea515a50e517bf91ca5dcf67a8f80693701d41715950b15fb1f59921686c600c705cad1b115d8fedc5f07980023f5b91e584294b5175e1bd4c5f613d26c7905cbfa865a239a4b129f22a5fcb21d981583f40b6b8ea0805939b1ab8f449b18334fcb69334abfc40aa803a054ff5391b5ecd9dcdb8c4b71d18b631011abd9157272d1bdaf147e845f3f71ce3a96d6c837164596920e2baabeb58f7b41508d4f28a92c6d26078367a8c3bb277c0016f6d1259a5a6e4088c2730b538fda64e055760d5792625554e15f07311ca491fc815fa9022e4cc4c02e85119b3f903f52a7d03213ea00892c81dd5b078938cec58cb960b7cbc22c49aee98196717ae34bb8fe4bc792eda72ddd689b10a2375bcffe1a824d418b9dc1509237fc915910706e48832c8f634df0f18016ca2fff7af5c136667985dc5233ce30c3101df17a841aacc11d22ae01d61404b33b5750ec989e96577124cc4bbf23a7594ed5c59603084217704be4aa6a685022bede83c6f5a8c701cd8e9b530cbadbe7a43d81e38dfc58634a6eda1a3a14e5d5d3eb8e912194c3ecb4caee98a113acf818198c0acc697f51cd1d497a91dabe6b2f43f067b2fbab63b10cb861d1a247fda2c9043931a1612f32e1f7bb91f8dbab8e2a86ad525dbb6558ae42cbdbb418bc962ddd9c7da0712a2172d746883239474292a9a6b04b675fe2d74a88ccd4f799c4d2b1a6b2c9ff96e24ba213a75b279f8b9843e53ea90d6db6d5e4f08036e784ed786714cbf7a6077a431fb1a1abd025b448d94a491d9472cd9ee0b94e9f71ecfffe3facb39de8a0c5dddc3b223cb418f4e16fbed4d628fdb9a9c32204e7be6f29dd6edf35db27f2194e708ef07f0ace929811a5d481f47e860105a6cebb36c54980a70a9085e35191eba7cc8e7f1545e66a3064f6e6f369f14be653029bc897a558d7d71a9f03f771aa84fc06101d68f2cd84e6b7be0a82e5213ebe4d9b6233c45770e377d60da3fcc350a49fe7d0772e935de6effff303d901c11b775366804325ef35f91b419ddaf16656635477e055328e2caaede16a53de9c3d5451c9ab039e60d113c4bb5c1e0cd2fdcf3fe5b76aca6c2b82274d5c236aaaf0af8f8bba4f1baeca35d6de6bbe414e2596faba7fd0b40320ca8195110f03e8a26c6196859aa1dbe7205cb0260008927f9e25b647b4623ac43827a5f8bb3819b918d2270bc977d5713bf4285a3f7c7d93b9b2309bd4db8ce52df03eff51e214d5e5ab665fc821a4ed1fd09a1841ab8538265502758e8e3231f7a7e7cbc7d0a18444cca8ab28e5a1f89ff72da03005d05392bbc925c8fd763cf9ba0cde80361bb8a0fb5e08b6665971b8c298fa3e195f1ce07c3bbba49d3297f3c1a83a66607ce5d54b295a3e6af20192b3c77c1b3ed381e6f0d9fbe51cf9fcb1de475b9fc69ca49bb729e9e5e91254667bada1742a6111e22b859d2738858c7f68e1a095b49cd02e636e6b5be7fe2ba216d2fa99adfad31e645b3355be745dd0cc838c57b8dfbccdf82025875601abf0eca882526b1342a415def537bc22674896a4023edb32eb8e77a5ae211e23e23733976cebddb37e2ae80d359ea3b9312d6e1737831c7eece0f43afaa0efc7ed5330875a6c1a948f5851805e7ffaac59e1a9989e8f74a253fceaa0898cbcb0624bb53cf8c1d5e0967708a47ac130f44afa46809a8591a56296b3748f2a85bbb518feb480e8d4c46fdd4cb6f842967cdc32155e45441c2c50195d11fb88a369b5669f45a59ed4a46398439bafb78dbf2816b38d70619067395581b7253fa766d91b305e0c70563e685d5f0bdb2da6461f6eab88194d09f6e0074ee5d4c910c7bae663d0ed586dd72c20bba993eb26836e804babcb78151621aa42cb0eebf6731082668197f72feacea4a98aeeee6c0bdd04ae8ce6b2abab00fb06088be4e04383e5961d58d75b242dc8642feebbf08dbd14ad2e91a85db6a243cf19b43218e37f233f7bebb50325e991b22815de171246024c1600b7140977f875487eed4e1095d698f580762a99d30ffda9c635dee8b98f149cfe1f387b8c070ecbd7d5441ede91ffdda379e5000475b3d8528339bc4ee0673e4ecd28950d4580e80c26646c355ff5ac1e9f158c849e16f6a1d0866151c73aa349da65d91e54c1c301a8df605dffb082e981dfcfef13a60e16505a5f5a20507f6b38bb33ca13a46c48decbcb29bd288d4ec58e085db207ab988a8c37d957c702a902bea0137e1c590dd6a7679117f7c7df1fceebda12d2782868143d20f8e04f660852016b5ba0802a5de0c8ba877bcc4cd6634287066743d05f9234e9296a8d2dead8cbc83b84b94be1ad5b76b5e97d39fb5463b4bebdeeffbf8c138f55c3b8a0aa999a557f0bec837c9a5d795cbe69455fd0b5f01d54d689f9414463333bb94163d829b8c921682a1fea30a9f7664f09540fd64160c2cf4e26458f4f23f2f98465893d7df84fd1ad5143a8cf6a82cd8b666e34184d9a829eb44e6997c2710cf3adb9ec2fc69e5fa40df20768df9ad10ef80d79db8dec6d48dde015d3e3e66b053cb4c59b544d12f86642f70d5d9bbe0cd7490307180275a98f7448e826f3f8f9d698be859c8ecf406c5575e91027aaf5675b0dbbbd2d129d38324585ee5c02d48cd81b285b4b967f0c6ce503798f9fa78124bdcee841f93a893c407c2e047e81c6f7edca870514fd4eab62a7dcf31fc9d2b23de4db7e8d6d4fd8a8b81b033e1959489e99b8545bedbcbf8ebfef79e8a16e40a4e15df9f2b8db9994822881c95ae4855d6987adacfa2896e8370d29310941ddc8eb3366e1bd0d1e3572a4154fc8af89ca19fff21b99cffbb21a2a10faeac014c0c5624e27412b6e4271c2f5bb009a58db717d4a336c88fd0ada353f7eb71fa9d32b795657dfd81b2d95db3b5fe96c8dc1dece75301d8fb9b3a00324d0c17caa72b7a89b68817a54ae6941d4ed3eafbdbe5cda752378f148a4d57637bb55171fdf1e0faa3d5ceedb7dc50f71179d731879b68529e08bddd80640ace7927391f682a8720d26257a29c90b1a5f2707bfdc8745b7db2224c571ded622169bb3b7ef0739a8ae5c6db7320f08346f73ff9ab1945c1253b45b7cb36ee691709f7664443c75b556072602fd3f19ed654436a0514341402a25c003bad8e0b3b6cc759f2084202cd21f1b76678e37f56d1aad164eac394dc6d0efa54a05603070971768e14aebf746e54ec7dbf32ba7cbaf329335216a7c271d88f435f34f75ed0549f81398dc16d6280de4b2faec00608e010fce97205d4e8d39bed570297c76557d3258347ed3a1e1f01eb2855fc3a197f29499e18b5a6093c5c6f80f80782f0e3565bd4d8a6faa3ae62ae9c449bb2bf93f9e368fc80b453a2a366be10d6c08805b6719756d7bd0a8e5e94c08cf14fce25b0d76c0417123445dafa4d6fcfe2cf7900b2cdd18c58a167ddf08e3c8b7792ed4c769e8197682ad1cd870d70fdcc6a4de025a7535c2f914200333e3decccf5a7fec1b0d9b0f84da8424a675a174a2627146f23883a42e253c9e8d6523a070d30ed18f7e5017fcf55a6858517449c0c4424ffa93c6478363aeeb4930a3668c22eeaf7b2569bbcb2c8f927dfcc3f5020e59fbbece628390f1f499c7795eaaf5d34680567a2caf413f1caba31339eb93af4beda654c0eac30d94a1b62f1814ae25eea0e1d7a0f141c641277bca7dedabb1fce91e5a42de5d230df3eb3b3017ab77d5bf4aacad8fff8da06832dcba14eea2eecf4236703d9c0d06b481570e7a12b4da40b4aef284b6c1e86b01d90d1d9dd6236264b64d709981eb65104e3c6c0337cd5bb9af9aa74f4b5265a0bfe065e9a9ea6356885910cc33808b7cff8362cb32af6b88327b30915e3b352c6176d3f95f12d48a63c9430c1bbeacf95e8bfc6a015df07e8a794e05ffd6d1ce06e8383c3171452c330452f93f398007154bd63d95239016e16aea9ed36f29a208265730f015683fc3d4f8592c7169b43fcbd45f7fd889a434c48408653b2989ea2a5e36e49b64e9a06388617e3432b0aaf3eddd9a07d7cd0034e2ffd060f1e1c22b20066df6f4cc2148d7588818cb564f7138ac8820024f8bf1abb93c1109853ba71a2aa483e135dde954876120a8adb77535e235fa8a1d78ad515bd9bcf4a414915e313a3ba9dd89b23cf3a81989bf49a06adbfaad87c79f2a58f0dc8d5472cf9fbc8094f9d2497b0981581217e7e8a2a2840ab0c9aba4721b8277f859bbc002594b9ad84b2e6f9ea2c6768cbc2bc5d8207c670d8cd983a3142074f637284728c56398b691ca076855ebd49589d0b62f79e6a02dc7f1539669b0b4e6882dcd3a3895e772e337136a23c8aa24994a80b118aa8807eef4b286a8685a6251b389007fe887b2e8e8f589823a98487512f952131faff408b4c6f8911ec7b8ed7a61d482b40157c670c219b4e8b4ea53c109873e13f2672c1e1f653d71ce3cddd785471b01224cda92da4f56b4d2435f95021dd7351046c4db901ea9e2ce10206af966c906effda83b5067e729f3d87665b5256f418af6eecddb386906653a57716de4612146e64d0d6d7ec8a562f0d32d8d08e517e367aeda23b4fa8e97e0b22d4a1fd34c1831a61e0a59bd2c3f528c27a657b3a70f50f875fb8ae8fc69e74b51f587ca6a1332b9639096259b693c963d843d7d7c91ecbf8d4f6d185debd1cd854c0f1a0206540e77d677721341e6243426a3d47018ce10c1eda94c3b7262311dad820b271747f60320a04761f0e472d0c956964abdde619082c7c9f333ccfe1a77f9a0d5b7abf6668288222008b70290bd5f117fab3ebb3a09c39ede0595daf5b9fff4955c7f97dad4bb18537ade4617a93db1b4c5c7adad6f2f6f09be425d2a9aa3c37cac8d45038636dba66a4c47a94d0e1f1f648ffeeb232a28a62c55b7508dc4f91aeb06aa181c7f50f76d449773f67b7e1419a3ec84452c6429e02b3e4efd1eb15d114cd231247422c6aac205ba67435b4c4a943fbaea5b26131a8d43cfdf42816bbcf639a9f01b95fc47a7fd10c96e408d565362c60226f903924819ddcab2adcb2d22c2d6bc8a229d0aa2cb3bc7323856bf1d07bef502b96108e3535eecf314837ab75aec51dd57a5560cbea83451a3b0f1b7350bea7d6db5e2a1cc891621a33c2e0208c6223b6ef0974eac3b7afc672b947b0681d85734e88c98783df632cb4ff29b451e640caba263cb0404a6cc4736fb9b87bda879a2231705894fcea97f02bf8767cbca295e90856cb7aadcbfff4669cb2fe1bc9b3bb2291cbdf701ea728c1df40ddb9edd32b84d94f3c23e2d434845191b9c96f7d1a4b3d64062346d98036d2aa781d53cf9004ca8c5c1a32630b21b10633287cf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h73caaa249ff056afecedb3fdd8e40c42074b30e0ce3a3162c7eb21f336bcd44d873d45905d0abcef57b654b5800f269c58a8afd57d6bfa88d139611da1c7ff045f31e4955759151ba896bc35c6d9a4069109a5fceb1bb1319340a5ccbe5039f6fd2e67843165d8255cc07a4ba2cc5de2d74c8968846ef8dee69ccfdf7b1d3892589d890cb3571356ecbab218aad7d5145922ab0727a6e1cd36335e6ee4eab4351afda07bb0d8c808e5f679b52caf76ffc38216e1ff03bec55c53961f399d31925ec21f43e1275fb51f66b45a54cd1186dfa57f06ff5e0eb78aed1fafaef340b609c74f57678c6481c06f5dd315b8c7d90c9a6d3f3e21bca17e7566c9c27133b78ee80dd13318f00be89fde37d9f080949e1a0c56b481b90266038dc8c3f07a7c45aeda15b5b185058b21e389b02d3e06066f2b7069b36a1c36bca7b0716db3a78a2c0a33aa62c4152cf479376704499016bfb60a83c655fec38a22c9966d314cbddbee0c2ed75a1f7a4043ffcc0a447d85df09760ae7780d2118818a007c4a306b6103625c9e20925d363089f8087b4007f9c3f7835e6eceea5bf1d1c8952523b603ce93a079afb018eb35b0c85358fe9a9fc28e37979322cadd5138485a98aca5412a84ed80a12d1f4175aba0dd37358a25eaacf812cb60737936f8f7ad794379c2430ce9a788b1cf742a4d6c667a30a86510e4b82d1b26db49c7a90f73759d9a40821bec221c230b77b0a39df58afa0a5e34e9b3512ad7ca207dd8cd8998b1bb2e224761f2636155cf943772e3dd39cb1fa36a39a34c4f28fc3b401f100e6c32e97cdfe767cbd2a9cff15b1fe12db3c8c0cadf5afc39168260aa0690de792cae2a95babcf06aead8b1fa80e402e4c1ccd5486defe864bf2d780c66739b661cecbb2e75163009251b91773c09ac14cf8043c818ca736b4b365e18bc4af0ba9e0a09b1beccf02d02675440586ac09d12c92712f07199769e361395f42a5d851a953449d53280bfa9f4f8cad20c3fc6c83cf3a31ff3f09198cc99cfffe6b1cc11e22a846185c547293868ea7f15437ab943d9c012e927eb7c14ba575fd54139c4dfdf2613ebc206a21e264316f22142980e42ca77644dca6b94b32752a02bf5d6206cec31ea1776462dc13cd856d1d282d933492880847aee05b3c01c52046c3dcbf8ed41a2c9245aa878c61779ac7d148c674092814e349da404a771ac1228e9141e132ed3f721ab1eb892b3f29355e7c65c3a29b5e879586c1d7577b38de55d91df1a8178a57dcb16006b6a72cc9a6b6703e45f52b48f58df7fb6794a36926ceb4b3fbec4c03b79ff3e9e3447588615f8c04c2040c3a32b568650774d0fcc60ccc4c3369e1890d66150f83a57ad5335efe00449ec5bd7debb2346b4c22811ec425882818d7c21d4892d1f282157254ca7c97de5fa3ce7b471513ec0b84ec098dbd1604a4fc3b924ba0665888eb9d2c934762c21eacd81b3f0b20ae13d800f2bd134e9934dfb637c4bee073c2c719650bb0eea66072f8a6c41c639125d11c39bf0853e7e6fcd36fc1ab91515dec6387f526b3f792cd1a78ae3b6a4e6873f6e541b802a681b4580246f1fa4efe32ebf5be3f356e18b0663e48f57190326b588fc117bb399fb90ebb65641120a6f5100c52c837662d1c20405a5dd017b486efd026cf20332b4517f87ed5d990b9eb9ff08064247313da0e96e2933350aef2b41389f465178cd2dcfb826e494266bec0e75716860505188a880cd4578d5e0e87fb91260c13d3ce53410bb6bf7a081d718ecfe9974eb17c3c8845bb9df0e85d726d00a7f623cec92dc7a9844af004c2362a823a07e2f4de8f8ae01456bd2fc3824899c3dfdf275575c657c6537abc9af6c6ddb7eaa353b51989d297cc5b110e3775d09ddbf3729fba764fe230c6cf994084492783f847901ef9016d0194ad65317910fcb25fdc831e5cb1a85f5736361a590b4b4b6ad48491bacd4f05cf2c44b86b4839d07ce315fec594e893e6c00df4a4b804b6a3c002ba3ab89e67fc7537eda2312d9010023ae2d014dbc125c0bb74f182df54205fe18e6002576ec2e9d4f14c939958333b82fa001239e76c1ca40987f7688ee77fcd04d4a1f09454636d590394a6be00526cc70df874568ac63fa53fded3563409c3562a1b146ac2249c1706b5a92f7077b791fe777f43adddffa939cd8549303d833b62b8a5dab2e8e2c425796f198dfc0a303a4d147330e1f647578064dbe3e11e268acf969ec270703ceff9e8b0bd1dffd0539828cc9bcac7f3688299a574c98b5fbb1705c6db9aa8eced6e35de70cc7e7f7372363001eb552b678484c599e00a77698d5c2c7d49a6317d614d09eab81427bc0745990f3cde194bd1c66640cd40e8ad3f9bf600bcbb4a20bc5e4940069d7070bc17e53084abfff6b3919407b70faeb88b7211ab5524637641d8d64dbc77554453f59175a23fab15a6818928b34127f7de794af308f056b5b5bee057b7b09401cfdd1ac59547aeb0483b366dfade88e6d6d127e21bc54e2c67e94b4b3c5b5663b639eb4e9807c1ac0c72082ab74e50787fc055adef2d04d0f5c6e83faa70309d222fd8d56190c2705a61ebc1b8fc75211505552dd42360fb485498e02add85f214618a3ea2fdb9f75c1cd22f5dd195ea9d876d42658eec31e7682bdd2da2fe150cd48585be1ac205f415586f80a1836da61d22e584a50da710ca0c403ff9c41a9b2d6689789c25a2d46879b61444000d1bce23ed7b88776c417122a284dfe72e95f48612c0eb8417642da01c8aa239c7b49b378518fa5cef3552f6f79ba0cb7695f8999b0e98d5e0468776c95dd8faac3799cbcdd9a79cb9fea79ff9da432d9e447586b56fb1012a37445b65cc3b0669281dce084e7daa00fa0d99dc00c3c99cba3acf607f8b228eaf417a01d485cda7a67329af3231168352641f91c5dc19213dc8f5ef7e556b639b968f1de6cf6148e27997fa6759a72d3e093f4b42709bff2f3ff410f3a9e8de7ebb99036366c08d914e86c8c4e220d26cbb687e52d175ff319850ef853c07b9e555bd4921bf0280759123df1332b47e69b520f57d19a625cd74aec0d39feef11603e80c946cd8f4d1e24a354ef05936b5c689ddc66001f69176e442d8b6f74d302257a0663f2d9e3c56af40c8d09099ebfa3155d992b32071ce3a82f69eff022ed6cce67bda4bcb918342ae7bbccc50778cc02e5fc5651c962f460a2bdbde0350cfb40f15c33cf9b20d6671b00206b9bcd757ba84f944c838de85edcbdfd8d41b1d9311ba46b125278d8c34f4ea47dc3e61d794c2feafd2d3b4b3c08b02d8cb468a2331e1f76a481943ca2fdbbbd6c8ae599f486ea89d3b931b96430f959f13893b859eb61ffc251e1fc309876702acc892c9924f2e0b3c3215f07bcc447d64387d69ef0c24791b12ac8190bd821a9f65f3153e92eeae1e4fa83107c7feb95ab73a6f82a85b450032ce33b41bb20dfb06788d5143d771fa252c62243990ae9afb01036fbfaf80968c2b2bad6c308d8d38f1ac364b0983a42dac0e8316b0118501255b2b4292d0ff5df409fe48573ef50d476be6cf8ed5abd6423eeb9c8f196bf46a4db349771d0e87310dbc7298c1052d723ca1fa11a85f22b3d71492e88921c0e1aa17eefc71ded338023c3a7789a6bfa7fde5b5dffbfffd1f953e2856f3d21f45853fd3e6567ecfe357523c1751de31d90f32a8cf34663e2e7c26dab0990ceebba582dc47796dbd5b475dec0e2fe18215560538da96c8d2039d167ef9c37623303927af2766492287363a05964a020a8daaa0a4f4d9db0ee618bc6b56caa996b52c9029b8bc80574f95d6aef371ead40d046dfe94b3ab3e2f4a06151158acc7c123ed406b46890c6cb00c5636eb300edf4b879d49975fb43c07416505d24bf3dbcce05b55c41c4579ddc5b63d2d67d722c891167712e7a4070428eb7b324e699570ac9fcf24bd999362a99b1909d241fa393d5fa14cb5dd3776a5b45fda80f3b99b68a77e27ecca091aa4f8bb5b1275677484c910e1c7e3d91db62ffc8f995734649cbbaa61aa7766d5ac02eb2faba1c6404cb16cbf4b97c6333a8997f2464eb25b3026a4b8f4a0007477015586f72b874a1b115f206e3896a196ec2ba16367a17d19203ff34f973f63647504607e4e2f92a1271508232b8c2a0fb73b4999bc994fcbec17963836949358f645a105028577983022af1f5f8f37ec6d758b7626814872fd374df14f17e034a5bdb730d399c946b8342ea5f65480937548e2429378acbb6a78a7dbce9b07e9fcb1ec83cc71ec43d212771dac787c0134fbe1ea4a53c3e83a6f09660fadbd1bfbcea6b06c6601b12d57c77f46f6ffb615c0d3dc6ab4820b37fc5313b0a544a5d92cfbede8e0f80322173ab62d91b0c1bfe62450a836c4c23ae00ef91421bfb277eeb05c1891a30123299ee77faa65089935c677b0b9a0ab3091e271aff4ed13d025153b307c723edf5640fe785aaebfef98761668ae42fb4810f7c05201da41675d57765761c21c0a5facd97aba32a3af0f8bc9d1fb79a9b428885bb23c60a0d3c73088a1ee7fd209b16136b0b3969727ce44557b231e8f02b5a310246291257021904daa8021482971d5b5f9723241939e67c79cb66a7fbf2f67b977f5693e05f3e9d2b748759fc437a08e9d7a39d75ab2ccbf3013582a2372be4053ae10fe8357d685cd8b7afd309c577bf35a4bf09e8c73401b303e24501cf7002a977baea3dab6f04bc9998d219d4df516d29630d4177fc9e7cdad1538f4a00ad2c8e385815622d1214bd1d0523f181639a96a8b5a8c8d2726dc5ac781c13fc75fba1cdc6dfd8ee8c164a1b0337cc4ce2c06ea3253af285ce076f807ba33b8bca4b14797e3ccaf703c727a278936f0ef4d765653565df944fb856477510f1936dcfabcf382782bda52f71439b8239f3d7d829f87bb3d76d02f53c91659a2af60c78ea5a406ef9574bb4b7042e9e47121175739c5728139899f76d4d33ffe4f06c9e397aea11210b76a81ee9dd70c71b69b4ab3bd979830c376dcb20427117f550d7ff88e0c64d74d0518c1251d959c3560ee4d07db781402e70f1f7437be72730aec25195a5c0c0ac04a36252151a47eb05c7e7ae1ab041782f367a7f28de9a1005910e0c14d4cf2b5273fd3713d8630509986b0ffab744f9d5eecc87b9272da8aa03af12422c1e470a447196d6ffc66626ecfc65f9b7345ec4a67c161150aeaac4df861c0122f2af8e0aefc724a151af0f5fb8808404f5787694ae6220b73f6dda9df88c69be76c85594c8bcd7b25ae58f9dd4929e020f5573c8a51c1fc2204fa3295d022af2b01899edf86eccb7b4fef7519e156154fdbfae4839b9fae4847f50fee1eb2b3752128047ef6317b10791b38c425d8282bccdee31235ee207afcf0b137302ba2a10a5a1734923b6102cdc42cb2d2cd68bf461ece11000685a6f66824c8cad119837fba7e1f0c27214f329c70bfd1973262ce6744d2eaa68586e7fdb38dbe47dbf34709e514c67d8746a24f40e1b11f5ae04de623ccf707d71e991f302ac97b3a82efb10aa74add5f391b77a1aca804fa7a4fc6b14a333b7a7ec08e550b7fd71c35927e95ead6f4cb7a208080f7735f137fd5e90feae052f0651135d7553989ddd0cfc6053bccf897793c314f47d736df3d5ac47c99aed0c35b748450908c646137e76bd15d4a0acf63e91d64e7c8b04c8c9fc20b0818a6e192112e2c30fd0c3006cebc133a39e23fae9f4412f79f9be5641c018e59fe703dc69ef4b58f8901afdfb7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he76a9b798a60f0c2e2de1b895f7f3df2576bb620e04015a2a5b4dcb84f20997024e2dad832b00df122798d2f8e902cf32a4b1174a675384e73dc02a0ffb4e72601451a825169babece70b022673e518fb54de9e505f2edee2305b367738456e96c935b20ff8eaf1ef9ffed1342ce2c53a864ba4f4baafa0281e5d3a89b7c98762ac350225f5504b6eaa37b52e44920f6ad9c4868a461fffa68b66ca336ff1724755108629103b0fc07c2ca4d1dd928db820472a4b559649a986a60487dc551b20c39fa190354caacd2f3d494cf2c935d550fb0cc594c877f840d7a87263a897f37c566b38a9c61bf1e686fea8a1ec62f8fc03a92af29247d219b7b8c5593b9171de36caaf59e0dd886a2ad351c4ad4af65859c52d193c6f4deafb9ea42d4256365aa78012807d8f23d9528178de968d49aa7f6b4197552d812e2261c5446f6023afddb5b746f817ef84691d81a8a249d11df78d988cbf64c4bd3dabc7fbf71234817d602e15210aeaaa2242748d6dce6135dfe1b95565f334b32d2a99b6899a6315b23e41bb6785bdcda1c740ee05c17d0ab10871e70f33ebe5c4a2df98c3282e262efa101c144cca2a5731ebe9f861cfa84493a5af2e0c1e31aaea43c3897c067bdc1cc309170d362d0ff34932b400d0ad19158bb7fd1d50fb20182acf11e12a5c01a0568fcfbe6920ce1b0906f165ac153a4b0bf08e8348ab57f95cfb46a516107ea65e405dd6c07df3a49e2706d7ed9e18cb1d2e20e5d8270db062ea45f8a146d3aa7922935f6f63d63e40b3140696e16670cfd03a75b3ed0b377cd0eabffc5b1203ae68c3289b9aa974de0a6da0212cb6cc46a0524b86f913ef79f76fe23978607fb4dcb12a780732f4fa6a816bf3f68d9d62d6143dba4a82cdb8635ef85570baff50e7b1cac735e456a1a1abbdf357df14c9d89e16a3f4b0ef53ea79d8d9f68946be97678a5c7a28abd20ace6ab093c873db8946eaa7a734162508d8db4b622427ccce2c3c1ac22590f02377fe8e9f2ddc02d881d13478b595ccb58398f6fffd9ca6f9eb37e9441316f654b18237c8096b7c2b43857cb66147ffdfe5d06d1466a9fbe075340509a28996aca1e6acdb3f0e84fe9f283051c0b5d888ac7b7976e896f8d3056bf1865b1e506b0a9a7d372e133072a27799da44712fe223fa64ced63d82d3e6415b2999bf54e8cf6e4e3e5c5f11e7e52ad288944cbef52c615b60a5f1f4648e0e1cb815b63b5c33fba2f5393a3efaa3e02aa86a233e47a1551e87368b15269c524722dd097270712799eaf7157db886b6fd2b83fcbf1885f7a747da7d3ea9f3ed957f0a645446aeb329e68509c3176da963bf18e0fc2263a8ae50336b88fcfd4806f5fcd32a543dea5d4702c56ac1a38afdbc7bdda942d54917a5ba7a853730d4e3f199430305be93310b3c62565f97a2bc115e69f4ec30b9e3d3f14d75ec48b58022150b014a1001b87096713574d7a929fedf74288b02001e8dc02fa5697b72696da92d85ddbae1ac24a6cebf21afe6b2f58cdd6de852b2c5fc272a428e56aa8ba578457fe4c4572a569267c0ebfb2fe098cebbc221d379331574d953affe19fa7ca93cff7a3418da6b96b5e99f3a4ad2b08ee51c8d55e9f564a9f3b980afeeffcc9a082254ad91f61c6cd0cf085a5d72c3f08dab1a2acb594a66bdd74a92ece695a9a16ab9037f29da139077c768476566a94765fd8bd3f024c6b18c19f1362d514ff5a77df0ea36a87695c85005f4b20500706a78e9c38e14005bc1583eaf623398960c5e96257a7559dab22c262c5fa59836a5562cbd1e2f80596ac9176b0ff4cfc5172510236a730dad85d7789524a93b540c4a9b0c5889891b5c3ddfa942e7da50d110b3fe85a97adfb6d21aaab1d786aa8d2b7e6f658e3904ff50c46eba9ed42d5db5dc08ad930d95bd22eebde35431d2aeb6c1947fb8217d6bde9e41e66ca75e27fb7dd0d7128b6857d728524bfc49f4990e5e0e060cd835d1a8a8b41ecba955c8d2f598bd8efa967a058c66f90c4866e00ba90911b6b3df37398b1833b3255ac3ed6b42e766ae5025ee338dd9b50f9c1a1f1c1a0d9714d6cdb2534a26391620023cbbe977ebd6c42481e8b78c85fa817179000ffeb334103dc00b60b21769648d361411099218cb89ab4617c813a88ed8c11d82cfc1cc74f4113e6de41b7ddc89c04f881cb6ef1e7c1895516df89a1e2bcff4ce32eaf05592b2d5f904318f3b0be4451aef44ecde6c5fa8069737ba4fda511588413969d9a0668e1fd48fb950cf27a21d748c2dae6c96477fc2ec33b44487fc21b67702404f3e94df09d9f15ccbb12d79e4879d54253192d35f78243883941b5b2cc020b7a51ec2dca87c30999673156fe22beec54ea0a6bdcef8a5314cef6a20cce301a273a6f8c8028df26c8621783c47d44487046686b86ec43b98bf0bea112f0c83d1639cdd4cd079c614c562154c493fe4c98cfcc53965c963d6f0722e2535af13bbae812e4ce60533d6cc71f2ffff5d8bed5e231fb47c522cb5151c536f847b8ce420e80569c52f3abe1944a98f4de37c9de16e21456d4a1707670d07c5a3914cb34dd7c38e0870695b4f3b2d548dd53a15eee7db95ca43fe4a0e0b2193e0885da3eba77c3dfae75b1ffb55f038e13986aa75703c64e2ffa88888a8112dee47080decc28288af6771fd6ba190795efa7b1d9822736bb50a8fc30e007e4d0fbf3cb15cd59b4971fce2802a35f682e54c7253d1d5845c61f06e6ba8dd0ab5920dc3377644cd669539d68874a7841b4778906a925db5500afc54b2bd13ba5841893967cd39dd5540fe32a54ad4cc08156b41427e6d902ca27fc4bc6467702eccfd382e6e0a347976e4c5c4c8393150b38365eff02e7a0e7bd5f9fce3aa50725c91b77613f93e153bd61e901d2f84c5816ac8fd2af1d4e8168c56be7e0934bb43983409190ffd9f041201d0e00a96960f001fe0db31493e6b88cc5a90ca4e07a9decf2951b73c8bf49151ed6eca29e048c43ecd6c3ac9c4f644c0e6f394d07827bd542be8d201e00845d636ac73da9ae2575eca39f7ce24e83a5471daf63c04588ee8baac8beef0e86d2009497fe7d7157a2c84f29ee1e2ae1249e43816a7ecbcd6d490770b52a497b9d6513339837096dfdffae2ba90ed039256c1b2ccfc268b9620e6596e46600070c64d180a2497a964d058955cfbbcef0f0fda22b864b2973b1f5a1d85fab25e39bd5d71a52bdfcc4c7face8979247593ce976187060ee6f57cfee43fbfcad2d61832d9adf93cca477404bd23c6cf8ef9b5e64fc8784d9d9e1d3c4ae35a5fa873009789b20db8d16a055012222fafc90ed1922b961f3f498b5694ec16de2324878cb3b493574fea7145b285df662a84e632d758ecd1f34f9d947548c0490081d5907acea17ab47bcef9414ff5d09e2ca1d3566335a0f7fef7a8b4865361cc271414b0a54eb056635125b93913dd129fed7dcd9a30681d4036efc6e7a6d7976a4bf70fcab5a6abb4fc808cdf98e7a8a91afdad47f075d5aacf6efb846bedb78e1ca20d398d72230ab67179e12e5ea0536510eac72d2c90db085a35a0b810f2f0af70f706cded12235f91e3a1f507cf880f3b5600cbdca9a852aeb2651517b66b3b8a0027d0a976f306ad6161ee3a2c74e73560b0f965d51b83dd168d66e1c0ca037e8db844b41aced04ba2739b2ac0ba3b5fc2f5625086576f596120783678fabd8564db659d9a30d1362081878b0079610851bb54c87495a3f49be54fe0515862ffe2e57c1a2a5690a986886fa815ede776134d0af9f75280561239cea30bc8433b284ff35c71732b8c20a98f6689035d8caa7add5aba99bfb1a7ae8a20b5582f55d3b0d3421740582a65a43726bb55495636d36d4a147f632072de1ac4c767df109c864c54f2c9bba85531e64e004b80dcba086a6b78f2830521787e989d87bbf29bea7bde3bde28187e9b018d41b32ed8512f7ae640ca731e386585cf40f7310cff9881d4208cbf920dd3dfdaa2cb122bb84ea4a72dfcfffce5e4f34d6cb59b47081dcb3dd8d7ca56f60958935cc6b1c54c1f3c247d291a5bbfd254e3b6a276092614a9844177cd540c377c5c7ab66751ae3240c2b984ef3c45993569897380e002309303afc116fb8cb9ede049ff147ce64dd45d7079a243ef5053fb57c67638cdf4f4ec4e499404d26ac05ecb102838c273810fd269921dc3398576544ad48b49d0d5574f3cec25792a9416bc21936701453651fc5c27344e2e593e9dd25391c29e36d42b59d01eff9f585ac0e86a0da4169746ed0d85e712b1ce75b89275d79694e0bca017034b6d84b293f9f47a03823025e4978dac67fa84c714297587fb19bbcf4e0009cf3a4a22ccac000875caf925d53f2bf84535e607f78c2ee7be73b2f069d6603d1cb24ea9332e620e8d7f6e97905fbf6a3021be957ce14cb9e62dd52aac683c97a7a4210e9cd4f7cde7ebea4da11339d9c27abe1623553d429978a818047d5a7b22f2284f4528146b8adf5dee1a4cdae9f7fee6201f4da98453cbf9421e32d07d93eb39bb960385fb5ffc969afb34a3924c8dee3b4a3fa2055a8d1282f872ab77e9bbb87d48c2bf1e752a996a19b2dd150d6d092f5333cd1d870db00d590a0328ed561be2b390def5c0b5c8f9dba14b11adcabcd65fa80fb8b296e985ac7d0ba8e4c5060c7f632bd3579cd5ed00d12bf89daff38344ed8d57e21a4c8f53583a719a8985587112fc902168e33b6b698183bdf779ce7f1d03576fc6fa448eb4cf42cc65c71013b076a3ffb668da94c93025984410cbb399658334ad31f4a2c8d7179725ec315875a63b136220119225894ad37e03246d936002fe4c531ccf57ecee9c05893b834fa9a28b67e39aec18d8c5281a69713d72ee0ba5c4c3f63a826c495f3ba8999bf64fb85e64e1baf2eed6f284bba4eb9a39fd87078bc38f1970e3ec441d84fe4d562ae2b4f0198260504f5713145f9d6d59f59492c0c733705c1afc3ef6263ee39444634f5545dd445dc6ca3811b594eb6ff4eb3f986d992265a07e6e928f4f5fcb0806dedf9f678c4bbc1e16eb3f1e4c438a6ce70c90f29faacc44e75afa50c7bc1e3caebbf22b1a3245d2f1b591c9b2c8fb74d556373f389383cfea87474dac261f4142db36d1708b33bc690c2feaf67c59603f46347507f44634457c5fc36cabfd9f669f19916e938d4a1b1aef86cd8dcdb6d2b62286b923ecb1ed47c4483cb89bb1a1f13ec8d45b8bd9b0a8d5bf0e3d96ea2e8948e1bbe8f2a2f27d5b0c613945e935662387cb13705f6ba06638bca77f44187036ae2bbad6a990ee2061ea85c189193eb30e0ddd09a934a5be4f1c24983d5560af9ae851609f6b9301c328aaca39ad60277dd2aa3fc0b966c1bc43c5eda188b70ace1610608ef889c79ef4d2aa2b7278d81f57776a161827607e9164586ce91b75d34cc7150e76b10a8f7a714c0c1827b253f0af421655c20f46bb2f622e40d080d08255c34583ced0f4b142c6db610e7eddf363ff6c082f308c5ef32fb5825787d08f26da6483ef7b1229f921bd1266c175997783ab7d0d222e225dd2d3c93e6647cec9a51eb03746b5e23f49837454e18249c2b9ef5b3b7431de06c1f31495e654551c93782c47cf34b39f6ac1a8908ec7dcf912ead58d28977343cc59621d372ac9e793277a16d96d159abdde73a56aeafeff47b17b3243189abebba727f5f964e1e89d24ecb54ffcf9b55741514de11750cdaf6d6ac814e9d52f6f94f112b758167475982514b3d50c3a7b23e661fc296fe2e338;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hedc8c7eefc0a1453eac10e6a42aa47642fde4a974bf69cadb5c127a1215724f1fda31cb16803bb857ab88793f4ec5983875fa215b0d6a02ca025f835fcde0fcaefa6678e4818cc3d987b8eb4fa9044665095e51478659851ffac5954d5732d0fc8ab89f03e3c3a61d28af9d6128af96ad2a2fbc36fecd3cc8cfee5d2539f7fa02d26da7dd52ad0e547a2c74c2842ea23e81341acfb3b1be5d48b1120694c744602b2c2589d28fa13d8b26bc92074d588562c2dc71e719f0faae94ec7871512f71edde51e6a7e86d6fa0c6f4095d50e6d2846f9104007c53418d3a32cccfebd9810d52e1cbb3d6494dbe0458578cbcd225c2cb96e6e9d583492d4d7357660ec3e511ea13d61686ff5bde947bab76af4880280f0a80b89a9959eb298201c3b2eedcda797fcad5c117130f9174c20521eebef5918249c9928e77f75ace4f1bf5d1e7e68a4409d9893f9f287b0508820a24ce2b2da0c198427836193c966dcfc2b67fdf7333ed7390d64a711fa25f3e86c52c1f21c936fd27b3a867710c17186ad4a56c0ca82545ba15a4ab482990c74b5c3cadd8922954a7b9cf8cf922d8efacf8758b043db71d35b7b740da3d8f38c827f8bbdf27371a00b635dc601b7be355c4d6c9e4c24b7b0d6b1aa948f10c1a374307e7ef83a561620329d169ca8ddacb7431490d92f72ff19700389d7f855c8c3901adde74e21e33363665b58f50fa34dcb5abfa56b05caf663085e48e1454f3401cb878b6c50a564f34cce9797a81984cdbfee77606dad7aae5728d58e23a63a8d9cf5929f49f811e43ff12b213f9447f016fb32eac7cf3f7527094d647712f157b361ade0904f9c5d23e5a44e85ee5b21cdb3a09afe033f123a4dbb8735b733bc028309963fb8565671682ae88538a4dcf52ed241cc2a09fcc0a06cab327f3f7fa503d4399d2357c35da9a87265ab15ed2e71a6703f74a69fec7f392908fd1f5a013bb1190745ea79bb405e353c2c6bc437a4d7b2c1b6b3c6dba8b6a524d087a5f2e1f0b19737d9b59d1f2b5305911acb9f2835b1a19f826efc9aa52ea4957f192fab030ab57c978dd6384fdd5af8533cd5bcd6d45a990dcc79c51a5c96d02782c7873598ad8f399a561a1c2fad7d3f45d53a23a316b4d96999f75e96f373e3bad05e5de880ab78e24820f4cd3c3d37bea167c704e57aa113a7958d59dfdfbe1f39294cbfc599391c79940eb578b506233d38881bd6cd8608ca2d09a6b4314e24bb7fe0c91c54cb8109af3fca9f4d99b93ae8c0d52dc95677666fb8c8444b5f28d74976805ecdbcf416b2eea57c14b879ea6fd5cbe7e61a80b0d3aeabf95d02412c0156b9a1943f17864d07613744d68904a734d33e97aee230ecec8dd912791d064b971ff5bed901f36919408e5d0e6a786fab0223cbd9fe8bcd9b02c588e8a99338c55c5f00bc077f6ed6269e7bf0f2ddfb4057355935e19ded458b171ee0ed9945a431480ee903936d5e7437c7362d0283bed804f82184f12977b69a318e5f11d62e19a7650bd6699c5ee85b14f5f8d1bd0665a45dc055929c74d94e54e5b6e9c3b899648be7ecc4927d494c2c5cb5617d0915d2db5414fb1fed0fe1ca450b0e2ee8c422dbf7be0c51574ac40cefd99bc7d47470693bb45dce672961810a65e995c4057e9a59d9b93400543957db8a72a21dcbc4a1410d3b154f0797960466c4c597a7ea3523a1e71a50ba182b347c62208a2c0196e0ad48bcd1f60fa7c7783ee714a18e54589499ba11ccf408f024803e1c45c69b2ce90e3498569e1538b0f544ac9ac9b5987e87435be092124d5dddb27c390e3c100dc41af1662f6a76defc765666a8c08d79e434ac88a54fe3ef3921907dc05637ee263134f3a00f008f36cddbf12ff681bf4a2afc28909b22dc4c6c06de88c820b0475fe646bc9a16eb4c3cbaa96e5e29a918eaf90bc74a8c413c6d6fe14d10734103d18386489a3451f4ed64dedd60123417183745d07f0c6b25935bf08079b1fde630726ed5f28517e9bccc7cb2d68c924ea52033c9ab1a966291de5774b458400c7ee07093f888862f0e443befc1a0d0e9c74772dd054ef975bb30a45ac307e5019cc74de72f6e87e22911a0e3f79400f391f79755cb1f13fee180bf3dcf2507ebfb8ccdd6f66b21138f1c29ea5061c769258584940c71808a9e9b79b554038299bfa20fdfc563fff92d64eb19298a1695b5845931560ff81caef104982b5c293a79f6e8e1992b39299421b7257d7ad4638163ff812ac61e4923b48f37d53c8b391b33e0acc9fc5b6e52b7d9ab01f0e5085507a3859f877deac54532ae7620470ad6c2b254917dd0a9c0d038fc68642643804c5273fe0a624556b1c5c53c4eeb33fa2de34616d919c1f64d627f9f3fccf2d6f4af3092aa4e7101053ef0b6e430f334376d88b80a548b1b5b15b90ad69f9c79372d99096842e60c32447c4588b684eabd30f0da7513bae7d16f6662a84b3adc22b02f3d7abf6210e94fe57a9af4d8500b196932ec714a3dedf02a2ead68f37e71bbe00a9029ada618ac4690bdc32e5ac47f290acce1c1588e68e68432bb4f3680c660d2be34a5eec4e0fc167f5d4fb5c3de1e04b0bfbf616cb576b1bd6704d42f93c8f8b571df01a1ae3c646216761e787bd0a4f294570541727e68a15195dabd84b8c6ff1bf6604b41324ea02bf7d57518e850ae842ed630669f16440c59f03bd4022bd4a8fec18d2613df9b1ea813a6e12c0ad0455d55736a82bb2fa2f17ed124d23282b50a29eaa00e5d60b3e8af83112fd8b0baf6f13b9ad9788a497c681cfbc49490393264e926517f80af7c997648176471a869cf192e7b0e1862d4fd3d6ee4bdc17b84ad3f6970532fe14340bd99aca3c9598a8eaca268001af3d9e512061ccf9c9799b6d343a2ec87028311c2c335b1f470ac9234693a53e2d49f1924fedc1cfb6b12066de4ebf91036b8d92712f92458ff8d621f675ceb66ed7773b88098f4dffa3d8f7a94117b34db2e299d735b2d7226d542cff3911da0293473138f83227268bcdc7645dbeeda99871b2afcb1176e09b19eca942cf7f8a069be7b5e534f2ad40ab75a862fb342d01b14cde75e1528d6c4d7ab63402cfb3fcf372cd36963fa511630b59f3d9177fecb38858159a36bf47fa9113a88121f09c3283076ce91730f3b61835f20301826908c7c4ec118acc4666c0dac79aff7e00d09ff3d39cfdde6ab166fff10fbb28a3a50e0dfcd703e0b00629ee92a70b37211d746296e7968bb5e6a20acfbf47c4d6676b5583d3947c17fb17e97d38f97f1ba9b186dacc82ed5cfc41802ee4572bb35e7d3220f39777678686010824b0293327e485f210d80f33b92f3d06304f98a61abd1c7d1816e009ade5eb80b0e2118aeff2ab1ef8fd3d999a2e9fedf5dbb20315506899bc4f1545b4718449bd40f0866fff610651873f659c441c4dbe5662588958662b66d71920f763b9bf57806021b321560efed3372c653e6fd30f6282277ffb5f8273a84b761d653c6bdc74c4495fbe4b28325e70432833cb5f0267920bd2076542fbddf56c8a593bbcf62c80960049ce51ac111bc942de5f2d5d3e2eacd1cfd523ccf479554510553ce9a2a50cbbb5978526608e5d21374fbb23916942c4d8eb04bc9636afae4899a266955fc50b8967951a641ca46e6a2d318f2f85aad7cf2b46f20a84756a2128763c2dd57bb816d1c6dad0ac59464a187f57cc696a753846dbb4fbda98c44a5a4e919e8251d62250b5f03039dcd496c38adc43ea5ac68603d4ee154db35d222d45414d768802eae9353afd46d5e6e8a5a7e00ab08e58d651b5d2f55b409c8121e5fac458cb3ff1eb37f8d825049b023579d04ad3942c8373d0beed804538764cdd986d72e39a696030dc5b60e99821ded8a1c4478cb471747f31824e975803ada9908f3820cac72e81e651fb52e7782fd18313b2291d1bb613eb4aca588109a5cc4e184c9bbcca0b0b16419cfc6596d98a024547bda03bb4c4af5ac23ef8bcba12a7e38162c47079656d641d80ffcd32ea46a287f8ccd8d91acd693d8617e5469f20fc02c3e8626b67a276864a87a406390f7d0d4392e93fdadc860a1f8bea74bfc746ac441c5f07c0163623c58069e882ea9180a665283698b1bec8bbe31830316186d8f9ab69c9de1c54cfee02185ed98a8612f473f8e1d692a9c2607c901fa50a6286b32133323869ece4c3b2e9c1e27f19f10451538060b6edb5325f9b2f2be150e0478b2542f9ae36974f7be3d6ad9f1b25fe76bbf5970c9cfd09a3680cc588ebf2321ca333a6d2cf29e68beff55cec2e578da044b4f0c0ce224fd155077b00ccf13938b811d6fc4c3c1a7a4ceb1621313326a32b54c292ea66b33c4cb633f934162bf543d143ec1ffe5630470f06a8d05ac91497eeb14da8f5ce76f9b17faf8ef74ff4cceb6c8b744a4ce7ca1b2298df0dd9562b362739f31ce6ef8d5e5c23862eb050199a288c00f45e726cffa0ae8d8c0dbc28004d2537a00d546440ebdf4b74b53152c04147b4e691cbeba62dd0ce916b12efa972fa92f5ef29c234284d8e4aa45d30ea5ab7bb752ef7e5a5d81a5920126d3f5bb69d5bc1d7df10a6a018e780cd90987ee4001865d5b2a2b202dd241f962e6c7f2a289ff05308e182d33191f2f409895d306f26f13dd4e8defefa90907ba81618b1cf350d1b9d0036afe4fdc44ddb226090ce4545bb1379be97dd3bdb9485a51db9a9840ac5014b5f58c045ce6ad7ce2d8189fefe477b44465945dd60a8d5154dff9124bbf1d1128e6e27dd913f49cdda0493fa8453b6a103e4e2b8e99ef7f30bd451189e0bf4e7aea15f982dc15f820615488cf7fb6999e1ca4e43d10021295659fe16095f2672620db8ed898d6d1e8fcf2427a0d01b67817efd07e0eaabccd6b5bccbabd122f12e5a80d1ac6f9d38747a575005cb885a09f1c4ce870c3a0583d7152c73494e5a50940d1cf8efaebe33a45d9232b08103314f4737df7a2e78a0843e1c259b8f7417a07ee39edddc3d0bcd3e20e11272adc73e049bc4562261ffe04d567d56b47253023be30020d6ea76fefdf2f12746c31b74859873a2382e596aa40e66b0ed629be9e0d23a013ccd10e6c4346e7b05dd251fa564071e2abebb53f9be6a2de3f6251c7c9a53c1f754474f4c750100df37228df3115f80fec9881507e7886f2b51b8a82a91b9a1260a5fc390ff3fa3f2bee6cb9bbbc574de62255eda654cbaa69cb3f510ede304daf5175ad546dd47826c1df3363d324c6bb872b307144fe0655d5e1fe4e2b004598e6cc5464eb9415674aa06b53ebcad272c81523c8fcf81479d96ec96b3f5195a31b1fb1dfa5e9f8d7fd9da04c2e3ace738ebb08ce01c4ecea4f0ff9a17fd7ce18bbe14be9fca83d60b68fdce3264ecf9930144c6157ca0caa4d21a20d5d9338f8a010fbcc8c6ee97b4527c21d7521a16111bd35044aa618e4e8313fb29d6788385d3f6182eabb6e91164cac7ec6a65e3074da5d5882573d0a7177069d315375d7059666dab60107ed784a82e862c89d60e98afe7e4be53665cab09da0628965c8b42f0aafadbc6a5a8fd9b892a56a23c6021315f8a07c2b75b5e6286819990f1a91ff99b900a8a004a0b53526d6b802b6ee29150d97633014215297cc2a7acdf00b878a38514b4da43b2a9855d38930a1ddcfd9b7cb8aa699b179a15527f6ea431b18fbb6c5d14c774c2ce0a77e5167e834beffeb513a409374dca81d8bd0617de58ac6edf6858c2db3387cefeabd7b07a8e7992e06e7cae22f84bf6861b6667d2f0ffaa5c346;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd5ef89ae006836975d434ad50b3338d8db8698e6c953ce4678e6d6ecb91d0768599aaf6901a3ec341b593b298c8bbcb9e9ff07288aa42e47b65ab498439584c43ff0b942df911d5407c22d2a57e6561a54d9452ea1f7eba668d701f2adce946d511761298261f44933a3236370606af2ce4addb10705c9e5b9959a8ddf6ed21062cb5842a6a6d08119e1b3aa5f0c2c51f747da40018f9d85947a0c9505d06ab91a8de6b53ef686a7ba01111e256d7b874a8534d40640824722a8028b5cd41b572f90d12424c32362ef008abd27cd85a04f6c7d75fbaa0a138f166ae34127603b4672891dbc213f179c4789b7f18e7aa44721c783da08db23898a8a33a51164d58caa849fb75ceaf7df745bbf49735d91b4d4567baa384a091f44ab0a6a0154664cc2daa5d0b38d9ea32a1336b9613fd331f3d2ed5d73d82a661a40bc323588a84d14b65938a4f30d0e117b43cfcd572523ca3c393dee49e56a51b49fad9faec36ff1e11d41f84e4e30c287ee1f3656c712164ff755ed076f1b2c23e464a2cf5c1978403aa859723bbd4274d17be24f69c70da3ace566c96515a5244136dc5a945f3d7b304c4065aaaf4cf26160f1773af717b1beb9e80290417a53ebe82d497cf0b7c867dd4e82b1eb201139cbf14a61b7a7d4285934785949af690e661d2816783d9541c18b9049ed926bf0db2b10a2b83e92ca4b3e9e9464c05d94d4e430607da138b3afe9ea379fc34c14e48d8d2361b264a4eca12712dc4df8aac2a71b15213cbd995325fd30fbb81b7ea3ff10e7b71367d866ac266851092feba96850cc292547094914a6b5cb289e7f29bebbf017a466726f10f73f8bbc7ca5aa1698bd18ea82f454a2be114860a888acabad07d1ea36effe239d2bbfd1c285594090ea0ddcea63e050cffb3f58f20350ce61a4c9cec9b05b8679552f6450ebc9f36bc93ad60706a473ab4015debd28d40413f4a4b8fc7d0ebf6e65035c176ca0c21d0e93a4c5004a4a079643fdd9cd95a5d8e7ea95223d4b919bcce67e24a91abb437378e6529f110c801065595d8d4bb7dbe7e7a0681039eacec906e038a4ab3ba6df18a2717005ffc736ccd3f8511d11fc1b61f864718a80600bf2383399b81554df5f3168fba8f40c6e034fa4e70ab3146e2bf066dd08c3c51d8511dd586d77a9dbfd79c8768fe5bc7fdd81bf1d07f005b6993139aa350a1f4da91409995b94a7386795f1bd6d038bfedf38c828b9d3810763315fe7c98588d85b5fd63087a8417c4c490d329248890e147b90eea9f583ef068793f81d94b4421546c091c041bc1eac9725ee9fa4198897bdf3c5de63d8d57d767742f0fbccd3cc1c8a973a4bccaca2f7c94443e749d16e3023ad4861fc43a76c0ee32f1b812a2d0c54671ee4b9f61a659dd9192523a48218a2aad84a7c0070f371ef040bc67d9cd2e9304b76eb521eafa9b60292ce5d4fb43d08f5ae8145eee2e00819b46896c0ab04e8f5144e07a6c9ade9681154d39fe96367c1a3638bfe88e8815f4347bcbbbf6571f8c537f66e4219401154ac8f7eef2cdcb17351e0d57fb53d96926f63c1dd812616a50afa1ec0b4b4eed310be288fee8d78a98bcf242686a2643ef7e63476a9a1526af6ce84c5e4b7e7c7e9eb4172a7585605a11228fad68888d5e085e7c69752192fdfdd6c8facb70ac27bcf55e51fe7ab6444b8a8fd0581658cf0feb93a6b1eb4f024d1ef1813ee5fc7cfe40cede1c68670c1e6f8cbdf7a527843dd193f8970b6fa5195d6f635eb68d79f3ac929e3c20ab54d53f71183d819b055c0ac48468f88da67d29f43dc757637fda161c31ebbbca7e7b09c5a152513d6040c7f11c7bae3271aec9537a09c86b3efd50e5e928f1516d8c531dd582906c8884b0ee3567f55f43468e5d521819bd89311fa4ce1ac45d76e94ee0208d686595ce7a072be556688391b93793b2dd967d29111d880d6ff0ef1c705016d1f510d54d5d5781d3d2ce47991b663d4cc928e67a968125145b52959e1f944903a48be5962292dc371ed9dee4cddf584f38eed71545d32a5fe085bc4c632c8599266b42c1b58bf46672714f40825ed57acb3ae4a25ae5945b0681721968b36d1a9c12995a92695635e686b728994e2752954be877977a0bb2f001d87d2c053eeb2c3caaad0e49cdac507b51e1814eaaa0822b67a31a269ad12b0be4da00f1db3db12418e658d43c15939f7407a0f0a615a8b1a736a7eeeaab5a6f59f52e373ffc74ad69f7917d75b7c68207473a6af2bdb136eaaab8ef979a6975c2c0e0ca33394bc0257bfab8f5a5516c2b57043ac788991e679e36103dede3722de0228888e475b3b82475892ce7e0dd03bcd457ae0dd490dad1f2e405eda2cb183335051bd0db2fe3bf5b356755e7e4e4108a7d4b95033902e8d7e4683fef1194d4d8b71d3f56287f8f7caab0eda2ed0b896604b146746c2b888cdf50dc562d092f9d1911b8a49a098b74ae7115d30704e7eecae4cfb54ef2e7c87a0d3a22f05178b03b0462a56bec1f5d5636758d4ec0f1c434b6b44645e3b5bedf9f9d5bebdde7dfa52e3229e4185d80b07771faf5c8508a5c947a6e5a07dad3d33ee6d36d6557fa815686a05d9d9eeecb281d4d0d8a5fab4b93230a556a60597d092b4e622ad5624b80aebf3cc021a28a670afd3a077916c30204b6ab708d49d2e58063d2455d209a146bf906a8254fcd9d0e92845b3d1002f704948004e9c0cd3caf3f673da989d5fe861c927cf3c8d78ff5917f04652c39db7efbab866dfc883e913e159463251317facce000e5bd41d0ec2d7cb380b1dcdbb709dfeaf5a7504bf890b903d71d5aa0121017f1e1aab442fa4702c612b1db80437f2949c8735876b8decb9fd8e2b8fd34a95ad1d64550ce80c12839376c6fbc11753541dbf43416ef97c7d216cc8303ce75581ce3f05ccb196b01290cce4569605a8adccde550717e86d9b8ba165f3f0a51bb164509c573aec5f91659776c742c208e1a8e5fb6dc33dde6c9d02d4dba19131bd300f1b6125132655213e8bdb26755edd61db42c61ad6c913969605d10309e73b914f3697efe507510b03756586037328f7a2aba5cff68681b29ec7884a7ff8fffb1e12d18c12a5d014377e9b7dab0429ed3b1f3b6f7ca87eb235bec0711f4cc369317cb950472f57cb72a462af20fd0bf0d4ce324bbbf8fd056f42a4fc01a90c533dfb2d63a1264d201adb1be3796d351b73da8a02c957634b15ee74ec2686d11b939a01a2d7571728ff44aa98fffb5b0bf306afac19bd6a41d1ba3da735787cbddc9cc723fff5fbfb0489f35cebdc76879e4cbb9d78ede3d858d70c6ff6f559e9cadb465fb03c1df693d8f2bc2eed27862e1f1a5af5ed632e5b0f4e6f1adee9645122a9eec250cb1f9e388ab43c8c18976316cb832baeb22ff0315ce6f26dd9649a2ef698b37d97eb57a20c051319388af6bc19762dcc2a2166c0aec848d45bfa41f450a3333bd24249e4b28ad6b348b006fd7e3110bc1fce0d7eb929751d2e0958da5752478c37c9852c242b806b30dea44a58c41b5dbc2a464b70d64fd72ca8a7380d3819ddf053ea4eab933ed3760fc5ff5a0afaa00376c0cae0f08c612f012f127625bdcccdeaed2e0261ba99dc5a14996fa6f2e50dc4dbc0d4e833e9fb170dd4893f4f91ab1bbf356b374f72f1b54af6fe5d4deb9df5a0e70d7c8cb90e4a6d27ddffb80f3f5b53b2778885038556ab374dc37d175a4d4c502d17651be8a96d4603260285c747ac03e8bda4f52152ab0aaeb0247965f136d304b6c180262ccc5c0e58304adbd57a8b5bcea7fec030c8b45e6622214ec292bd0ba98cf8de635db6ae6d2874ec16ce019c3e33a0f0e8bd03d83c0ce1dbc05e4481505ebcd35fb04b3746d3af4d54bab9bdb8740fb5776ef47a66f2807cfda3322372a5beae6cff8d93e2a53e95096bf0df5036b31f9935d6497517f72feb3fc3eb1772f39896bc2c4f678caadfb951bac3cf5ab62acba0e8494ddc2f89ba22cec6871340008e11ee4a7bcc68b1d92d1fb7a7af37f3743671484c51fb5afbe8efbcd097ca76708c9d5c8705a51b4cbd8f349ece9d39188c894b1984e563e0f38407aac9745a2287011e4d130d3b19b85b987b3d987c7fb0adebd6eff9dd3d924575e977fe4a8339ccbe1a97df2b4082154081146a36bf94d4f141b1564ae64ea47962c49b0b88b01b97edb2b35517641905978d2b3e62d6619d3d42cc9c87fcecb95933397f690205ec854c034c2f1177821b89e22828f6e3277ab224c143da68487572c2722b0983516bf5d8bf29048d5942e7404ee97830f675bce0b5feade4be922fd2226e48cbfd92bd359909e8688e8d10ba0524320c3f1dd27a9280b1b74c34169b351fd619f126bba190cf79146e362969ff2b192f9b394a25e6aa9fdc17f43a4715bf354b7a64b1fd77c75a48001cd3da5530cb18a3402336f0a638fe3205cc5a0c2a8009a9d2235e3088118031dbb1f69e068243f0e9357069337c35f55323b5ab1ee2952cea3aa69741d8194cc41e8d3c485ec67293e402af481a6908e1e9eed0dafc4a022d2d29e3d4b56c67e36198b867b1684660a5a99a09d7f74e2fba1fdd8b7652f2b6149f2b5154645b5fa9640678657746887701e59d4ac8ad9e3fd83314fd87081ca3ca406fc85113bb96f5b095a18dd28e0d4179df6c7a14182483c7aab11f216fa1424eb3757e8f977b19e0e335dbcdd9b87a3e94bebfc4f45fef4063d62ed625b2a11e6158f87e9bd82699dff3bd3494997cb22d3febcce98882d37cd9b4b8a0636a0a3d773a64bfeeb89e795038dc8f96007b7918766a2f5842cc1aacb0fae7461ef2929d5e6d2f97192e6333413c7203bfea3d621f50d90e7410f08a1b2e6d1b60bf235169154797834c5c6a047489830bda0a75b4b6ae69bf075c47c194fa75c97d50c850505746208460e678e45dac4c662b319c170854b76c98f2894cc2d1a2cf53b7b72b576d51a963491dba96100055110480807aeb78c4175ed44f55f3c74135b00928f82a8aa8e905a565a0337e4172209b02ef36785998425ccd413bfbec0479b77b4ce13c0a3540c9937acf539d1f54d3a10ee49ab83442fca55c4740151b4de36b04be0de8922d46d399d79f5c5e150ef146102eb679263e758776d6e64b75130dc132f0a47c901afdb6466cbb6bc665dedb19d594f5c3e73477bd9010838efe833ee8b4b1ec5814acfa14052003eefa07427df63d2a97a64db0af4c066e789c980e41e365ddeedeb931fef5a33f9b1ab3d012868043053e7a2b0d743b253da367de280b2e70c904e42a5e2a335a2f9c3b77d14c185fd4e126708bf904bf6ccbda3d849aaa384eb2c594cc8c310de9e2330d6f89423be164fadc1383776325431c5847350a324eeccf0fc882fab1492faa655fac954f8922a252fee187ee1a0fc208582cf37e938b76afcbd16ae8df1e48161be7a4e50a13c93d59ed28f81de87c1dc12f9e36e24a68af12ad3b10af47737a7b363ac63432a093bd79dbe9ca97f739b58052311882fa686ee43a79298324a242a65362ec311d3381638e51b539464ff4e3b0dcbb41aa062ed04f556d6e210cd60569c23689b0d388bcdba898dc8ba32136ea3e2af0ec0eff8904aaef0697ff7199dfc34f1e4a9b946a92831a97226c3952dd46f696599c39320801b77757b387b74fab6b10e368a0b3b0ff6cc4a1a5f85ed6a322fb33699b3a701fc2dbeec4f538a692b56a145a085791b3f1b56a1ba70dc425552a1e67c9bc7b15089eeb7d37e960ef986461e9c064534e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcc50fa3f736390ccf392dfd5dfc7cee7ac4705a5d4242b8271ea1283bc3de251b384ec0d90d77932041dfabe2160f1467cbf93143e2e665376a3794bbc0f944272d9c13bad003f245a18eacbc1cd86cb756097c7967bdac72093128e6e82885537a7d9d388d840d10838bc49466c3717b3de155f01756d098db944ed6f2c575a12f5e6c2a63df60a694de4dfd155bcaf1e57fb7ef6950dfc6dee3aada308a3e647d0627a8ea6dbe08cc1cb003ef2f084bb5f3ed07acc49d42961c75be448e163817a158c4aeb107b179662a04c29bcf8ab5a8552ee89aba744441465c4332cb86d4d4be5a135538856438ac0d4cdeeb046b67fd3bae66ff0e0d67c12cefc4e288541782671340badf7353f0dcb1dcf7e503e1c16ec83734295893a7f2284d3a32ce1dd9931382858f5b01c6abdc9d743b2e6e8b36806c026833c116d3b05685bc42514f3e7e702ce1df742bd92b0b8323cf0c67483db62a5857f0a77ded369f15f399868a7a4ae2178c0689e1be44423e523d9937d2bb5f00e461fbe7ce6ebbddb5de3bbab44d65d0bee8162d61de9ba42bd31700625f74523b1cf1ef05a8f99f986cb9b12bf45d2b60f28d6ad16084f510924708ea86963d2a7e4139429d025386f7829c2464b71c1a0911163d2d7ee16c205596edbbf9d9d49ace9fe7cc63dd3182a3b43954f9379241638faa4fc7c6d2236242f70ddc622bc2f5fbb265707e7ba83cb49f38554ecca04f87271e40d43e27a18288550aaeff982b649d977beacbce3ec917c5f70ef884667e37e4c3b0cf052221ec51926d703bdc86ef0415c952dc9a51cbb23ced5ed2c7ad562d44e00e26cfe0a8e13eaa49f84fe7dffc306e591e1d49a345a9cee3cbcae72c613d69f6bc4e6f65e7d76fc022b3683a841eee46211726613f0b6fa6f20af1e0dfac462b004dbf35d1288a10b6dc81132ef2c171439e2ec9cbc352203c39ee9f038b6c6ffe6e3e531faba95129c3e8bf7afd7baa7d6cdce34026aa5de48cf77303adf4fbbabb0fc049ea5a45e8590a7db00f90aa27a8efc4cc53d9a04f2f3230fb2e9130e94e3064fbb5a8224a25101233baaa5be4825baae4cca120e9e44bb51a4070e1bfbc7e3d63823a27875b9c2fb8b30d55f8bad82962940eb956ece0d4bc83381082d0e43c013de4e6dbc39ee294d64d62702e2e625662de527afa3a86bdeee18077184a1eceeba51f7a1f3b47ea1086311d9b239f90ef4476a94fd2f015eaff9e0fdedbaeb998eb4c2dac13df3f5f43eac05be4bc428451c64152817780345fb8898bc3afb9cfc14e16099119b5c894a2e94bf76f6ed74f2fedf18d768607a2d564d6cb69bdaa6069cfc716bcda88cecb36bd7e04ec042b45feef1a4d02b7ea03b2a35e25d1d04a5a2f896b53b459833c956667ce03c48ed0d0d15b56a0b7c08c0e82be0b73420d22734c62c249d3be85b83aed95905f82df75db926c2d5c68218dd2ee051315f218682011c4482bda0cea1dd0c0165a4e3610fd8918193bba98fe13ec7ac2ccf19582865fd934fe002c079e5dd1f74aa9b4042d5926b58a9ca27b71f42f4163cab2a3a293230cd217d13bf8c49c27a1d32f55508f3a2b316064e3ff7800d7cdb545a38f1a1aaab863b93ab1b7940eaf079cf1f9f142054fe1b2b61ae1d395bc008345c71be7159785c8da5fb0522f11ada9444e1d657fa78087c8edf7bbda6c66f53179dc3d1fb5abd120668139346e31303ad86e09bbdf447bd47e50e9b9a41ed0524d05f2b7646705b1996a8719c161d0365fbc963b0768ddf37d7f0a803783011bc2dbec5aee5f05b1d2a5008e2a07a3bb238a1e5f7f2b27269471f91c55468d193226301940e4964cf604feb4551f38ddec90904aee43b7b9a625ba1097b101394b286e4e47605915e550853746cd30e9b3e1370f659a186379ec72184b240cd00b21d1dcc1ea548ef24b928bc60e33b465bac09869b0bcda16d1511b0b06e17484261d59740c05bd594aea0d667f6b2333e8a2b55e5bd21782b909572d91978458f55c31320b745621cfcbe18adc1bc4c7bd153697a72cd471c2c971725dda6d869a11e6e6627749276fb4cfc5510248b38a38ca74f0450f470586452356db331ba8357f95bb08c3934e2f91394fc892644c0a77c6099caeac7e3223f5425be9aa0fbe9a483548195cc51e624d01ef85c746532377fcd43ff5b703d42bbe2c1d4a9ec929f27960b2f35cc20de70940e4554706e52204307e02d60cf36a16fc1eaad2e2bcc8520ac619ff36c7c4236dac8bd8955799fc4c74dbdd2e644f14b4d45155dd754e5ab9e3d761b17a745689d634eb6d6fced7a33d5268950893eee94cd7ccb74eb176544a21a2cc2f215187b599d54175761c0636e0c295df59a6e648d944f59a3d290b9e0930f760f4efa05c106fe1a22f59d04465943b6cb8a97ec65af0ab49aab9d322e9f27eadc1f2b62fbc0b098fa735bd8afe92a06876cfbef8611a754710899a473434831e3aa6bf99d9f09f069b178f87a262124820138ec594052066f7cf548c8bddc4f46fb4a0a35065a7d96922dde378cb2de17bf7e4461eea46a36c9276e0c68cbc45858ea5927e83d28ea1543432efb29278a28688cf458ebf9c5c7df340a6240e9bec4c267925bfc3758e3095a11a40dba8061e215bb2d34a62095c2898fdbc090875046bdce58d12566a4522f634f39740162c944618cd518cebee57bbcc61decacc17a25dc57f8880b6c0a92c5e06d6207551beccf1e4c2255e6d2d3e7fd42bf4db451247ed0bb69995c256e032740476a92f9cd9b0282374f832115698e1478f46f4961c7579ba4912c7824693d6cbf8fcdd2ea6dd76d6ab21f30ebbe7e63264d334b00694a5f7ee4b0713720e8a1b5dac041621b399936bb206e4f814b56312ccca9af078fcb1c96c6d0c0d8b17d8fae71adc2dadae7bb91f1dc4ed57c6e074422d7fe76ce498183b1e31e4c2035723c5f6b3c4692b4c6e5b6b916c1c87db925ba39db5d894a11e0e8db543a35452d411332da9baf55a9c3f1aa9b3c4135767d3945961416436bdc6759afbb5b0f45989654ee6d1214d1dbcf9ceba5172e77b85de62da6e521fbe89cf4a078710ae4799abb759bd058c87b2bdbb9e0d1f8f64b13e19d5583ce015b4cbcce0d0828df0e7e2af8700451f904d5f1db0375484c7bba70ebcea92bd52e5839976a04765ffb4405fa0610980e69d0b3fc92a19f2eb6326e3ab4250e2df8684261d1ced6af64b3e4c02e76f1961bab9f6720406d43261cdbc96fbee848929ca35c38b09d72add27903a094a0a77a511aff49b22ac9023c5dfddef384b1e72522bec547547590a4ec29faa4856092ad55dbbcfe78e99e47a3abb24bc705335cc151ab1a3810d0d319a529ede122b3bee4583d09612a7c2f8040bfd1d128e58289fdda34f0902f9bd5420da5067142da85c810c8fd6978e79ded16d92014b3052803c97e166c18a3c7a39b974b4d58ae72a2cda415541736687d0a29f7e609bbce11c200495672807d47cdd0d0f2784fb7b8337a68d7684127db03982cf55f98237c6133165dc9f798c961d3dd663653effb5410ef941b972147aad21a903a2c7d88cea5f5ddb69205a5b0b53a85f22fe85baebb883228224cb89f234b0b1fd1e3dd3aec6698b09321e960bd9ae7da814e2dfa73cf311dd92a30048bd88ff3170e4542c859af74a35866f3321931904da541a7982d9fa7e90be89dced27366019aa205d56598e5031fe75fb14d90295cd52243e1a358b16cb4db0420083ac08953d9190001f7f7a1e0353064a3f2dabf4cb8ad93c053500e135488e4742c68d8b78805f971a45f5ba35821550ec7f5214572bb9fe066549bb6acc270af4f6276c4cd4a5f869f43a998dc2540ed35c95ea3a92af14df5867327546ccde7d1de9c91c40897cf4a45deff532f58e797206e19eb85576462e355974db5a221ddd4ad5d7019d89e0982dbbae20a1345f61a3eaeab2bc3dd4f2c1d31f581e222d799bcec2184bdc95b2a93f27ddcf142ac833ac51c1c84569c7e5fc9eec78e18d5adb9dda3a264bed690bc3f0fee35faf248f36168dae747723a8ea2a54aec297aa2ee117222b6008e9882322e8e409e3d2da3cdaabafba0f9bca12fd0b79f38639ce265cda990708f93265c4c70365ae92c552c2a5834ff73f7c974b5b99a5caf304b5e8a0a99f7b57c5dd4feeb42e5533f9cc4d920e64bdf68fd119257d25cb4e90dafddb755c9405ebc2fe7ded35779c5cb0a2b499d722b9f7441c445e2ebc1308386212a96fcc5c824e931b266ee5779ce24a5ab3a892983d22bf1ddb504b1f7415a9c474d90c03bade13dc2ed6d609fdc42205012c48a227816443102b8e46f3b5fe92655831b5e206737087254e5454a792abc119c567cfdf81ecc4415e436f380732987d685040d4d9eacfbc0df86179e18d47556a414a94e966b98aad249ceacd48a6496c2e54749bbb700f6c8c10b8f4c362f69063a4a3e81fb8e86cdb18783493656d5e8c6af913d769f8ecbce6fdb6c478c14d7b5c6ef5a8b7c5fb72a71ffc1e29a9854bf1b03dec2bad3971c19719eff6fbe90c9159db0cd8a77aa643eaea3c93ecd30bd37f8b3747ce3cb37bd0e3e8a65f62b9e0c5860f5a46cf329a5a2e228fc861c32ef1d8365e0f1c011f0913fefa6d7e800f0f628f9f30263608d313860b4894b76cfca91cf486bf681135f11e1b2c227e6940c0281bdf3695979c3b81faa1d84a7b01f4c633fd16d5a2d6274433887f1b7b0088a168be70642023588d355b483b893721ccd8c44ef1d8a8f5987dabbd8c50528481b5ba9de337e04083c721f02115157f7eccca3056685218a14b57f677946cc807c859c8836b0d976eb9191f6aaac63c800887ffce0d5d92ca19f5ca19c68436e928d0bdc5e789200984703b9246839f9c13c2fa38188827d5a65f50ea610ed41c8b58a72625a0119026c1a772077575a540e6706913efded3caf88b6febf4dda2b5029473e5c5a07a0041c5e3173dec23bc984663548b3414ef24f7de84ba771c59b1420fd3cd16fc596af17d7c06a0f5a14d07a5a2df9de0e44f1eadda703781062449b78127b3c55d75e3767ac8724959458aff1762e450993884a0fb0ee0b29bc54eab9bafc66d00abee746e4b9337a5cad00d2bc2f909a277108e4addba92e521ceb62cc3bbc713e460f2a2eceaa098166e4d6abe2ed00d198e900262b20febbba150618f6f551e6bf8b384aaac5cb92f3e0a9ea13bf99329d73cfe196bb28aa28a91a08cc452d90b7a5e09133d0be0a00ed2b41f8f232c9fca13451431e04da5993595326caebdeba1040560e3d6669eaa80005f8af22dd547bab34d202638c9a46b515bb8a0c7d919087078af0a9fbb12f36a131c916417d033007ba847a0db4d3b61a3e94de85c2f63a1153e101532ee464009f549ae7ecfc83631c58e452494c9a0be80d6f583c8b75d28a9f7a50456e7b716f39a6254b2727c0859a6c4a55042e73c811bf5f8f12f55380e175caf789cc685926068bd599255e6bcfb204548684968a5460f629ac47d5dad2129e05e9d2f2112fba9fb46ff7412ce1b2b96592f042ac16ab8783660723f6d867a57c067cff0f911be60ddd2129fd7f570f95d24a50170d5537b5e4831fe8531e996cc3c98e22c94f7035be415c7e152d6f33060334d64518ce2d0eb2b4cf105ce098a1dae36569adf4768901d4e4cc1ab8210b762fe490fdc6df51b1a17c6bc6f1783e12e5f37afd2653a2976d461992f2bd114dfb302b0d946246d4d0dd822fb1c7e1b9c9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4b21754a06214d87ad73bdf6a015f45f6498b90bb173adc5eaedcfd1f68dc8c483da68829367660534c264f846f1a6fa450a8ad0f24634e4ca5b7cc28b8041e7092ca2d44cfd5af1f86ece55eab9d2b34ead99308939ae4e20d92a71c9006a9eeaa348ad42adb4c2eebf25bb308142c50c55d97014ecdf50ac3a3c1dca829b49de70f3e5bfa972ea07a1c34a1adaca40d90890386c1d18e09b195bfcb2b94fd4540c533593ec6c4c2d00c438695a6a107982a830dff5d4196a070c293aa8dbb7daf15754d02b1ed3b36e560c0e132a9844b0c338d4f7ab6edb2a7b9e74aa42bed307e018ea58ed4dcc91c290ad48a1d67468827726d52e9d96b5e7295372b24bba88806ae1490a372951e1c519d85f19428d43eb895bf5644db76aed805b9bc47cde3d592f3a71f83ad0da07fb8c7bf63737eead7aaaddc8e09a3049ae84d592c5a4c30509ba2c7438d7e7613f031e351c91980ea9b971bbf85a2fc8d7ace83324c69ead7785e796fa73ce48e56a60955fbf3708f240ddc6c73df2bc8d22ae95a4ca11eda637a7e650cf5dfc17b15dfa8dc705d1f640b471ff7e47db05dc9287421365b87ce3efacb64ae567af953ed7c38bb171315c8610d978ade0eac8123e51826d59c19983bb38d6cae5c4cfc653dffc21f346e0acd79b659f6e3cebce3ba6b2820dc90907b32f9fd5e2f010429d8e49665850b0189d8a972cb15a36abf9ec7b2eb7be508124ae990b7d90085d7bff743c5d1aa8e341c0c74c8f2984c38911b477b2fc0d48a45f4a91458fa934aaeba7220f9c1f17a628e659d97921196253e37af25af1418ca32a9e41782f1c06bc0142b4023c7f6b2e96e06dce3e0264e3d6e0c539d2a214933d35f217a5128c98961bd48369653d5037077ccfa05c13d3499045a570d8f41c9f1047b2590271f831280eeb7154d1848141737dad41ab7b0c20a8f782c50b267c4d126c48bec02da1a0238ae455709655b98ff7f6d549438710edcfdea00ffa92526e8ed5d977ff1882c67c15fca97b9d4472777247bfc97d5490c7b300938119ce1deff53373b0362e08700d7d807ade7a6eb747d205a5166cad6171027cbc6c9e261dc4255c83939a8f2831ea2568ee956144beb21e002ae73f47d0a8dc6fe2e7f4161eda9f1be3224212212cfe7caa7df339c2f8d87bd666f50c5d13f54a4186fb780502444c968f283c967d8790ac93f7ebd63a73a4616b73a87ed9a9d1c6288b16ccc40ed75de39d22d087d38482cf7435584fce9967abc5448c698408e55c4ec59326fbb5a4e52ff164430ab9bee5209dbb98cf4f9cf7b22c70bbe79160c63417be95b1c03aba10839e9e1553319b9ff130b014a74e8aa7cc2b74a1bd805f1657977c595102bb5859df9eb157bc10bbe3c7641f7c5a9a2a17e316c42ec80758b862c3c6943387f0593f0f0683bb621c04b22219292620aed99d6dca872c7d515c320794aafc5fc2be99eb06c2490c9673c4e8e2763671b156b4284d356dcff9ec4df5ec3392c4dde426f2af3b4631abb4536a202007bd07d1fa62f0161d775d73ec698a0927da8bca4b30d32d52d10f1c081d7d7d0dfa135c5b27ffb89abceaafe193e0bfe290cccf03a800011957b8079aa869da2e3d95dbd5a06eb38915d3fc7ae2860e9d54fa68621dbb48f1c699cd47740f2201c2b65f2fa7c07a98a1a0f0772b148172e3f9cbc586eff1f9e70a3311adb25c22470f9c01e6e668f0029beaa20ab94a4a056e2e511f19ee3811e2629fa0b5a113152cb769dcf06e2de72575bacb901d812e418c068dceda875e385d6ce8ccd2fe4d4bfad1efa61ee34ed8e225b12e5d69baebc62d6b2ff6030b30b60f71ec89985cee0f3e1ff33c08bdf84159c8be8e7c8dd11c86f10571344d44976a6d3c0da61dc64d656913557b9e390649c1742b87691919229343e062e5cbeddd5d0edccbcb56e5cc9c91e157c8f39c04f0c7e2913ddd37ae920b398973ab7bc82678da2ebe674f8579f76fe1a835ebc21e04190acba290056a4abecefe63cd4370849d2dced4c62c90268e1ff23176e17f628b159cf809fdc173bb3a712397d66901bffd7c2c3b5fe91988f6c2055bac98e34b4c675aa5547ae47c45d05f3dfa030ccc4a5fd9b5352d5abad7c5ee00b50773e8108052c54580232cfdb9f396c4c0608794eceb8efe5d1488df64c72e3d17be7226f3f931f6862131ff5be181913a2528270d99e713079e5d706c3fae9e91a88dfeeb7482906cbcc5338447bd92205af47f7aaccf103be15a2b55b47ba11be70c8a3275c9f5d8f2f117a4b07ecf24d4678a8459b74f9c36e4d5bee72a48a4e84a22479a6df15ecca958da8883f51090750f890b33d0e87fb0fd1ace2df2e335a86601c9011aebb1112793fd78fecb35065406e0c89a2c168e33e6ec0621e5949b7680fcaeb6d3025103d8ca875fb28a09b8bc3cb97c3ebb1cacf3736e1ffbfc823d73931027c13325b73c644fe9cc2633d1ebd62a8a9cbd6531e34769d3398d065baaafb09f031f62e9b1c706567668b3f204228593d1d2d34b98c12b94ef2fbd5a43ed317f7e6aa3e56f1b851bdd385b8d7046e466b0af42d9a6d2db60f1ed8d430e58c9a46d9962ed6ebb37a28c9835603c265fe1567a6518706b47bf6efe11268a3c158361800c5fcb01322bb8312f7a142fce6e0c986a1cb6cc1ca32e986810367c79978ab8be5e597b93956d17565dc6ff167ad073dfae3db60ec3164e761e4cb05a4489736e62088b4a66d44ea73159ab86fd9ac3998f4df2d55663031baa0ecd061489dcade06191e4bedcad2eee24a80aa35e38931fd1da645fb89e73f22482e5459dbb5007fd0da2040459e940130b22216705c964b196da6b71e8b73c2753b4491e4e90492baff651bb1ecee23347978509fa65ea9281c93b812bb3e9ce81dee49eb76dac34dcd8f79a48786b4e9428a9791a48c97c520d240049aebdcbff9293c6af756ea9165185b56597342cc75e6e3295433f4dbb1a49596193955e5181feb2d1e77071d323f2ab79218d5d71dd9d2274512d946df20402a8facd56fdce7f2f8cb89a05078ea993b4b0cf5f6091b7698b74745ed57cf965e6d2b6d9f8c6beac13c6bd0b0947eebd177d44bb66cf5e2f23c436f0e1f7fb9d32239d462181cb6e7971b31451e307bd59ece584b63185b7d93ff05548938342646689f3f193ad2a48950716115b4419c52879a47922a4ea254977d56204efdb26ec04a4d3dcdf680df6f1f843767c23c391c11eca3f768d740a1df78ee2a0f378ede0c7ce37898e38e78a19d2a558067e2c4e50c122468888175ab7a8985f02588db44c85cdb4a0d0eb8d0567cc8a8cb572bf8348e8372ad7bf1764276441bb19863664263fdd0a5fd1d9d2d14281f3fd88c8dff5d34651162c110358271417cde418a56c84a1777efcebade5f981dab59495999fe596a6c86aa22c933ded5621ce6d27918ccb3dc493d5186172a4c8d28e288bb014f2c54d1d7606b1d1094210be80865ff7fa0bf84878f9d8c77f2bf6a0648a199b838c12e075e4a5af0e9cdb98f62524a0feb21d11b7c268b370d51a4ee9403ed114c3a37d20fee311d982f16eb1cc2f0989098f3e77bbeddba5072ed53e49f094f93f3db9445ed088a61cd0cd6d7a303d8a96157773e6a7114960e4a9e836d1add8fc4d2bf2815382ef821b015e0add031423386cab02cc9e11ef4643b1da05d9c15b67e1f2488ba1146516304bebb755b32dcb63858351550f4d508f44cb5fff46ec6d0e20a57120d38a7da4b266e879b8bc227d2a70d74d05406045500df0aa9f2a1994710092fcbf44f904067486b10aee38bede8e14798fe573a43df0432344acb84cf9d34bbe35c3db75c0771ce11a0bf99756db0b1fc4b151d390c615aef6a24b4659c00286c21b1dc2e00a3188efba2d3c82d6884913f818e3843bd4e5d6d12f652fc40807a9f4d597c1e2bb56eb8fa8487a2c25ba8153dbd0c2a5fc9d42e670b77d20fe522462f9bb0bb9abf7570cbc79702eb0054d8284c34bc4ff1c2020bf434f43ed1804abf21888f6750748c410040bb1f93aa314589182b9d45cadb96f04f51d62c289ed2faf592c04ea1fa96554613e9ee816d2be1f64606d453c3d6cdd8804956e4378fb895a80956dfc4b84d72e7a0e3b3926f10a0a60dbf481a604c1a8568d1fe216935c6f7d1e8a96cb8e262d2a570c9a18e80dfb897d93f2c63632625a385481ccb35342a6f803f5a9ea68263e7bde39efa6e4d4af141feb2948fdd624b54bc9a149a41e416efb5117f2f18f354d3b9dce7f21d862d02bb49adbce5de8dee253e1224e51c463b7be0c21ef6e84ec9eade52eac613479a120bb2f45a42bfc61737a42c172bd833ba982d59c8322c172cdc86f386573e7edb8d362d4ae346aa012dbd602901b65f1f83dcae6e7833d8b2c92947ce4fa086f2c7a217f0777201421bd1c0e40c9aa9b0b70c367eb122e0b316a8528c88bf26b081a69492a6af8e183810b671803b3cea6c34593c5f9e5b56dc7cfa157468a01acae73163672e3c739de00cd6f3fe73d62ca2ab4dba7d545abb100d8da17ecfc2f03dd9edce404f4aa317b31efac6c354f5ff769024a989bca3fa36d4e8832a1a257fc8a2f5038172e3a095954e3fe5f103c03d2094ab2ed6df71ae933ee4d877e0b18f89fe89184284ed7a47725d4fdf70195266b9f697f0dd435d5392ba168fb0a0e15bf7ce4216edef9eb7cf2cc5bfe16f8aed4b43d5ab1241a4c73ca903067ca0f03dd72e50802117d20ad7ed85483a9f7ca8de434e9c4b8dde7a409d17c02050518305ff676064d70a1678aa6bb3cd23d3a445c9a85d8073754b15dcae916baef487ae730403e6c522db59c751f92a855c2a50b4314803ff950155d382850b1387c58955170376bd9b16ad2a644e1d50480b083f4ae8bfabac8356f965e2d9464b79c4a112e63d705f2a26a78dbaee047360437d0349589043bffe2d8983abb6c6fd9747218eca87c08b728a387d6349722c1b5b4f91943810d2d4857488b9f46a7ea50c5afb24b1b9775ddb78d036d879265e9cb119d456a80340d6c5442ea63324fcd696c3de93b606854af4e81aa8dfa89bdc2c1af56ae8f6ea6315287c700e7421489ef48f22f5d4d9aac1d7ff20766c02dd95e859c57a41c20c786f2d950d4e419f5185ebbd5792d7a026a55443e22626065d6bef6d0920d3ca7058e327903e46562061ee5c52ec76199e7e2dc9ed1ccade5e992d50d065b253238c193220c6d8a34816ed2ba307694233de08a8671b33f96e9fefd7c0159521f4afe89d6075cc27afb78d432268b2a9a5ddaa6882dcba84ddbf57b378a8ffabf455403fe1b2682597a25a620c275de3af9ca2afada526d81c993ce6d09bf3e884c339beed945c6fb9c63c1a7ecefe0ffa483cd4260d10d836ce4406f89e2f8d8cb0e9a58d9180039ae497959f53d40057466b826e2c05baefcf08ace27a04d88379ea94d08669fead22ae3c0e0524b32942cd8594b7d8ad9d7f7e8961368ea08419580585833bc97382e6009e1a9694ba33ba14f445d58c24cb1588c731222dcedc834648365a376ebc7f0b6e14eea046ccc36dc596369e6ca070b353bc4c828a573727c34f394f0449fec8f5ab85bd0f35c03570b9c203a695ebc50db7494340405f21be679131d1d43da45e54f89515522ae0b2d24258e6d0000fb8c21b4d8399ddff973971f3d56fae8a8707959c174c159ee0ae57ff007c943e4a04445c9bb3736957300f6d3ad11ad81ef269cea2b5f2fb7cd3a75d0864deb44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc6d7a5209c6fb40fba412c9178aaeeb2bcf016b075407672dfd44edbdc58da7e4f0b67c2f3a28e54e33d444dea72a7587a0819bfc34ccdad27683be5cf4ecde0f00f439dd84835b9f0b8dc5ba0f45ac1b00413d0f347ebf1f5e44b5781ae403c7b79efd9500319cc6a9abcbfcf89b52d56f226f1178dd1a9e17dbed1bbefbce2e94b4f817e72c57eaa9eada55baa61d24410425c9d862293847506cec52ca30455ed677554e59ee17b16a19ac6bf4316b1379620de76d58c8fad131341e08d11cf66e8f67cf0202e2bd23b8c31eae844afe6e78f70c14efacc177d9ad769df2034d0ddc7d93732d9890a441834951e7512242c1e47d3be1ad71ddc82fdb2db306b875a19437b0c48eab64b5cd7237061159f25db17ac91f7d2965b1f4b7fa99221b8b76f231ebf7e4797a37caee7a54c2fcffb12f06d5b83c41e2079345013993f16cdea9150360051ac51499b7075c0d319791a19c20cf0955c3766426b6b5d4e7e204c03d46ae14d3d6496f0d72a09dcf2c17fb7800aa49133784eb74b5d34e143a1e07b5b19d2547ad307d1e381a9d6509d63564a6e3eebc64e6586314e70f5fb9b9bb3371f8c533807194fedf41367b0313b8228313f13840ed5fc96e2b093743a74201e2cc225db8bf3609ce53e8b36b972496538ecc25da28248fdaea61313fe87b7b47e321fef28d423eed00a4d00f2d646935b0875117fdaf7156626bd36a1d0be25290eae5b19d042465efeff0cb6906f531754d5d738facb45573589f54d6ce0f384e172174b83ec1b3f13f85cb4ce08b60d685e9480fa8db25a9f8d367b0f9fe2cb4783ec6e11f2a4ffe3a3175950c04931f1925804257efa328263f8ab8de1358c60afd258525752c66eb097c61d99d7ff72c2fa11b09e587b0aaf37792820574bc229e8c43e3493581a6b7c64275f694160d8d0f76c6f360b78585267b90aced33c7e43df86feeda36e4429c794e9880a2cc32e774a09c81597fcfc295ad5d8fd83783323400052ab9ac91d9fcb49cc5e30fe028e8607b7b7fceae1dbe48e117051bc234e7c91ef07346634c5361c18e673cb6135f3d8789dc9d5d6f1d64c1f84aee1b0286f4cfb507328ffc68c78255e9226c91fb5c34a7dcb4281b76090032b77104f5e5f82cadfc74f81cf309b8ee34d51bc603acb10a8be837ec3a2dd5cd72997df5e2e5f4a60773415b9dce10acabb0d5b84620af0ebc791de91774df6dd97f2ecd12356dbfde8c3d77f22dbdda40ffaee18903378e8cf79139796d6eae881e9dab095aca5d78831420f6cac71daf88b140939dfaa1382af0d220c86f2f0f19a1e208e2d1ac6300241f2d58d8ebda9c33bc97cad2eb02b58d446ac4bce73385eb4910cb94da6621f7660db857c250a2283f0d307a7b3bb092d754cb36d875e59c84c054e157459ce19bbef061cb4920c91dd61295e36aa173218b0d4de5d9d6e93d433c37fd552a31605291e4d4dcc10cbdbc8d001df17c6e57407bca9430361961eb5477baf4c2a75d3be081568b6e92af83fd1a06f88ba22bd6dc914c3a499c59177b849ec229111dbf3322b3165dca4de715f6b1136ebe832caa0d4334f4994cf4bbbb6d08c551128985baa6bbb41452348e63e55575e78e0aa3fa8f6abdb016d72acf08e44bbaf96c3922f04d3cb43d682d391512f504c8e608ad9d639541d71d705bf68d0cab772cb3c1f67496c0d70f393ed28901c6baee9b86bfbdddb1a9bd38e00ddce769787c09b076ee95ca0013ccb8b5e2f7815966fe0baeabeaf511c7315fe264ca2b201c895c058cb2f4f6593afabc7d87abfc7ebf0d794144475e0ec46044fc17e59ca36dd5f67197586e040c745c550bbd65e99fa95d8682cf21ce3ee5ef0c27b67007e83422a71c66012b4b4bb0114169b90a0af99d4d61249b0795c87811718dc0858b6abaa50e2edb55e372555dde9a814a9a787e4e428f03271a69f1abc489113138dad2f350e592e21676cbd5bb889105f5aa4943992758d777db19c9c3bfd8625aec1162ee9e795db8fc8b2442ce8423132472ee61e6328c1d52b4f1bc700207ddeb1392dcb38c1c30944ab640b4b45e438293e23d9cd36fade05a3e0788bfd1998687b38e9fb80296c77a539d022cb1d4f2b14d5fd7a0cc1edfb3f947ca78fe5666bc47e6bc9ae3061bb0f96ff0522725292cd07fa46364bc73c134309cf3e1d85c4f345b50eb67a3a36efbf877bd0516e4c57764e222cd1927094821270dcc82aa6d916ea58a4f1a646c3676499d656469d25173687751f4d3b710e15835da2dde0e1a5497bd13928dc0d647778ca0a81cf53fe3fdf217813bdf11da2b0d5089ab072a85281f59c315b155b57fd65f8cec1603a70aa650a2177d64eac90e2613b8227e2dfc5e77933c56c9a297aab41b2ffced64252d263f414cc54a95123945c71a425ab0a53deecde6c44d85645f0929fba6104a38b400b5c5c67710779724940f22a16445d622a76fa112a1ac3cb65b97a50680648a1317c3a22e17c80431094df6e915c9d52e97f3b9de96a1255d0e780d00385b31cb47e7f2d00c4883d0eb4ce0dd230b0609fa876686dbfc18a1e3dde1b2633533e45e90574b06d1871355ad8e6be2e5f9d2728c8d2cf5b0723649c458ee85e3b76c220264d61200aa9f4a3384bb74a1f389c51b3c2c778a3b45de7b550815849d0efb097bc742fe989956acfca74cbb708aaf23b6ff425c0be1f7fa3dd8f4280617664258c63032f96f850cc57c816c903aa5169639918bf75fba0a94802b8a7345e89f2f8a5524184c8b8102e0eeb61ba768550e0ff49da4be6d2c9ec4079aef9f7df0b43d584a88a8cabfb6b096f1cccb0239bd73ffe737bb47c5bd53c16fcef98100c7e0f9b073aa79b9eaed5b01b21e0bd66b6636441043acb4d906df867056bbebc7f83df075a22640c49e7920063cc11c8771a1f1beedb8b2123629ec49e00bc1b72074225be4e87a48173698ba0207c71a8774da91f25022988717be9132dbe7fb03c7fa98141fb06df8cb6890eb12c0e39e16a61e11eeb6e36c1fe968d3908a7360c9691ba0dae3bc72d3fd21de5b652ec341a878f02390e5d6bda8437aeffdcbc3910b975a74e892f36a1242f64a5f30d6c61e50e543fdc49d4f1a0985cfaba2f6870cbb9fe2ccffd3cc7ff4cc1f571c55addd111976a8d27b70f37dbc0ab7431ff43fc613bae1143ada9e5b3b5412eb023e99df24c2f744f980aa6deb8374a85ddbc4ebef2feb01cf901c47277b77a9b512d124b19d9caf26b2475386fa934a17b7646853546bbfcc68f298c4f7e1ea74952f14af56c4829b0b2e3fc48f50960a2ced7034b1a2e81e753cd35d3b72b6255a6284c855978a2f1dbec0de4688aa5c96827fba599b5b78433936e2c88d72a84d7eb06b003acd497735c619c953154379966945e5ea4e344af2b7e7f024560b7d8c24d5342c345ce232975a4dc8a5622150b7906134c6597645c5e87f706bfb1029188e9a5854eafb3d0c2b3df8d8e802c3480fdd4c29bf6d075ccf894de4de5e0523bbec1a97ad5da80ad1017bcde9326881379efadbd4e7d245d5a41167cc00ac8715cacf829f213e57bd6d5d40f322057d40ffb3784fe213f3e032fc4142294e8ff6d5a900526c674bc49c10a769780a5bd332eff0fa00b1fd077436be73656444d47e75c73d36e0f4eb74c8232839ae39944c48eebd315664bc18029cf85a3c5748c7f60a55af185385c3acf83978aedfb1a0108e6f2086d2eed253a71ee1986639f5f640faab0e027c6649890146f75e0e65841b77aa4a1f636c0a40fd003944a17c36ccdf39a44ab2bf2665a6a1c5573caa59b70ea9e858e75ead2dfaa30101c78cea3a481bbcaef0349205fefaf334c649d5abd194d938fc1db7b763e93fc59c259d9d7913f1cb9eb3d20b3e2edac76c10fb7a82a0dacb91405127dcb4ee57ee274bda14fc63be8a72f5a5eb9703a997f84cc8004e9fe0a9a3fdc5e241fa8e4b1bb5fe8afa8a97b7923aef805b1eeb86d1dbb05fe87a4f3edf7992f64ccefd3334f19858babc90131c5aa01abecb5699cd80f632bbf9bc1a33c34bd5a0513c9e62aa5b689ca4313b29b855999df9265793be3fca18318357e7e74ffff86862db7410eaef41f740e0d79009709465b2465f89065f580959c31ce655eb6fad2ea47cd831ef53947a552e9b8eced2b2234f747f0e2070fd86beb05f071ab066711ccd3e744c70999cfd979cde04e90ab0673f2b572126d698948c6e16ac579f465c76cf6eadcbfbd34d9ff05a60f0be0c729efce192867c5f1051f0855e224615a4a39c1937d2fe97b000cafdb477872b969ba4591ba80a6d5c25668c00b71fe46eb04d551cf42586b98e2ebc8d4a13ac45b9ef1bf906159cc2faf7dd9bb37659d37151341d8f9e35c522d2f0b05f138959e6dff40dd2addc683ba29bdc788f711caab1959c35a4c4a77688bdc78d1e15eefb11996a2f7fcf71f97b783b00507a414560b476d28ac2ef5514e160ebea44152212078b47428ab1cdd2deff835ade246a0b41897ae9db84f8a7ececeab170559f2fb792d68c3f40f05e30f94b7884ede122de5c94f453442c929de8bc972971173ef8c4077c672beb5c9debae118734294e3a7385a0b0e785d9fa7cf8f70eb3fe0ee37c56bc407d259eba77b72203370cd3f581b49e3814e9a44f3fe5b98812212adb1ad2419ec2e4a5a9a997fe54427ad1dad932a28e777a52750c010f7ed7008bd05fe131332a189d71908221d65751623e3f190455333c401db55dd13180441e6153455295f4bdb45b7537d6ea2091a4fc02e9632be2cca144e492cc5c83b3f829e2f482c664fab0a7b837e2a0368f2e75d960d3f43193eb974c5e2bd15a9b5fb5b5621a08a1157b3fe62f2d4691a7dc39a8c066e2573c848c073938b1b4f86fdd4de5833ac3ff96a5059f548e12a406bcc9cbb5e631fc98e07083031c95e7e2090fcc62aba2454aa461655217e50b2bf84a8bf7fab7824593f9b008b0bf898f413a80dd90a76e9bc72bac93dd2968fdf91c4c0798628a740ede5146e0267ebb732c9457bde5e0f8ca0bc0afd97cb3a2f40fbdba439ec28c35b7f34769a2650c7a3fa7ab500ce8e3d3726c894fefecbeaec6051904c0df80475b5b4ecf480e27bcf82a941ffb53b4d152b403c9a428ccce689e80316a2151620ee6393683a849915987da77a80586b5900e7c07a4f75443d5fbec876c8c1738149e329fdb1528224d6a886745204e54b5c842812c2b3f7c459f45726f932be714aaf411ff1193865f4c2715da6e31216bfd624eb8f24b6df2c731ede026f87c358d3ca50fd1eed6192e7d14c4591edf9026d4d29bd5d675e7d0bd05ecfdccc7ec04534209333cc9061987bad9e6607f19a5543d729b28fac92f9197ca0ae0d15794e64cf86620429924e6ad756fd2e8515e71ee9116d91ddd392eebbd1a0247671c6cb14d992a1b40d037ad041b04f7bafa4f1d34bc0f2befde104ab921f4a1614a92804cc0421747ef61b4c9fb554133f0e11c132a0f1a7ed0434ec0341a99492c47a23c4e0378bc3a2eea5d4cfa00dbd32b4d110ec3807a252e66681df6d00c30ef70ab13f00bd4910aad865aff979210da8c148e172885bdad971fc579160ec5ce7a726027f075826e3a912e8d5619dcc162843977a33e1127e3a2c07f7587b98a1d9b1e439d7b343d4c9c132fcfb1991695bbc201e7effd96172a8db577dab436e3b339b3d48b2f163163cfd3f41639ec2ba6088cd5f5cc4e6eec7f479856eb19254b6ee35603f077b88feb6fb7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb60f4da269c053ea586e866f77a6922fb2acd3a107b533079f185851656a05344941eeb81baa76f42c54788b919a6f80c7ca410cb3e5090e1ffcdcea56986a9896ed3cd247702365ddf7665ed2faaf39fe42f6fc75af8371f3abba628e7f605482e9a259cf3bdaf33f14fd754770a64533730e5d210d360ca932844d9327bed3e121056aaac58a976e71e586b49ed753daf7de73f6d24b449d5e498f267915edb4c153b9301358c75e8ba70eadda7c87d5fc4d772e03405afd9ffa6d55213dcee0c05333ab856004f46a0d734e3bacee02c9e7583d2b60c0742567ce2fc8dba7fc125975f47b055731c0034c71159a1308291465fa35d1063ecc1ecfa34b0732e9268490b5c15005f12848d6755594fd82509c94414d1ce3c1c64e204be3e8ad6bbe1fe2cc2d5e12424dc0d7ffa35644f78323aaae4146226bea0269f664e97e90c9ac4e71ce4ae85970f6af4034d374c68be11df1726d51d527449628f3e91e32c89f3388f55853e67bf4da5a43b6844ace093a3d4c0b4c82e386676d49db38d06680b324627747470c4ce82a780d848b293eba364516b268709240808ba37945f0f33b3ece1ad188c0f64c66d4d906e9d9100bdaf9174fd8001f245a1870deae0d90a59c2db3b181cc7728820a142acba4190d309ca207eb9545f5c8d82d1e81daaea2dcbb6f941bff4abcc434484d596af40c4259bb5e0729ef61c12169b02098e5eee417bf4c3efa9a07417589fac46465ea299fb7cf46fd4e6c36a4244f07d2988010e1c98f3e7608bc6e8af8b00a1317ce36e33508ee4ed1d773046d63c59cc0b0d8946c6da09f3dc3a065a25b218d330bd0512c360e9e0de53b05497693f90ba87581e50c5702f19778c74dcb2ae9afec532685c5571b4ef9a5f39a96da8bf9e1aa0440600a97ba6d0a4e3bbec8c420f2c90205520c22140dc9bd464d0539e9449c0fdadb2ba177a96424ae87c8746e7c91f88bdff706936667020ae48282696635c5da93e4296d33d40c62ad4e9ac387f29d10af35eccdfdc1e23060d995797dbdf818971d1202bda9589bf0bd1c6c5d8a43319f53bba03f46b682ed957d6b88a743d74a7a9727fb2324e7636e7da07166e1171165c9f30b924fa00730e5d2f5ab849113a2760638a493af6b2e73830083c9f4411c47946e34146acabb7161b26d40a731e7e7cacff9b54ef39751b7c9e1bf925e522daca21aac3e90a0aeacc58fef1f704319b3d4076951e154d5079b0d10520fc8a8eae7d361b5f52ae60e76737df88fa358995cbca059e8405fc984f8b7a990e117bfe5c65c88f8ba3d722b07915231e6aad2e974a267755d7f3e131f0c7c1edc6aebf671a65d6fd5655d3f7da1b6634731d4d98a010ed91398eb123b2b9a7162968f5711e33f1a0681f26ed8c165e43d77afe685448d0ae0321d8f8543fef8724b1d5d568b116f0acacd2877f4b83bd9059b23188c9c493faf6001c5d465b469ac07e9d8c15c11d196f86a2e5eab2341528c0084d2916a0d71bf1e38387420251586f7e9f09369779d9078ae793d7dbc633cc158bf6f74744b2e88f892e2990197f15ab5fe4778c19ac5b4add3fec1a33a7f3e7652ac8862dcb7d34beb9ae0eb37faf7ba0cdc7d1b69fc8069d7aaa4b0bbc565f4a5f10cead26ab02d2f6db6580bc612c2bed38059f274b19fe4bf3986dfed104f99279a2ccf3104608dae36c70ecb38ad491e66f4a8ec28a36c48fded9c3e4f5984bcc4ce750cb883c229ecd7f6a3df5b1dc673da254f1b1ca84d42203bca541a3b3c83cae32527397bf8c62b919356f61cf0ba643c9228af78d3c7bc6ccf2255cd6a7c91a10896c1f3d0230edcd96f829471e7ae9c452d98ed079bd5bf5af92349f45bfdea2076547fe4a7b41638d37c1ca31923189f9cc4caf13a6f6b5369a8b2d2a57a63557f83412726cbf6a0f1411248b5b19e7c429f3c10130f63484fb739649b32395a1b3e45f1f2f2077955c4d95232f1d4fcf9578932fa95074e45d780600c55dbce820576e94b41c3b9fe06f67a953fb43159eca16737446b5e0e7e7e9c1a43b0342d3090ec63995e97ac05b293028c997f3a10cd613f6094d0f94815d0bde75bfaba466724acf3a24d82c6fc5e01477655dc7ffe67d0af7bc72012403c70532372d64f4efde7cedd52a73d422fe651c1a4a245e07f2d8c1fbd30691214a92b36eea98aab77e48f651e7bfdcfed60bb54e334b80bfad1bc2a0bffa1d514eec8bfaf652ca250ede3e819fedcc56ee87816fae2a6c4f386a6ac0b4645f927def5c652529c7f5ccff85a03002d7370d95d3a0b8c1fa2045dcc4b6d7015a3fa1ed6507a5685724d5eedea0385b606b26ce8a17ff35255398ce0c5fb21c235302ab7015d645777931ad97f5821a23008bf8d10cc488052adbbbf537373613bbe77fc7fce4f3d7988f24b281e1fb72745f496ecaa2c1af8f6f1a8d7d8a94b8ba33210dc5251f633c5b62a3af59b1b55d0aadb091d87866371ff2be71381b54c340db8ffdc4c6f643fa944cad03d854d4f609ed77dccee9a67a93eeb22ba39be5a166ce8f28e2a950c7199a2f54a267b932f72717be1bacb68f0e78371842c352f87cb263aaa9e5715523b0f2b5e38aec2fc6cb079c758cfd2ad74609ce9cb9f3d2bb618670a7fc349b5907307f96335c84075ed382f00f260bbf576394d60c995d950c60c9f61800a5fede75d36a4cc8455a0ce84ea5c231f1c289f074195d99a4e7b2cb7ef6ae71f51fe8ec9d1b8f2fdbf5e5c67a4ba5b49acb681e8a2ec172977918903c96ddf0eb716e21e5825d7990fa77867edae217c9bc8048b450e8570015ceb579ed1217a43f29c534774677e8b6fb71a4d5d2113734b229b87c3c0151295419603b0e10015af534f56105a851305cf0c269c656eab0f9da1320ae2f67afe34e0acb3a2acd980ff78031404cd36812a4fab68725789f73e88d7ee45a6f86cfe4bfe8edf9401ff8f801809ab668e3f995892e2c2abf427fe7927c762f54936340a4b9ec8b65e53fb9bad2aa32ce30924943362aa16ee9e76f4b86264c027172cad6222b56cc736b48cdbbe2183b21188544be21834e5a11c0ff3d9f6333c411d24e1645d1f334b20bed20d8e1ec5c06447825b2c85c7175f2f14beebc4de54aba6e22c28ae8873b5b968cba762dc38c0b92fa3b0d268476078e31ead6b1d7c6efa5fa7bed9187dd42e56e0a9824ce15d5fa98fc5100d23553749d1cd147be6107ca23537f2d52c1e69a852ff3cfd55a8dbbea7f025df5ffe1f4e8e0d8a879f5abb92ec7c80c594f9526fba185dd4868e284f7dd7369a58bc32b066bc3f1fc65d9297e3e80698cd763434d65c753794c75d19c772353ff54e4b19f97f9c815c3c5e654983b4011e7b4fcc61d03cc188db9fa1c76233d8b23a26e6fb70aaf73d64e3016669844b212b2cac5f57fa2b01acb59785dcb6f26ffd7e125a85140a6b75ae425a9c8d1ec0768b8a2e8b914d45c68c4d4a159c39d00ea734cc417cd7eb498e6f7ac6f05febe16a17803d0fdea644e39062dd3d3621c7192fa3244503546a8307b5343748fd39781458e449401f4f84e521d5b861aabb0e3b3a03f6e269d49057507389335d4aab96adec711b75fe0d770b0672e20a0cebe8e7cab47c0c9f6b9c647a88b544d6c447e485bf4212ae44c4dd21166b50a64996c34f17d96a7fa8b49c4e739d2e6c1dea5e631189ec7a0f14ffa5315f51b44a9203140d08df905a886059ec4f0695a2ebe4b1f7825c25c70b29827ef6e1ea28ef2c7253b4dfa97ae11bb6abad2d9dc5cae7b2455c6e2212f77d2275f3de6513b56540081866981605989b0ac2b16102126cfe3ff6f230d8c5dc511b58145ce1cfc1ffe8dc7e2c65a887db4b2d2e2baddce08d46495335dc3cefcefeb008e009c9f2b14a6050d6314e96e1f91bc5b9cd181ffe941d589e927b8f835dd00d6e95e6321d43e94a50b8660b0ba13a042fe9149f363bfe31ef06143a2cd5c7dee9251f5655fd907e40552f23ac4c8591bc1e1e366cb511a42fe0fa403cbfb73c31bdd2a1e1359196a9035b2597157bec4fcba60e87b5ebdaa1d178bc8b25ca181f7f83937c8c3a201acad500b0c8c7a8c1baaa39cf9afc85165f99fc1ab40fd7a61db1771dd201eb397c19b5f9d726c44c074409e0aea734456aabb2d6a4efff7ab104499c65cc7456038d2e1e521f9d0bd62fe4f4d4ad389eb9f853a2333a13f58e47b9757e7846dde4adac938b42f687c3cbdab605f6d3a7d50164b2c9f37d77b59d886945bf855b3f6e9013888f290f56356bd85e950a76c1e31a1cc9d9f19393a53c57215d362b0f40da4f6003b01f247a6b1bf40be68f2bebefe748c93cf3d16c1ca47c85d4d82e7092cf42fb60a6e4295bd3e80a5a13586073ed88af95adc9ac4ea49bfb4b07e8ef17dc05a279701c67ad7d0282ac56540cc35f69db283b6b8203f0324f575f93b02a415fbd77fcefd05ffacc4e60024ba54dc5bd6af824fa8f629dc8c4f0798b8159f06fdd3f1746441a909ae9955076c5fa440843bac04341a0a3df6089308959131f31a1a5ff8c9827b4602200593853bf99e4826d1eb3670914abb897273b727181e77175518ee72a94e645a7286ca54739777db5e7fe50230766faf413df4e0b001fed890c423691ebc70249a425acfdf3e46e13dee851be09cf41311a9a0ea8b9bf5d61b682d8b48f6ade922c1096ab53575e2f227ccd97a9ac3df16d4e328b14db4a0ac3e0a4fdd1b4950279656edcad5bef36171f6c3f2f8c632f3b4cb92d84a37797bdd4347db20c00f689a5790f46547ea9338388c3adf7bcc3fd117fd04c36c437e6077db36ef687e38b5e1c0abb3127cca92fb94b19c271542a15e71958443384f8b042f69e58723f26a8d4e3e54ed8fa1bfaed30e28bca003308533a2d1161d3ab5b9cba7473561200e8744c9ff62f5c079329096d72109c4d53e2d11e7cf1f5e605aec4147241dca6cced824c9815c22cf03af5e4cf395636ae697e6531fa1bd098a10cdb46cc13259176321b8f2f41e89e94d9933586ee8fa90b8eb9b3ecbddfbdc6072c25a69ca2482725926041e69c2f501444ad805d8334db0549ebdbd995b8f53c12fcf6b2b560f390bde98668192b3a8fa89e287964bcd408e9992a315b6492cc1eb6b6ca057e72aa0c8277189ad486062f826c59f17fd65f772dd7b2615064b65b72dea2125a9566071db069bf0e61fb0ed0e4f06e7cca4066f867507677447c4227b76033545eb0bdc5a7523fcef1fa0505cf048b5deed34c050caba15f5859481f98b3e9a8f9ab69563ba906c4a4df8202b9d8f4294ca8203338aaedf6a9dc242a57d4b6f440fb8b6b5940ac4493858578c2549c99bce5e07a513e819a30c652b35bac26044b5a2f9222b143f5da2d122c36d5f89bb1ae9cc491807d2b5508071dd9df7035c5886c7180c3646a9eaf35c94ec054f805cb478131896605833bfd24378f363c39a9a4aae5fe97f1c37a9dd31ac38f011f837cc03117aee38112ce5f228e3c6ea5aaa95116055e7d2d1912969ae69f00533cf9ee7d8be5cd84a40019080e03663f75c3ee0e26ee8bf1473c380d9031ffd2a83158bd47cdf93a920c7814b784172d593191a4cf83ccb5aeefbd885e8cc7f4d219db412cba12034f439984d4a3eec6ebda7329dad00cb8fa5eaa44cb984d7605e7fd5363e449ce6a25877bad355458cd0cb2deefe32b8db927bb4c3c7e8ee811df784bf225fd53e8391c42851de888ec4734279cbbec54a2eb560d637a9845adfe23755796876afae98561;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h860a158cda1ba1191901eae421955269b0a1296dd5822ba1c91010b558a5c06da7f65903689b9aa05808326430a013dd4d94ae2a92edb8400a64429ac8c1a17c9344f179259de0bc2e6fef665aeaac88e3df2eb51db04cda4e87e32fd1f9e8923015f011c13ebbc299e17a7b93f56e75e9c24fbd3bcdc96e33bcd274e3e62b6d259ecaf8f599154d7e5c9630535e9c952cbf40976596a25d32aab6ea1a86826582ca34b390d4898afcddd78e1de393911d9bbab91b793f8b9065a4d4323bcff74257b0dcffd38a6aaae09cc00ef9d698a3cc046abccd8a2b71637cb5c6e9f770a39c57c0d65d6bcdec33702139a170a831f7ed934d54be42a45f002982d22c0c37c4442b313f08e7e2b9f5f97905cf2cd1cd9fcb0755cb9389a1e24ed43daafa4f76bbe26e6831f10427929c8fae5a148c869a1cf6a775aa95e0500a40f807419b1a5e7f527ae0ae4bc004f32ed35af9f5a641feea917e85db6566874ac6807191e383693ac0139e09e50ec74ee91446848624690442ce5e5a9948fe6552f94282f20cbf9dad19ae246d0fb82e9948334583472219539b60e195d3ade43820f55e4f451dd0aee95db7ee3aa6e96d1f2128e50ebe2f908400759b2444956e659201fe1b68df5880213775095f7765bf6985c3c9d2883ff0b84076239dcdb1215e2bd3f45a046c1fa43ac5b978ccb4b8ee1005f1cdbc091b1cca2695db70f2e8339d1da279cf77ed6b0d3a9b94b9bcfb00bccace089a301a14fd9fa320a1a99bfa92f2c714b2dc0b82f3c9d85aa058b64aefe10598a14379f1cd0b25cf9f32a66fae426909257103ccb96c62fd4850b8acf620f8ae5ca83f51b3640297c53f6d16479f0c2e47677b3e88c108f3bbc7cd235a0bb7397e967a3555311e0c657dc271dc15609d786b0acdc39ca0f3a779aba924f030fb3bca4521c7130bfc5a53c25f7408acf24e6eb506836051bcf5a55a0db5e25460f4e68c26917415d6d2f05f2e79830519b33ae402e14b0a92f74996ec546e19e7c3380dfe4d6a482179f8b738bab6538baa099472e7d59093f2c7ec05d31a51457c4c0eb5ca30604cf7e1f1cc093beae8130b2dc63349413fdec14d44c1a691d9e600a16e5bbf42009ceb53c98cdb7764a0e028bf949a973cb792cb49a5f36f1fec70470f6d0697b0c1a7ab52729f13a4180b96590d02dd0894a1de2e51403dca61c7b98cbbc366e3b6036f44cc410222ae6fb344e00ed58b24019da9fe5542cf6146344b13050b593c049144872092919646fe42ecbcf91ebd1a9e7250047e59b3c11ddeff3e3ddc4bd6e3a93c7cd57c5ddb906a13cef51929ac589782966ce4059675736c12b21171fc19fb67a4b83ac76ebf813db3655be46d6c805b9cb9c33d723caa8e2e31cb380612d2a5ba57c7d0609cf2758a85ffe9ed5a2716967c5fabb0a3c4a3a146d4532bb14548e719de5521d326e775742aaf6b4ced1dc1b14dd4eb2fa3139b8b1e033dff896d384f3eb3953d1ee6bcc6ee1d68b47ce04b20f3ad37a5ef51079aff54b2282142bc03c374c2024bdf3a30ebf1597a5829b6b0a090201704bcacba1bd76dc35672b2712c18bfee7997a5f6380d5a00064c37b8bf813e419dad65169dd008a90e770869fa00c32f55b77417cd9a72f0ba96b3c753a913bc502b66ba4ce67b700a180596aa028d0cfcef8286af9b7cc2b0b8ed09ece0507cf79de94fb571516045bcfacae3a3b31281f3d115436f803f1a00f89cfa835dadd0d61d59b9e6d79def73fa0ebb7f5566d4539554ec588b702ffb7b7d17d9616cce4f893ae063c9e7f64312c5f137b01861eb3fb1fbe434d1efb79ca062f4612d1e35d84dc802d91495f6ac47bbfbaf6c1478dc88aba1f286d72ac0166ca39314ee06bc83b4537ae1e2ca66562f268d60807ffda3057f9fc1acd0739293853a6e3fd9bfede1f01dd7db42119a17e0db1a7121a1a709b5c82870ba9f727e436527ee5c95dc27cfbbb64f85d34bc05f5982c740decf431d0e5b87310d5399038cb700043834465f6d3c3afd6da07941fc7a48a0fb304ca87c34d51b0a11dfe6f8a2bab68988367465d815f1464b860d06d8bb0f28e7c34c43ae55722e6d394aa977ae2bcef10260a630ecc37b6d3a26f944be054f274ad0146d47f67859ff259c65332ca7491f568669160af37c5b3892b3b117157cd83b3cb031750fa1754cb059e2e60d0e930c03d994067cbeef66302e1b9bdbf8d81c48931f2652917ffee959eb63018fe3a172314bf378667183422a2dca0ac05b2a0f231b7763ed19db2c859f93e16c2f8bc5946d69fe1a88aff0d1563a10998327980f0c61fa67967bdbab93b3f23144de1db73c82e41f5a02fa8fd432c698b015ea655f4ad667cf6e67eb4979d0df86c490bc748793c6ccbdc27c9ba763817f87a6fcc002552e895e340b8311f10a82e8da6cdd39fb78c8d04aefc8b20cd750051a17f0d875812a2c27033cbc2580bc623625050ddc56e38a5fd9e010ae8ad132d9c35c7ebf136f2e72a4ad769c029ce90fb6cd98a50e98175a9656902398c46665e629af30be977a2fb0ca5c3470710c2cc29d466dd6b7eefd0dcb1f39215e5bdacd5b8c7a0912246291e6bbc134ec78b3fc0ecd14f55a81256cb69dc5dedab99220e0e7e7dc656b760f63709439a24884012c1ca11dfee9a4a1fdd9a6c1c9fa95634be6a3398913e12c674e6ce90dfa6a35c97a3f9473234b149df86ea804a4a4f7c23513386a56e434ebc97bc37a748f5d320ca9c6acb716c4fbfc123159ba317d76dc846a8b1834a0c63b23e4328070af2ca9b5b87c0d1dde10a86642af3c15e39d8787f96b28a4d47b0fee88045d8e0a0256f8207449d1e149c736343b2a905790677cb5c8d4149fb56432756319ef6706d80193d4560f5df132ecb3307cd29d7089a450264e2efa8acd3e7c21867aa187c3805da0a1e5e6350149ce6ecf0480b6af46f71291de8185fc68b630dcb04e785e64307d22e9b02b0e64135b75afd32dcfee9fb0b35588cda87901efd8e9e14cb40492ab537fc6b231453c1fe5f4ad66059672631984d90ba1a01087d990dbcd7a1cc8dd0e19c5e0dde233a7b7e051d8f5f3ff512c95cb04f4e7205c15c08cb3d43a76325dd4c5e44177a4045a8337456be2be23518d81f231a3d4904044b8f9a983a9f83118e5882f21f4f9257c25cb39a7260f41d625db367338632ac11b9977270dafcddf91d5717459e15ae88146cea1a398feac459cac2adc34057ada242e5f27a3d8be42cc801486affd281281a3823588f4cce927a4a3beb9ee67ffa34c1a39d5b00e3f5733c9b4094904dae4c4fa1c39622f78f1e4f8cb9ae409cec288556533820c41aa7ec6a2f38f58aea59ef293400dde5c62b696b44683e5261345bedbc03b1a29357ca3c7f29a1e4e24ba3116bd9608e999650a610bfeae803561d6f9526e7e29ce9e954884ac237be0a1554bb177b40c2cf54705737e3b1d897a717c9eee74fc223851110e80d6a605ec7909dc58d4f8f84470bae1d77d7e8125b53af7d50dce46fe642e8dcce2030a7559bc099d360c8e8c03f5604ab45ebd1fe067573f21660f95b5999d556a95e6bafe74ffb3556867a3c0aa1ad63a0df7699f5eae1e4e98a013af6c1cab3227f03a5af4b5e8e162ef04cff1cc8aceab00b738f130ccf6005b6f01a2a8dba72f40ba358669e4d8f0c3ea4966555f3b0fb8e281ada4bb4530a11d247828ccd85be3911532d682aafee4cbfc4def8a240cc8f201ff0e4fddc7c85588b1c837e8ad6142da0df831ae8309750a4df2835d644b4fbbec78a5dd22a7bde17f574041f4390b0d72dd316f54156d92614b8a98136ee770fa0727f82c18efcfbdff001311d758e1fd555c457a815bac9ba1bebc596fa714bd77941c5b9fd65e3f520c0f6f5ef43f11eb660dc0591d97b2020612892edb9b24adc4c56fd13ce2dd587c883d73ae3aa0239ed3d0ba0eadcf13300f45b335901dbd6a475da5618fa3b5b26a5d124e86ae563811fd956e13c72639df944b6fafff09b62869d25d62fab1add69ff78eb256743fe1b17b00828f40f96d9f8380608e82b2f821f689d5bd1c00e61dd716ac9ad4b666dec72ba37c33726635ed2a0c58f95fcda062fc80d9f696a347fa7ddc68ef585ec72b9b432eb89fb90c76017c92be5b3fb12197d5a79402923645a0717047a9abf0c0a622432995ab8b06d6f62048edae8a8d4ab46213bb58ae12741b885bfaf89221510b0b8aeb84b90e92a6bf445d3d481aaf694b9fc8cdf793065136f7ce98966e26497e53690531b315cc0534a3fcc6855c68a8844465c7de9b61522f1648d6500ce5594305f497feeed06df5b22017dc313f2ec89ca554f08e5c6986f34bc37ff99bb3c92f964af45cc33b04a9038e4b3f222c0470279f2ef6ad3b48d28cc9055fbcab9c987d54d70d263a9bfaabea32838c6a2326df2e2f70fb2449b2aed7e8d9cd3a9bec2c88f9f06c81cde07ae676284bea9f7e64178e2dae552d4579ae984ecd9003b9ce9a8218bbfe39b33746c91fb6a8382c3ed7d1db32bc72d5895fe928e98f93d5e43bd169ed485c15670c6773274ed76e5590cfd06f11ba6a0b30fab7282da4051aa17eb5e89cbac33e7aa1db2b00c8c983c3bef3ec43767cfd913cf6652c14f0ae2ffb52da20bc3e5b43b581c128c5f9d65f78568991dec4c98653d884aecd1c9ffd6a46dbf7695e664b77cda7ea0a76959cacfc1777cf6e282c745e090ed200f56d92d4dcb4331c614344bdfaa045957f9eecc020915d798fc77d92be18869d51afae07659cd18600017a011b2cc0b8db71a0a16bf56952e4946cc16eaee589cf61f5a0729b12c51d7b73b7355c004956dfa590030002b0f876c3572ab4a3c85c059189ea0cd46c066c14fdc9fe628d6aca206cbed8590ea2f13c7554c297d56f0afc4d4acac506e59086accc16ad7b5c1383cdd66ccab089c1e69804d9325f82bde13e56903f658ba83cbb1aabc52fcf3e94fd84114d00aebc97bb23a5c000a3be1bcb164b56d7ac3fc32013e3b8d8bd89857ed067ecf4a383c2d934140e4c86e5eb3757cb13ae2a5040b7ca0611a1e6be1d3974c3d09abceaa9cedfa55d89e93b0830b0b597834ab21b8785beb5340ee9b3467fd1850a3c91f20c7a7f33fadc2a42a3a63abba8bdd419ced1c13d967688408510f6dabe82ca1b84b2f74d2dbea5ef796cd6575c286f423860549fb641e1a0cc29fd137e3a560c25ea40dda61b9f961e9b83f455a52e21978c4adbbcc140464524653d4385b451181ac70fc610e536b4cb3128314d9a898bcfce0fd4fe89f211321dc20c79c4f833d66349d6a6bf92bb1210b10e61f484f164df4570fcdca721eae739a849577fda708e6a47bf1607598d2b16ed95044c74dd58bbe21211dbcca6941da3cb2f5683cd8dd31b19f6819761d664f410bfadc2082ece7fb0e984910fb34ef6dc5ec5bc882ac39cacc4c4579ec91cfe673c17a29a85e3ca2e55da800eaf2f5cfd80ef556d2a7f3b9a70007da186a88c4a95d3946c52886e3b8456170c8fa6d32160f61e7508944915b5543d52000550a12c37c454b8e3d6c82c042e701bc732e27dc49409dd99d0e0185396e6b3aefca851101f785fa867ec5e79b0b1a2515894d70a3002fc269fbff44a888e49726084c437960b16b3127efa5674b4b7c14be42b1620da86335caf8b2ee4d98cf963b6287d284eee9e943bd8568e4d7a02b355ed92fa603d8148582098bf98354d71be1da213e1723171857a3c05392ac6d0057d7f2c655b150bc23ef;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h98e4b8e6c37c600011caf994b6a5810cbaf88bb5f05f9e5558ad7c9a2897ec9f5814ff03108b2e55332e5d94f3f3205cb271032d137c70575143b5c1cb8799c998edbaebe13729e57dc61c275ec11cfeba5094b0ceae1b7547a6786aa8866f08d4c6d8b911c769a9b545c7518e6ba40e85e71d4a0493565e77707f0d236763b9d5f5eb5031b7eff8238640bcbba15f7451cfe91a8aab65f86f8ffe69da536398da44838727cb8473fb690aca8f7f3ecf79c4afcdfb383694fc763cdb3e8fd4f5aeb4e7823010ed3619a00fefeb0625a50b9df1988983d6612929f4b115982d987bcdf81ccef64c819240603dcb554e4b107f2deedb577d1363b9e094b1cdd8ed6f35fd088f00b633cb7199f8f632f017d49b94448c48098a7fb28f3cb6875ec384e262fbaa0a7ff3dd812c29ad09cee561dcd033e869ba4a50a3af6efd7146108ac4cbda7c3e6c5c9be6fe912069c9e4e3e30e595846a1e996ff0325e415669e26849237ac61f15a1da5d8fbbd74aa66f666aa9dcf4d48f32d9e2247c314c7d4bb8023977518de2190124c9e30684b0d6a0b399d6eacf5913390c2b9c166dbb79015c9f59861453e2fd25635137e728a6b8de6e16cbcc43c5da4fa988a260620b26563b9d5a1d284846801b568c7b8efe7870607aacca4b4d24db506cecf574e6eea365708b9dd4a7727b3cd9ae41378e374900e54f9dba8714996a108f7eae3cff71e0dce37dd0bce3debda5e4950db10f9603e1bbca014fde9200fdf845ce706ce81281667380d7230d1a4b11a3124d8b78ab2e4a3544a0f3f9d68f2c44f3091c44c6bcfc1dd52c573b491b217607131ef52b5148182fe85048918c84e024f34f9cd44a69d99eb924b3cc6514e6a02ee06849e59eb559d98fe24c144624ac33aef332fdafac9e96c01618ef6d4bdae3261c163f4072577a23e8c6975a3ef69a4db080033229a0bec761ce6ab52e2ade0b9c52845228c83df9c0f678dcdf6828a567f4365f1d47bd98aaa59545cfb6653fed21a07dc13a911bf6609d99a4c5ac16ac36422c3395ad7e62f1da4e8d333e996601fa879cfb93845ca55aab07e8f4bc2c0ddd02205e8594b969ffeaa2ef69618a04510a6fbbc72cf3ab232ff5a032b95498752b7d4d7d63cbf2cc188f0b9a070874977ef39b17ef457203320a810ff9a9475ad86dd1d96485f23bf68c9d42c7362474176ce0b96652ef44b185c2249a212e613e2741125dddd80aea560ac3ef3ca7f331438e277394fd0fdd4b7290a36cb707d38ee1ead00d29e1504b9196e6d5b387eeffe73725b0dc44d12c638bbd6de13f5def1f3bfa5443eef789337197c000ea03964f5dcb768c7c2efb4fabbaf43225f2df3a049127acf5f04eda9153973d6d70a939b74326f7f1ccf6469a1b425f3841c9c650346cf2471816067d5189292c0c6ec1c4d65a65e4cec4f158cdc4b5b9dff8f47de926490e19a23147471913a314bcf1b72c54e4198463b8f80b0833416d62e4bb0546c05bab46399d5013712911ab6c1546f892955794a65997f1754bf3fc4ccf8849345fe7483c729b70434c1ff849558511199b688372e992370d786772e4342b08efe706fbab0f830b821d3f102da747ba44a502a1f7a9f53bc628848dcd43d392fd679da778f770613f0e815efedf9b4e51ae18dd1b96387fb0edcb8daab472e9db712b9af1c5bb97177b154fd84e6f2b9bfb8cd1b220e06855bfa78eadc5150a9a7e6d039d0cfb8fe2c6456424f9db599532caeb97e3abd31c84db812bf95f5c707240b1d9e97b13eb928e437b8b87f27a89e5db71c48aed6e82ec80bed88628772c0c41c58552bc95e1906f32827db80e087fcc2a1b2531859b1ded2ab13c5553b43c590a42f604bbf1da9382caa63e65c1ddb9d6f985a6d68f1619819956aa5616a2a2a558e8d0e9b84f408f1627629b46f35a90694a5b70faff46e41e98185be724acbdff8b5b70917b7ff3fcf6b692b48153d27b8fff9a244067e30eb9347f9ed5f59979b8fdf4427f42284665053867a408347dca37c67464da360d0888f55aa5a70afe7a23caeb94d544164fe8522fe7c2e23e20631749e55597df6d3be7d1287732481fb8e8db4b7696a7fb31a938077d4b425e4967e2bb77dfc40dff378e179ffeb29eb97350ed45dc5122bc4f168bc2e0cdaa0fbdd75d2d441550b4a3447e7f0149ce869ba9242f67419dec8f20316e1ebfa0b56376a85b7e1bb385a8e5250f03b4196bd2689beb7e3300cf09cf71b2a0c2583da33ba87780e85bded9f0a3c41b9adc56a8356af56c271cfe2e7950b88c27c859558e799944de90cc3f424f06715e4b81ff924a436fa603be5cb49489147cf931fdcb0ad2c4604362c0e8e9639ae841797fbef4e7af233d03530227b3fd15883cd8177541f8844b9ca78bf2a3100a46c14d8d21ca06cd4b0d9080ac154aa6b685fc3982bce5bf9c0a16205546553a8b869680021714011fbaeef759c2f5464da88625ffe1fb9ae0ef1d1d04239cf10fa9fee8a534f9f1de477e3d96681da9c79f0a4341883da0026a3d69c45f67ef02dabd02194b201445dffbe8305c5cef362d30d26c782587ff5eb821d3bbe60c139235af387c42e5d636b963ae4aa514975e432ae7f7567c78038766e91b0993f18c792fd239010711a33661a004ee0d95ffc51aa7b4a50077e072880eb65103f52c5f0f6e75d2cf1dc0ce62dae3f408de01c1ce462930c4dd0187e31b3513c746e90b502cbc65627e50382e3946d09fb04516aed38829e5e8d39b8277f8386a4a96d28e8e459239c96f4cb9890ce96dda049c0e1aaa758a9d08032a701fba2f03113f0eb04a87337e78ad36e4729bf31b106019e93b5e6da62a647564a2cb54e595a8fc2a6b5d33c31e0c7ddb1ba5d154e8a5494a2cea16627b5d5ec6fb063fe4fbc002c460a9c91005ed08a2e025e4aa2d5a086d470f5f4e023e0ac088b624f58734ad5801743c69f9c74cd417b030af66e7bad4ba97684d9caaf83b8a55d8c68dbc65b7f3ea9cbe6d216188b8bec8f4f27fd713148030598f43ae0e76e470f80e5b0fb5ed42872c5dd2d3f75ea04286ad54b32d6b4d268bbd66f96b5a57f55c20e3a2651ff7d47330ddecc13e198e61defd168de30c55cde36f3307b379453060f3c5da7f19d47346edcbbc01e4da36d4b646b2ade7eab4e287297f85cb45e462c37758abc33df45c3bc07b268fc087a6591b371e0925f4cbc13fd8b188b6777790623ebd23c066657b13f2c3cb9e920354cc069daf09d03778b0b312124b3c9716d59d47916f7da9b38ddf3d46bb9346ea60c5e8ac4bbc28b0a70fd3fd8cb58d6d37c52276320c7d5892bd4bb0b8540c1bbb7d3dd6d3480a7954e6d1c3dc41c379600e8c2e973b7ed3888a8c85521d825dbe81a49d7f663de4b6e6252365d72721f4bb2533a559668199d7033735a810f932710cedc32e158401347d3dc7936e3b8d80f3cca3b4cf9388b37dd08404ec98638da023c6c7ecf15b71fdd5b63ab5b2a0b4d1f7f579352d910324283612e4032eea74a67b2bc47529e6634f64412144c3353f13fcafdc165cba1b9a493d85eba5dddef2cdb86fa758b4d85b28cc1b3205971043a231ecf1346aa645becdfa6441233c5130aed2ad2dd21ffb45c101d053716a695119dc9df54e65eb52a54f59e3809a8cab9ae584d714d26fbaa4f252d5683e972c8ca121b2ee239940acd8dc6a42c4c3034b423f5b1f19e13be4dad8675b7f1854bb143c7fc93ed6040a43f1ddc41693e37332d88f97a83c23f7eacfca3d4dbed1e60d9fcf1d74e8c51f5212ac947a10a55224d1bd07ef76bca6fed26aa1d69cdde9e91ec3df3ace7159a0557b96ba3de33e02efea50a6d401c59d7771e1dd1ec8eff8932048727d821f89e68be47799bcb44f788207021ed3dfa0d839aa00d83579e92c861e05a89babdc0ed98f72b8c5ed27cfce587124a028487b55275a986503ec562396034d455e979d9d49462d3a13b745cd18fcd8be3ce51de52c3f2b4d5824cb105b2766b3c231e26889616106f1f8a5e70bc18b0b3965330edb5f180cb850e0459e64ec4bc07817523bf4088c8e32f3a947f641c8bca870f322c6c89ba90197ea3f3b1a507f286ff4414d70bc39b54c4830677f71fe2a531109a27467158a46182c3c7dcfefe198540eae17d0d46342ddf0ae78b2bf1f02c1aab27799fb851bb67962f37f40cd183b081341ea06ac67adf1749272bd2b3e2260e6395db0f5e45c3f3fd0e73e4933ac2589ddd364fafb7cbc1925eedfc338516c8bf2ce86e08ea882b354e914fe465828174554ea089c48371d99a2bfcd050cb2b39543f13a754120c20bdd4530724a460439e12d69c2284c3967ff3065473e26fce0bc30666f488ca66acffed856f16ddcaec1c1632c3a9790426e266d4ae7930a1488bbd61270c6e21fa15d735db700e454591b94041c31a386c29eaa87d5d34a601d6a3f82a4c28e2aa97bfb1fc32d4f8c9439a9b2a43390d562c0a0eb3243b1d434c20a00afc27815b9abd4e452e0de7a672f65c77664a2ed98296d0794cc5c5abeef3372b3ef3a6925799e18f2f72f2b24259b49cba8414edc0fcdb93f3ae7e2bc73ce30e230cd91d8c96548b89b02a267e6fb539934caa599f7e5fb70a4e122ba560bb1ed08144e278a8bfca96ef32b905ca230d213a52c3fffc2e59289383bc48aeaf3e55499b781d0757b4a3a9250bf1acbed40882dc71c24eac16f34ff2963f7b94b25f04dce262dd774427318234dadb391af24a98937bc0a3585a056d05741649827013dc331e80c137547628e8b9d599053a0e8ec87a25f821ba404374032cc1cd0c9658b5107c482caa4914a2bce124f7efcd470000b9e5876482090482196828e48e27d82280ebde4a12adb040d2913641fdf69c5640162e2f4e1728163d84c60bae2383491dddd8ce370d4dc04b58aceca367d6f6165104226fc6ae1ecbea686d012aaa1154dd79e9b7c1cd59c5def1f52227cff40ee5d4969bd3e6369108bda46eba18077145b6b2e903bd335feb635cf441ee5c8f64fc6e8a1da2084c727b12112b569160b534d281fa1f8ee1464b50069f6e597b68d136e80e373657ca33dbba511fb59ae36990c759f3184b9740cc5e3dae7428ad5bd23ec8354194152e9126cf54bf0d67fb470ec2e9819f8ca6bc2492403a7ecb5f3ba4ca949c4aa884bbd0a2ea6b0999f0ecf7bc83442f9f5be0caada682e3c91755a0b226a2867ea2f5b0d23fa1ad88c52b7c43c67dc3d5e725dde2fdc3819d1b99e903983e136b04d2487f212672a40c7a316d14996eef48a1163e4ecf7d267f4c63a0b83ed67ca07d4565e10a84a50a46a4b5afd100af37fc8fc920bed8d2c8f16b9b13dd4b28666921a4542ff2032c8f1814281c30da16d2996c016ff7b89dad6528aa9467ac690f34572446994d686a09514504c93a569d36871d702d201ff81e445b3edbd532ed50785879a0b7a63ebcdd9f0c6e83c29bf66342a119116bcdebc84c18c49062bb3937a53bf0c1a05a272be71b1184595e0ff1f0d8b2730852ddd2b4dff8eea4b2d05565ee9b07d8591273579a484b026e95cad5c9877e12e57e60576d55e4c63210d3a3eb995086eccfc09542354c2d53ae15f3c8a00bfc778f392d53c523162322ef08d9c840d691c01b51da230a1ac4d020e74c2c5e0c00b0ed6b9ab3df0982350f6e45acb86a2f35f821c1501e585a4fb5986cc8fc51ef70d6d14cf45975e842c05152de2aa481317887c9b5e7c8c3824c6bdfb5dd075824be39dbf87d90f8d786cc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha8e2659297f6d74f3df27055e445592da59f74d25650f82d7bc2dd6bfd858922e09d12eef851ebddf42b4def93d5adad14d8d1216fde544cb840803b8aace55f3e7b7ca73e26a0e6113c43623147f4f6892b87d987b556df983cb4973567e969454d915b0272821ef983d56c07524f4a48ba164a1dbe12f69c668229d661bdec0f2ba17646cfb86336b037f041b64bdb7eb1a4ed8a290e1d9ecd3c2df0eb4f11d30bec4713f851c6dc77c8f7a6c2d1ba2a8a8b224bf5db7bee0df6ee85678e9374238af54e7da0b615ec2b12375df0c32cc0ef04d4243051de739aed2287d37a2bc389b83de1b80d50330e125ac3519c7756143d1e55c537de62f68646d4d5ad7fbd7a34e20e798a1af6bae3233137398ad1ed9e9415b1e63955ddce65ec29ade696470913e54f893cfc395052ef09da05247377b7070fe1e185179debb727c81cf5e89f17cc77501c6e2b1a38c332018dd1cb40187562c2c2bcc570c9833ff6a779e90b78f96731c6b05539d6c2a7be336ce3897986f61e35456114845fc805a4a0a72f3a647f7748c3bb8068e58577545f48410e6357f78e7845195c92968a0c17655db6942a0b51992344461ee9ab628d1b4e6498719166804e206947fa05bd24c1cd31e2d81ec990f86835792c2ed7761828071f41f692fa5f8d385402aac5465d4c946d5b7f1f6f16dc905113a56b101961d92abdc861c16894f0cbc4f218166ae3349086935e8211eb05814dd7dad16f3b09bab14e1968f01969034f5d18601e7215721bba6a8448375bd3581429199684876733ea84739a78e28ea3be1cb5647b613390ef7528df3827de8feaf4c7c19222178a4bb51e8c37787ef461bceb8d5d95c684ea56cd0020bc709af65be9647c84162eb4c6a3d9f5ddc81c7ace335bfdedcc8414f3e14a3bdae9a3daf444ab6f4e2bdc0956c176c39aaf3e675b58942b445c6567ffacb9094c6e3a08341c7c84276c94e80b70525224d053d10dcbbabd3d053754dc3af60a4442e072f5129cfcd501fc3807cdde08b467c2db0875998412833ac96c7f9eeeab430895950af8f491e36f84b28cdbfc104eae6b05c345d25243fa8e595cb0fc0936c53e425efb5e3b4dd3b2f0a307696e65612861465df8e02f8e924091d52fb07191714eaecd504bb910026b4db8cbcdb1de23c7da0cb2e517215d92776e4fc123d38ccb9b0c6a88da5532faf6ef3a490444ae6129cf7fa92b2b4f6ec8e040c187503a770fbdc89cf10e4a81706946c4aa060aba6a3bb2371e65290d4b650b883d5db0dbfbbc7574354b59216bca1085d88ef62d5c883393504021a07e38b1e612ce1bd24fca53b57c7567a32d6283ffd426c0a4f39778b99ab3124a83499ebe3be2c79ad8f57c2ca2c471d46885d536dc846376bddaf8358ad64c87ca726fb608da7b79e015b9be0ad0e6b17405ac07375ba086761d181aacdc6ee219df1b1ea2805bc9e7ecf8798fd372ff62ce818d7da1d40369b698fb056b74343268a5fc9e9cfc59235961ece69b2fbe3d98d9fe66d230799d8650bcb6163ba045fb289d573ecc86cb7322239a85331bc2db204a920e776547bca65c7707bdf97e697e10e8833b23a29f2a296540afbc4e2568c8f6109d3a11ceb7a2d4b72d47b8bf73df6f5a1b2f3b617705060517c510fe585587888894270d3d842d3421d8afc7e4665c39cecba88118c3a4781b7e2992c7ded015f07df6c329e81497cf89723c8bdbcbd37cc939551d2a1ea2de95aae30f9c2043960bfb6de37c027d4977368220c014b12f59c92cb99030194502983de314f5766b1dc37d72ecd83e3820648b7f33bda9160bbbe4b6e5f3fc76ab4cf173b0235c4ff645e151c6c80121e4f62410fb4fb3cf98e0abb85def75e4683a18fe73d1ddbbd1dae2813f0fee1cf9073f0a9cfab2d0385d0bd66f4ddf0207e2f74579ed13a8efa5668e429502ce21f78cb4a59cfc8086e1abc9bbecde3a5953fb0e0515ca16deb4ee872fe3b615d53825ce6d2aa80f3ed5ad6f69d2f0b25422169c6048ed60ddfab95066fbbec5443ac71f6a86243f0bec57de9b77c842c87eaaa9448180ed8b7b2a39417b8e95b698453b44380a4a63dee4b67e259bbdf6ef6b053e111885b9f18349df9b6ddad10bbab2751d091d24016c71b4a25f6b8ccc043fc60b1b34a87c27bbfd7849898914d63f8f4e4f763f67d1096d9c85e9874afa178cd04cf4124fe822b27afdd718982310c7c49498c413c7245530688c4c6a4c0d3c1969d28e7346d1f70a1b8e1d7a792d15a4aac716175c00650ecc0a211e3239f656dc4e27a8ddffeea5a94214e458cd736024a4cd78b719bd2be78be5dce114b894cc30c1158998aab080290ac90c7ec01f4341e49726a52fd40ed5f6492950b3462861b99bd92fc70f87f498466b76e72dfbafdddf207b0fbbf99507c2226885258b38c1b579981f708ec6df441398c01548986348a500a6e3e78fa91f5d11a17f19ce4c1746c9c42f9da6710dc576e5c535964d9a24ef4ae822c11089ad16f5b41a93ee8dd98f7bf97ad19633236b7d3aa3b0984514da7d1c8dc183843886c9dd174273de5780520c4a4d1df5649c2a7bcf19ceec46d2f95897b0cffbe0457e6096e13a5bdd657f38eaaf0e513e46cc873eab4b9b429ee3f9bcbea2b544273d4ce38fd37c478ba8044759513f864bdece41676005baaeba734eeede34129e5dd3d1ae5294fe9bfe526424f0ec58aa3c5e2b53eefad4e629beb30ad67d7bec4747c0295d4bfb05bc43afbd962e77c45aa32cf2a42f6cadb790fdc6690fa67d04e497f4aa310be575458e9d73f3db2eb79ab9c94226964dcf964bf26a73a9e0389a8d4aa4445c3b9156c16aa14676855f816305de6eb6fc859faf43b941412238c7e36305479cec113615e69e25213b08133fd6cdf61544aff4d5aa0a55e56a3419605a04e53216dc8a2397a7ec16cd0b98928e3e40901c23f32ccf17e595cb007c2adb479e8bb7b291481e3707cb13d6afed70da3e319fb6c22a532ce49d62c430e38f05c6b75d677e5dbc9639b7074f1e5a449e3a5de53ecbe41d5f17d78fc30aeaefd7eb307760bb90906f3cf6c9d6b57ca8d415c5831c61ffb6543941001df1a396e297bbba129e2af9e222a6e9e5775f8c79b33d7c5d12390b8f5463131efef51d8a6a348be9d254af561e6570e0fe05fa4180309c4ed123d9257567a55037bcf7ba720e9b7658f870d70a71075b84f5fe61ed2c5f1b9cd8f23dffe7bc0c8625661a113a11d518e67edd8f33e09e9e40d291f860697d46df3c0c1d061c223117a7ff6ba8bdf9c89ee61eb587ceca4d489da04346e3f61ecc37dfdafc86797285774bf27076d6e0fde24c5f3baddcb95ca9da5317f3a5d12671dbcb4920ecf8981783dbf0a25d169ea80e9aae1252067830433a393685eab7d1d89acadd52d7f8fc7b5db8e316125822d7a3426eb03f8f04c6d16589504056c64c1afba263df1b03c0ba0468a7bf98bb77fe61081116d1b6d640f55c6c67ca914fdca5b39ea9b512e3511234fa329576a5c87c0cb53f78255647f2b9584f32cf90f8637617ae8e541ec0d8a2031208ffe306cdf2ff5f879308b59a527a0aa33c78f28ebb94b5294cfbff8527d1ca3789e902c211bdafd7771a46e4c9323e2d62faa378735b2e882938f7df3ab64a6d4201e625264c2545081b5b2f7c313082a666ffcc7ecb4fd0df6c1347b5e1707c54fcb0626096a69c3d2c516fbe0e0a34d4f353f0c3ed0497fd6881dc901ccd23d818f6c0856b87082174008f625fdd048055a29f0fd0bd48e7bfd1d5078276bc77bef9cda4f947ac1e60de117a160a4cb2594e96b49f69855b9e8336dd0cb04a7d2d2b2176598b6be1cebf449e0add5ea8229fbfbeae6aa0acfb0ad9a2216a135955bf9d3c216eee5c3d9325caf8d2e1c4b14b37e11500c9aac0a9432e6818febdcdc13ba90aa6d8dc8297accc1121322489d8d71324d7567ec0aeeb4a64e9490bcf54f46ee7b98aba66f9afa8a87b97b30b12bea0eab3a1c082c704abd1bb3c444df8e57adac06d2a95a09b81f133464847e1d6034eb3dd431d5ef9289f0a4437cd58500baaeb820ad3746d9083649c70cbe86befc0c1a639f7e703a50c349177ae25063167ab3eae7cb1232d4d42c77c437f49607235e34a8fada3a56e625f22fcffd92475147f09ce85381ea105c163bf554db8bc3cc5e8d94a2cea096503d50d9bddb0b6594e7a53c77a33f03a4c8ece60c00bf3efa03cf7368617e019e89dc5d00c32707c5ff61fba77f24eddead4f97f3047a30ff6b9b6eef9bc141ff4159baabbd4bcbabeb1ca78d7b72b0d098ed60d52832b8f8b55f31b5411101cca8b3816ef507c28095d1c76236a6c80c6ab148046bde5b28f050dc560a52bba154e967be252a723cabb9aa3d09109bdb5fab2188371ef1981fc8da4d307d5a04fe1b465f2c188e008d6371d1a31db4968a654f3f7dbfdeb8341a7cf7d53441bc5c39e6ccb93442b8fb768b6f3c201354cda98d59e8bcdad9d3bbc047c218e47a118ea42d7bbe9ed3aae907d94d65ed49d147392299bf9cb18b82bd954aa82ec8adb850df78ee26d074f770d5800e9625b6dfadca4ccfd9cb0af12d77d08ce581c12eb88cf93a47e6dfe2d67149bec1f53ebbe87f19f07e824f271014eebaa874752f2a37042652c7a5f54c41a82e0086c8727a999e602f1b19ce872d81a450a1a1a057fbafa171082fee601d7036b3fa9093449c82750cb71173a1aeb9e467aec1ecb934bbb0e041e784f10bce2b841a669b7c00d7e6364fae70b36178756e2c494f4ed4919cf90b58b5bf7ec29b7db947ff99f47a5a088c6656d74a0e4882118985a511dcfe7b6ef9f9e26180c6b24ae09edac11248f878efcc9bcc3e5ed589cb9b4484e87fc4e53be2f05fa5ae9f8f1c238c6e99148a211bc32199d16c18c3cbd0f802f272ebd0a18e666492d624b5e8212de81ce62670b8956b30485c6f117ded018441571d8fb84c45d52887fc56f8b47f77075b58d2d536d96a8439e0824061e013ad8cacf617b4b86880c778aced67b84b11795a1464b0807afa5716e0395ccf9077585081928b613a77a0e9619fa983a2100c028e3bc3c560c880603320bbd466f256d1d1df503cf65e4a447ada28fd079515816efd4c0b562eea72121cee54cf5bfb690436e586e81e9075efc96ce9e4e0a84a46a823689baee0a56327e339d87b0061c62f879907ab21ed3a75ab57e15e154381710a32ba7ffc93030a5fbfe8855e327836983938e1de81c5f186c6207a4ed178f6a7b856f37078cabe63546ef107de53cb57ac6afb8f6fd2dc8c0303f3e61b99e738e14238621263758f0ebac5567862e85eafb4487a2df394ba0d2b56b5a3290bdce837434cc5d5441067d402b15edba2cd12057544e3a60591654bdf6cb3bd6aa339d2da15a8e56efe33ddc623d888d074cae6b949a0db8a7dd9cb74b57cc729107fde572298a67daa5e2733094e94f56e8bff20686a03fed558639535758d17ba0be4249ee8690e9fcf26a12893d28ad90c6fef2d1a572e82af9128f12fcaf6debda42f5e0fc567dbf744d124690e42ac078da27c9307b15e04fb97c0743c482c039e756cd1d07647d772762ac44fdc14f1fb8950b256f6fdcb77347b0084c984a72359557bb9dcad8bfc6ece55670b7c98e0a9e4c652fdfb5e3c48a9c2d5155b58be124e481fcf9e26db19925c2f0aa9031b91d601adc242939fc331ad03630f0b41ea637323d22684bf65b7dbb2dccff61d20ad649b5c9ebdcf7a3213acb81;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb6e5a5ad15d50985cf066411789aed123c27400df3e839c2f77140e348e7b15c267ea37e2305a9e1c29d88b97c88e622bbb1df1e7389829acf954a95a2812ec2ee830908e5663830d6720625ec2669977a973c4880e7ceb1d7e335cb8df25fd1389c5f9c9881fd25b738e5df66228cea17a067d2e608d8d6fb301ad179d9c232ddf7d5efb72c65b478e98c22d58544b42f003b5589fed4cfcd8517944ee203dcd55832430402c52dbad76e2b07e7da70e1dba21cf0d31ca082146b86a6f0c7fbd03535cb4c201384526dd87e16050deb542cba1258ce6d9632988c4721722950fcab7aad8c4874d7f2c9a9ed4c2cc2600e4410139c3d307320fc4b85e5e64c303a8b07ee76344adc27d904eda2477b054e426fc58d6cee1afedb784050a124d47092f8062180fa6ffa1a950300e409d6b6ca61d61a9c5591e1a846307703a8eb8245549050241464538c7515036be010d1b3c7ad236f123b29e5322a9208cb69eb495248f84572f72af523c4fd6483647849e69f7caf52d7f6b2017369a4b1df55c362a8845f4ea13b503fd1d018505ed7faa4bb15caafdc1258b86e7524de70eef3691d9951e6f568b44866c3f44b8c87d189e29a9f495898c77395bd1502590dbf1d8277e97e51429e4d7cb1d8d9e96c9f337d8394bd5b88afb6dc3a7b0d2599af6cfe93d88c0898b9bcb3843e1884b17e2269f70cdf84eaa327eea46f8e83ed15ed0adb5bdfbf657f196dd16f006c7b2a8b3b6d185925ed42185f1a3be0af094f097c6c3a4514d13a828d4ba774b4301f644d1b3e82b6fde269d17225fe24d11c8e98c6b77275339c9e45b0fdbea0b26d639706ca5025afb0a71184527bf3d374c603626a2797dd02a5fe2ad253bf05df25d04ce33df8afa8fbd5f575067af501190fa80e7d021560545c473b3e0b1264d3396384bba49a2bb5fd1c82bec22cd29cb4f4fd59f2cd16d2734ac22fda9fd3ed770887f6e49ac8f5d4db0a3d5523369ef9906c5f31b07482cec786e115dcaeae2ecb4b50144241d3d4b49c061c1377ac6f2e29ebbefc8d7381d8a5d7b10be4987cc7e8840ed6306c7b60d7d96a6a2c135d5547edc0463a8b47b36b7c7fa1f0d63ae5297f47c423850946f5dad4bfe7cb74cac6ab9357953947ec1a4963971ee903702e2906004a85c22317602f5993847abe9ae39e94fcece289c1acd05d0faa8b6bc6f9d7977ff844a7e939c8bca645a0df4c0a2c753b141a4c2d5113203397ca0cce03163ea66ac219bdb0c3ca2a16f8a8d7764675d845e8aeee312b8ad0c6572f82e9292ad1dd52093de722abfe6b1e4e5d56cb8239de72dc59ff894b1583ab2684cc11370d0bacde1bf3d3a3e0c426d08ba42bd9ef7a628ef1a9bb778cbee62f255c2893a4a3f23d0c35afc18866b0505ab93a750be213ed376a9d38353538b5ab51823e361971109f03b0c486389db3b8802b9a3599179f761df8219e0793c4c3f7abfc6a31de89df08fee14bfda94296058e84bffea45f2daedc604c678299fcaa2c1ae58587b1899eafb21a0960a470dbf8b9b861e47f34c63191b985547e2a6903de3c2cb31ab471d5f038c11caf1624754fde9995da66c120eeb8d070d341dac960fa84dbb08654564f60a8a08b7be4fc2dc95a0f5c1b2c5e61ad442a751f7bb7f3257d2c3b0db02b984b240564ec20090c07480aabd2bb866f09b575077e67deb8486c7e48fcc8f0f0c96021bee7e914533a4e40b2d72d9e366115742fdc43f7ecc6232f2acc3312cdaf579bac833a297eb1ba4aac03b85f7997b81379d0ecdfe350fd442cb563cd7e8ee49e2666619c7077a644a5ce0736fced6cbfc89a9619815d6c1233ceba87b777a4d40ce14d7a13b9b97d19ea016e2627302c83dbeeeb7161fd742ea69958388dd9e7db4884b4b9d04faa1b53df9b8438ca8311d8640d76efcba1723d6922ea5f5eba99313a17e1738de923638dc1cfcf55e51fee7390ae6fdf2731163af9e1d6c4f8eed4b76ccbc89dcf70eb2645a8a80f69f163edc7b1c472c3df9746645dc90f44ef7cbf410fff8b65588a87c04733e56f2d865072f313b16d74b6cd60783844322c003259c9f0d73b0e31a3834985b4b41964e9d0df30aaf84f7b577774ef6a2f60160cdd63979240146e7972d7cb0de65a6ab5081f14a7afbe8b4d462b492b0570d7bca9954230339e07b8faf6eec92ed4c979dc0318cdc1c31b5df20f5521c1aec224ad6172dcb13c8672f61d86e47cc1f83d8021d9be526ef0547a286484fa1dab08a13ad26fff73dfbaa6afa76e64f6463eaa34955669350ec9017917d7d1867f97140a5ca35b39677c95c9a91e327d72eccb5184857b62a12d6c759607c6c669b507c383ceaefc4ce9046cbc463bd71472058f83ce9e40460f90d22ae33083345536cb6ecc0954e57d7a625a5dfe19d7d4f249a34e87d1cee92e5f5ec7cf95072d6ec6d269d48551040e3ed82a0dc9cc0f2d3fa67f94beb51bd7e1277dd99374feb8d8aca2dcb32a116bb05bc1362b45335c59dddc748e00058e7c04cda273f316d71c8b72cb5d0df7b345a0a1e5a4e6be09fbbce92afe145581b658dea2026a92b4bf977187b006db3c5faa5839ae3dfdc094d6415407d6e4975017f143c9ab217b3df1d4dc45b1cd56941a76000801978d1a6aa79c6ef108a0de39fde76024c17b12cb611b8042e8513979c6d884f0bf1774bb0325bebcbde85231d9b9c2f67b9d08a6f4476fdedcf599e4d95a24b17a955cecf0cf695c4c092e86abf71c6a1ae7c8878d90cf4e51363c7bacc9b19927d8181e97dbbd53020a0466ee8c2f8f378e5722c7c74fef6fa51cbbf5b198e05c71fa183c82bbf614f7dc9cf4a5c1c52c4c83f72b73b5a949deaf38fe1ab2445f6ade065871e22db76dca025b1318d256806c3978a7b5b74ceccbdf5715dd7af6b7f15bcaf76d5e17dae1dcbe55aeb6295abd8e6dea28ea01a0d5c938303e6887211bf28c3151ff87b549da80bc2acc479a2729c2734422578c2457392bffbb7d1a0bd69f10150ad077eecc1ceff6cd718ac874ea1fa8cf754b12f813cc90f21cdaca87e185b47d4a0544e14e15917721009421ef7946344c47ddd05fa694dd8515a7ed008a019d7cc2eeb787a7c156985bba4a9b0dd52c3640312a5beb396e8d6958a0bf999efd1e99ee11a0295f5a117de6a34791a996d9261f762e16b4ac6d4ac3a600b2961251657e9d9f9484ee48353cdf6ba6c4debb81ad32227397706826419df88742c01d9785c8d334ef1d902f815cf7a4793da50ee2afcae36e62dac9be005c1d11e2b64414666bdf6449e4514447e9f28a36793894aa8e22a4ede704f09fdce85b7d2b346f3aab92f5f441265db8a37678476c7c7a9617abcf2c9f65cec0927cf06b032b9101b76a2c5875b6a746862400be0d8908814fd5d58aaac7563544495f8312be5f820a45683d8fdf2381b3941509de8af784b38833b7f7cf720ead4676ef2a02fb28232972de72f5a767a77091bbdcb62e86dfcb639a52b34ee747d9f5d3d065364985ab677192cf485d03a4091e7e91c9e7e3ce4b03f33bcc3fd82b065704470e141a22a4eccb574b173d3f91c31611d736b8997c2e84c5eeb8d7544d7af32ff7b51921c8e1a28b3ac465b4b70ba4ee67e94862d8404d0c795b21ae530285370336819cec8e62cdc1d15665eb9f99b073b4653cbb972f4148560da0dde1b61470d7a2069a9207b395abb26c51ba30472d5b1cebce983922dd67b1bea7e2dde510380b70e9ea9add4f92eba308798a79938ae72ef6555f65dd56b4df6a51e3d834ddfe5feba6ae2f0f3c7566d52a1ca23f40b2b53d6878d2e305f7247e84faf97ba1b6c9221a3615a45443254563b6b719822f58dc81241c8343e1993c198203b331e2f1b85220f23aeb924f777260aca30ca66b61a525e00eddf56098cad48184b66059363567bc7ce0b113998f63317ff0589b2e0b334c87ab678ca5076300e433b9309541cea4f8ad6eb199a46b8456807191eabb0120287916086d5de4cc5d67da68c0be26b2f4f25f4228d982ed2af1960fdb6347661201874e2fdd28d73730b49abfbdb58942fa29b4e74047b3679f36b779aaba3c4d95463fcbac50a388e59820f1e9adf11e6feb243c77e3f7e377819489a8d4cdc333d06c593cb114ceb8baca30625758939952d0a5e52a8e1f526cece096096d1a279bbe76138a9818c4b3e9234dad2fb7f2feb1a1591144f10db8ec1f558dd986d3e1c8b9ebf72006cc39fe289881738baf8ecb6d24929cdba4124c548773279e5eb3dbef3077600df7e615e2b8b306ff8c580745681067a604dd187d6370b01049a3cdf1dc59dfae66a9849faa4c9e8f349495d4b4fb4b6bf82ed3ab60f28b6ccf73ad2ee75ffe420e0ea17fb19dab3793260b299a7fc78e27d483756e253eff13d27a8e686de73b3fa8d73bce640b61b1acdef44d690b0c9b60bed2c81d440bacf8e459ab5ada224d260bdd54aed1e57de7caa644a3141a9d6bc37e6cc6da950459cf988297d8444b7d67cecb88792dc4ec16fb7c356cb488d2a01bbbed6b446174f5f90172b9786aeec1aede2dcedab2e6919ff70841d58c0aff83d97a3837dd52ee07398f716d0021712d234076b1144ffb94ae26a9f7e9e682a5c51a9bfde89d3c368c1428480693a50dac1f2f548bb1057e1cd587e5eba3583e4e1d518d4c825dd9c490eca97b407c0ba7e3f50b799650ad968805005c845070fea3d0f23f8c230a7d44c94c96d3ba253378e5f9954f79caef0133c963e666419077c3731ae36265b9a156387956c32be54c923ed6b424dc260ac03728af1501b7c3f2e12bff75840a2d9bbe5143b6af9e7bb72bfb2318dd865f646ebfd3630d16e0845d7110af6b0693117716e2ed656ccb417d7a895a4eb26b9273f72fe2bf5f822f3e86f9318951c76b61a13b3046e8d2681e9f0010d8406dd79e8b2d2779374cccfadf654eb1213012996990af0750c0b7bcb0cc9b066c52dcdc7c4ba4705a335c08db9852d703e3f88c0647cbd460ed7435dfe5dfe78a6d59a0c71e88e5d057d0cc92f2a8914d2f270ffd73123531e6c857ba920d0ffecd8fd95c257c25833e458b64a32aa4bd0b5a17341916e7f252c365f858c595071d283604028cfa13be3cca8d2c20f53b8181c68cb62419ea3f49e42252e34c227a9ca97a42d9656ecf79ba6abe4c41c80b6dfb27ae3d7745db8db1935a3fd8ff05f2f7bbe551c4066796b280b65c435635f6e0de7c3d2766c1227bbc165425223bcdd4530a89a074e0580ee6d1c7023a8eac36db315f5acb64a6df17361d65c4c290caade9ad60c959b40796ede711ee08a5409778adba065b57905e635636becac8f73eb5b60b23736ba0adc7f911ba50640c7c90d5170110973b0e02b46236198d0078db7fc484870ed9b656c8b6b464ad6bd54db01d66cd128daa6144703f8ad4bec9e7280034df1f489af178bff35bfdb313df26a43a60ad626b8a5d6e0b8cdd07696d9172d7cb31c4d0bba97115dbd48c047f1a1f7ff3030b7cf115e5c95eb98a3ebd1655f56a89f9fd7d87b309dafbaa6f2dad3bb6d290d10b7e1cb6a5860ab903c1edb81304c814616c849bfc6e43fa55b712a910919f17274e5223739b1b08552273095f95756548aec74f362f8a3d302420544d0e228718da8198aead909f855abed5faee13dae2e4aeb4c14917a6068c7edce6e3a1c3f2958bfd126028bd878d63eeba0c1d5a053091502058ac53dc2b3d5341c88ff6572fcb42e144a01694370c5945ed027c0ca2d32e981fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9888aeafd15dc59f5f970b49b56935480cb0d744b5a7832be8fbb486f47d1d7dc9a69dad775a30bab1ff7df50484ba9bcb5e4cd5da67678624781c889d85ad98cc1170b54dfda9424b21d9f1237b99b1621ff760e44434c5d8206fddef4d45f53e18d8ec89df76ad7b3cb3ae60aceac1581cd9a7be02b4004eeb844d73bab29dc50e646f6a25ccdbf15f21e12da987d1e82e8f1396a77db005a371551455bdfbb9d7d384805dbeed5847b39d552a3da8819a32157f4bbd999ea5a0b24c4a8a7cca7d463d638c681f6e0352e1d9e63f8f1a90be6ecaad4de515d55a0af22a3c165567881d028ea5defe50d09c59c6540b3428b55394a19a1fc5259f5b7e7dc721286d7e3df614779de1e532daa1a847824331938bb0818ab37f6592af572a4dd49251d83329c4b03e0326c6851d497dcc9d449416e772d7b7f5b1f83b0fecdece08fa206dcaa38e48edb9c4819e2e5a3ea63b68418c1b8e59302fc6b8243fe6f5e13940b80fd693619d0b10c9825ed70875bbde0735c2c758c16b73c546194b28bf5f84901f5161b2025c93479d51fdbc52bcb5e9f233db213648ae424557551d407ee67de05d1fbbb7089764257440adc82304df486993cf1adac3b1d16f86ca3745c68b172bb7357371671d5b74f59cc4f0542ef9065126a75e2974da464c19a0dd688d8a87068d8f09af1cce6ac09e7c50903cd25a30e49bd49ca49176b80d1df1ee90ebd890a0babbc0585d4238fe418ca0763abba69a0732782e66feca0dda945f8153add5e2044e758d339c337c5d23fba29da9993f76e06c46ce9677ac4b2b6588f4fe4c2f09f312ea914a6524dd64a21aa982a31d7f20877c3777e130f987c584427bddc5949346d9bd37653464f5773c1450f750e563bb3afe2862985ca8a99b813080966bf454358941c599d9d478b7ebee3003f881be461eb6feb0bd8b76bdc00184a5a4f05e87c853279ead77322ac7dcd51ede57f1a85e4b8e32313f7d613e60047344c4e4df863c912ebdc0e4306535c72873bb76af4f8d289bdc879a48de676da0674567ecd04e2ee27c9aa67756ac4ea260e90b11ee44432f283919b2d8f7723bba78f69915f0a5c612afb9c8c20fbbde1f4869ab0ac6c7f793b4d1f82244d5a640bf93ddf9493bf7e560b571ab3aa3a8df52d3dcfdf36a54740e1ec66268d59c6647b6fb385afff473a52aa2a3dd28da12c2b1bcaa33e5d09146451490d1baac9f212da59b8d9cef3bccb81c1d5005202164a37a8ac5fbc5adba8c0c3142396cc3551ec088209412f270de0ddca70dfdf25bfaf9ce37dcc9f1b1fdb3b8dc5431b6f2da6731507e1b95a5f9becea7b4eef1741e1a8f960bb2fe29a14ae5bde5fbb81c639b976238a1bd743b62c2dcf8b4329b4a0310197e54bc11193017de487a8e318d8aa40fcad7dfe9db48e51964a5a06299f52d11d60be45ef67f6b5b7b44a3f9ead4b17716e4486cbfb6b3c2415f74b93eb2be2d2165d032166c860265e8eeeec832adc7a1d103c0b2bc2c0df310c9046409a5a9eae69644fed98f40079afc0ab01d7fb9801f808db7051addcc422451ed479ebcb53344cbc5a3b99799529f4a11eef4719179e102c92651da9123eeed36f8c495aac811a3669c07b59e2e55fcc5b2a376628444164932c05ba8fa557a16021c288538fc08698c10421d7e98f0269023db28bd1a45ffec6f553837092dde3495c5bbb7b680a043c7a8855a74b31d1a770eaef1e1f742ce57e7d91445e5ce118f9a2350d524061dea820b328495c13f409c3e866f035dced7077afd66cd3cd5ceb48917c2737dfb23b86c439aab2357aaa7717c1bbeadd164c196cf67fef71975bf441e6862090d2ed77951019fcee2c6b97e3be1d5ec0dcf84209df7d755cd7ecb6b50e3214d542d15094ef102e1957664acf00f1cb9e91469e24067e8a2df09563f7d123d7fece990e3c79ba4357e0597e88ee3bde2001b8342c4d101674c377cf62f04a860d727d690db65cbb9220ddd22caf456a33d124b439702d16ec08651ef3e5d31f96eae57d9a9e5ed0d45d81fc3a339b8e1b0b9f4cacb9582286490576d83f0a147adaddacc2f02020a20b76c6616326e0b8123673c6d4c30f008d27ae1166280597a420a5d28c81b370c6c0b15ba2fe8da6b8264625b3fdc1eab27d07eaeff5f444fec3ad8ad7a40ee30cf17413487283729466a55f561a290f106415fabd0154106e8b3697fb9ac573d46ff1e555c797a07c10a26421111d3c7ac2b0338a8d6affd7210a24b883378f91e74761bf9ffdb53c5119b92609b3a16c2cb2b0dacb8296322226fa1260533f0b33b43d0a727eda5e57a29a14d5931954d9e2e36e3444bfd742ec683b1bdc33109901aedd013f4382c33265d4104f3bf085070eb6190919f6956d6e18f944a6d54eca9dd63c3505f86768d143c2026f1153f75d0de4d556a1b721cc1445bf1656f25fec22483301150f369fcd161509c1bdc4d991ed1492a46f17f8e6da3e9850b585ef8bc829150a382edc09ac6d6b603c390cf9e05ee5e8a68f1fa93d7568384916ca62441da997e22a1d888d9f51b588ed892eb0ff8cc02deb12fde06e7be9a9aca83de45f0d26e7cc0d3037365c1beefa2a01e9d132534bf26a7f8cc85bb26d07b0244736c60e84121c8667f6061d63ea3f0d1b0012ba6dcd40de6aeaf3432e376014e490ca0e995523be917974620bca5182169181d02b21f97d1a611db3a750e13b6fae9407453048cf6b31b6c4603285e84c0c8d763ea8056451075ab3febcf9db9e6c3e4f811cf2acbf0ef682e2b5579b7c2415b7fbe7880ceea5842d2d5355d1239b302f1376db1a1ed6b9978a7b12d2acbea0e76470d218ef99a0db30614c33f461f0483e114a4f203ac69036db05635af48ce048c002e0b16249bb93b5e9615376e073a66a1c72a1165ef177295ac7bcbec62ec9105ebcbbcef8e5ebb6c15a2fe2d36265d341b00fd3df52b5f42911c21bf0cb25f0cc003cb917f448894c05575404e8e95f39c49a404bb9e45a919b935bacef693a3dd598788f635e0ffcdd938633614753751cbedabce03027189e19628197fcdd1e9dc8a439e38f93540c1132655f645d351662dc96f5d450047b7aa03bfa8f2be8e16a67020aa41e45a5991623bed17090c587eed1ef290919cdf689747216ad4889a62e696f760b986e4035a9908e41568eb307078a7a17c18a2d8e6ad9dd9e8cf1144569afeaab38ccbe32b769df6003034d0969fc8492eb3b364ef767c119b5cb4b176125722c1efdf2df700450c29dc7098a13ab09ae5ff7f2534e2a76511812599ff7233d8731d2635cff8f5af0b38e9b92402345620e016db5458f87a7240a18672f23a9b4c533432340da6924d55df45aeda6b1f90810759a7661c1e06c7f38e82feb9f7e0d2cf83223ab7370bc5a05035f1e40fb3dc556107e79403e285f850527bbc807780c6a9b0311cfad9b94963cf5cf5eaeee1f5bfccd0f776891be71f5a0e0c676d1f8d11af37b000bae2ad2a8952bee641973131906ca4ef7e59d2ed71c0b6c5107b8a338724fe820f4e3020f9e8e237889b71e6a79d66de9ebf7f9a360ffb1443ee4be0b5d4a12edbdda0b74766e1fe4d6e47d22c623fe4338dfacb5ba7f0d926ddc9daa5378b5331f6d41ed6546804c9fc14b67eeee0295b8fc41e3409dc94797ac0f071ec3332621565d97bd7cde19ec0f89bd1cb7a6104387770838150659174dc963a5654a6ac02b3433a8cf23360bccd4cd83fdd1e97f869912ea2f20e87ef20ac792de4dccd86b014f1e720cc6e868679342a0f0af778506c8dc3a9cd4f4d3d3303f27ea9873aaae4e778962b855a92921792911f4a6f0b39462e061af6ee17249e5c1767546813c0e7976adc9dc815ca8a2c3eb3e0b38f672923ff55afadeaff43046ba0494a421170f3975d740f4db7c49b922a26440e9a4c7736413400e36f14d85ec097ffaede712301dea0a6b33f73e8c129375d3e3b13b51a9e7d55e0a58f3f6e0c2f53adb7b73f172b19771db130588d1d82bbdabbea5cccec931c075ea75a67c065156c0515b478340ebb22d7ca053fb09c3361247ad432a54fc74d8b42128688d058a70d75d89d7d27b1d3d6604e10278dbde48dd12185a777918e79020cc020d582c119cd5cdc0713f5b3fe6cdc591c576261cfab2902e5e95f6dd5506ead2afad8cccd191e2ec2eb80c724ecdd4e1b78f3b74c06d060d74a1706b9a2a319aabb94f05e441768d95b15a0d159db7ef45cc95f9f2dc19fa78205665287b83232a2a2e70f7edbf2438590543b783243ce7bb0f9d240cbbe667ef3b8a2161a0d446e0cb1a098bbc83440131c1ae193784e74d691c7121419b2ccfab3979e2ae1a8eb457fcccc2e77464d7887cbb1f443f78a11faa14a70f684d4961db4afc6b352aed7e740b326843bf90fde2e816b52be22e156b29b8d88111964e14cbca5da024278870c8946886c3f71c6fd3ac7e04ac0e578591385f4489e19b4b44e6f004b60e5ecc60f09b77de79c2f9995683aa28859729f2804e699e358a8a4d9eb0e7a714e396be65b124c10ef26a2871166180602000c426764ea72a88f87b1b8030db204cc109f560c82a44a34833fd594a19d848fe8e5725cb710942b3cad0262267781e7dfaaea0362e0bffeb0ef0ee3cffe97a5fa294710c94fdfc8f69d915c421929a2fb9908dcca533c57d62d889ac04af760d6736a8f46789b5169d92f346981e73bd444164fc682a63b9aa736b4df7a2ccc482c85958ddbd02e65b7cf8ffa107897a012ff35673818a944b52885c8a3ebc310412bd7c84db2f008f526dfacab0574d898c01acbc4553297b72f1a5d2f2bfcb7209a2c3f030530e56a32adbf1063df3b4bf1b532e4322706c1023d1980dde4dcf339f6721a0f3cbdb5267ac6909ce4d7a9af139bf7ef0d47fe3ceb51ee6497118879592a94c16ef420f52030e4b3e893b25ff2b62272987b0447d01731e055e7b7196219c3e14c4d538391876201b79a78653fb62bf0dd691531013c2680d97aa8b7f72ddfb5c897a3d41e31a5d1dbf716155c230248ca46b40ea00a9556e7d871426f26490c8a90bf36193cef9a68c3847dedca92476f32d51bb8e1296a789cef3f60a7936d875c33a5d06f051529f1429b49cb7db8b51aaec64a759da814e87d5ee54b6a5dd91c9abf6d60737ed4193b32a0c2c3dbf6be67616c7e415ff4d8073431cbd504174cb30c422aa3c9ed718d588237d21d2109e885837468d03d86c733ac9f78d04a0dab4c8a8b52125748eb834fee92ab844e02469874b3a267608562a003e69df026c2899e9aea4dafccd66d851b376796cd1bd893c628987d32dbbc1a9f567644e9f8ef2c78af37ab4a8ba3b0cdcc8de3b16d898779104668ebe3121feab5fb17de60a7f141bf8490ccc6f8fa567c02f7b90fd9112a72d00805acbb3b510be9a0d2bbb6adbd39c51f82bb26062c4d9327dc43be7579cd7855feb17ef244991e77051956c035cea5e1b5b3f1547fa42a4c66c1d37ba607e5635f001497bb981f71118d0b553091141249acfd46b8182f427cb10deaafb46203867c6276f451f8e1670a687809a52498228183a2442af0057e86fc0d940e4608f60623b75c0cfd7e8a5838c6da57ace3bf9dd65f3bf8a50ca1a8dbf32a784fcb9dae4ea790d5f9d1866d1a42d08794c180b78ba8c254c1dcfda85c2a6596452caa46d3ed7aaa3c1838debd5e42b4af3b3de4386c34ac07dfe6ca2b5bca1a89bd3ae5b9ab0bfc3e4f37270cefca38a235d37df50a157081;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6190a26f4663b21b90c026e3fc294bf6b9f0343ffa9c88fc05afeb61a21db8b090263d92dc1bc6b2eb84c2f2c8058cffcbc6cb4df344b8624067df51673ff90d77ec3daa9c872f6cc0d5ba3ff67a8f420382e6cc98640c5c9b7e9fc96b26f984bc132e582c18e2761d44e70af5522bbc07f01a966b7e2603a9165a71c7a883c27cd22bea10657e03850a68d9a8477c79416d41ad7b3480fbd41ad7239bafc00a9c0694e0f5a41c6d1fd2ba3050cbfc45a093895d9be81289c0866503ee885a2d82d9afac9dac5233401fb2fe323e6b349849fb432acb0d1515d0fad685db19d07ebf2940acec115a27e5a692e458a6d2211f8688bd70073c9014a4e6a2aa43d311ebd5ba061653b94d53fab41b5dac1d6fea09472d72fea10f19620a9064613fc4c631098ca0aa8441706ddc9a12d588004ae6a9d711c79d4d73d882d34e97a1ca45ddba919578f66a6b6b01716b9fa9786eece86ca435fcd808928d6dfdeecef33a349bae263c7bc2ed25eff2bd74dc4ade4bcdbc5ac1d942d4233024e0c0f4d201d55930eba08162fc6ce0bbea6bef20bc4b68d229b6b92c76f0157819fb0b1a50bac1b0786f04f523dacea3f7d5fb6001873cf4e4ef9958357fec54486d9b702c76d04ac64ef3ae0036b24cbd8384fc24c3262689e01233e545c04588826de1a501b1e9ca1203d9a6809e7a8bb9e9d90d4023d5576434b50f23e4d09707e2bc1f3fa3758453f23386fc642be6139f4283e0775d447ad140599693c981c6829edb1991880e348b105d3e84950e942a9c7d2c0f81cddf5c19020dbb8b209890f65672fb34e5ceaea3c2d7fb76fded48c0aff0fd48188b324a061a40411c28a4a3970d43e23ae3f0b720b499044d2ede9ef7b53c4476324c7090e7f7c67a393cd18e5d4787601f01f210252847b689744b95becb6cb768a5e410fae9f9f3782d0ce99ca08e32990e6a3d7ae71cfc9403b5384cc09a4fd8bc9e1ada16e155034b4507ea49c0fb6c9ee62fb86e84fd32cfc47f8617978f3402ca61090ffbe3545474dc09341d25cb2758aabcfef5eecedcd956ace28b4ce8af6752557c186990cf47f2375aa9f412dbb8eb5f397d34d51879f0a987410018e7bbf640e0aaec4cebbba622d22bc1d86b2a26659ff87c4d792586c014f14f4de60ad0cc97c6b88ea6bf118f71ec43e592f35583681906c74f02ecda2879adf967c93fa42798871b4ba04c54bd99c79ae9a162d6c81e99a7386a999f96e0943b5fac3d651821476f607b9006922b12e12c09e39cea5708dd5778f1eeb347c7f15cc6552a3f4e168571c34971d83c1ab9ca0b95e8bb5b3bb10ac75d43e23abce4e58d6c33178d92d582ce6afd3fe0278df9bdd57bd7091701016013b85c88603c9f7bfb3510d06e3a032ed849c456d01964897bcb84bb9a4a45108c6013adbf64cacad630aa2cf457f53a2e6d1376d1c34663b21a33c137760c82cba76c6254bec0f2555abe430b3ca415f02752b02f8824f94124c568a85c3f1acde3423a63ecd0e50aa11e942b7db2b208b32ef5f989c0f22bdbc2e4c62ab517044ca3d239887bc2a262fd1a465d3615204b2bda054ef0fdcaa818183641af134eb3ff268653c4c5c91cf866952e1645eb34963b753c3cf992b6437628cf61f31789b52ff89cb69bc30e2c96382fadfc7bcc072e24ff424fc2ff07a6dd530bac8ffdd3773cec8f1841034e5c9b86e169f9552f9be4edfafcdfa17f9314d79d0ee42d0341e5201df9b4785eee689e857519e383f049594a194a209b2ba8237ed4a2cbabaec2875f20b9475abc29af380fdb8556b22184cb0f3abd15457b0e5d6143ac0667e38aac78a9f036c584eac6e5dff2c5fedb36b16d5c88ffae17bd2e67f71a878b42473c841a2d39fa696aa5b83c151994af2dc958064a959cadc62c115af32654c548f270f601f8c951175ae6d77f5776e787584c53ce6f383a4b2141e6cda74a43312651f56403982669bd1d18a5ed0aecd7668002888562af84a5c937460658de2cc8c799b5e670caf497aa83ac189ed7b03615330d1c965ba40045198513b4e43d511eabe14a58d322ddb7a10f88ef0a10e90ecd4a2ea70678b797ff4cc1d1ececc73f8970d2169c7c043e9ff0877c3ae2ec2e496f44fe1d2ad49b95ba5d4c18610db727a4f947af4e2752a0fa8b2259c5d891e8ad5ea32d83ad2374fb5f8dfe763c1604a173299da148338d578f26e318fba9a2dca5ac385d79fcfa32de4d984f1349888b44dfad04add83a82b07c7b59d75ecee4c21c6f433addbfb58d53953d0706d40ba96ad3f30e4d6a9ec4c3e7a666071103ac1a32736ba90de82246fa56ec01f6faa45143c6082bbf7957ed0745ab3b07fbb464a9517f7562c7a53605e708de7be27585289f927aecce4e9832a08cd06d4498ff06d2c21aab02c031a591c2ea9e5c279f9dc3c2cd03ff04cfbad7a1b8fcd99ed5a0f3dce2737cea0426a8b89dc69f37388cfa68b3f29af04b5a9a41eafcf0d268e81d31b262f4689c872cbe1d167d3ddd92f8110fe43efeb2e8529f21ec91a3c86194d16b278970487f414eeadee7dcc8788a43eba8fff123959a895866a3d68af0f24dcdb31f71974e48962dd2537fa02fc78a999a906ac74664ed1e755e8ff60b9afc04d6ad14aa691907ffff3d41ab430360fa9ceacffa079ffe7a0bb04775d79f620b9172bc75880366072004696262c3930475d2bdbb4961f36c2645f162e9574fe1d6fc3fbdd8d102f467b5eb7f009aa8400a899ac7959d371941e10f8ab7f7a36a2e8b86f1ed2afe497d3ce09f92113db6df547e5ea25137a739d21981debf32691e9f070ad33ad5eaafc3071af8f62e15868f96a64032c1ab8f42d66acf07e241cd18e9522c6699829edb4d6a53c41a998fea399b9ffe270d7982153bf2cd9851163f0e16cb14e8a2519c759d080c4b8c397a5f0bd83dad38a424fd242ab9c9167f7a9dc9d6ad0ab7ff54d9fbebc769fe24c1a77acac6151b1bccf61c07b31d943d9b1c7a549fbdf91ce5a287cc0c288159234a82d07f7874259bdf74d7f38dafda215d78a947a4ac43066e61b0d966ea3e824ec6ff2ade6706c7d4658a24c799856bfe7e07c409add95cc464a77393d04eb383219f5dc7ace58ec9355061f7540faacff91d8770eec60f23ae340254eef57c890bebe2873c6b63440cdb98835420d8ed4c8514107a7d4d6449d741153282e82cd7d35bb2f6428c57c3980afbac8b6f4228d3eebbe2e118ff07c8d598ec445e8ef0f7a8294f6342b8eeceaff9242493d33e6b2bab5282a6f3d7ec64278ee933ebb052db20f49e715d3fe17cadf5ecf879c068f225efe3c5dcbf2ffd0cd039f7b76e21d79b73b3e2e7a17f6c153e451bbc2a1648e402e28569b57beb93f39f7e1c926dbd2f96d256e4bad217e4bfd5b86af87d39e3b9b6944e08cf30f027343f0a413ded8ee4da6e25379c364f32387cc5b72973fd295ee0566a803597eb45424bfb3c942318c244cfb807fac4993fc987040edeba0d881724964e5a2ec7cffcf882319e70ff9eb3ca465b3bf82cb8571ea39b30790d0b7d026676ddb1b2aa49bb501b8a26e442b5e627452e76fb0eb8ef3cec42ca07b1092c1c06d02bbb99ef4d26b3293705a6621e0f0e80b8a68a4a4dce2b9a87462817a4274fdabfd13d6e4ea77aef31489e4848935e09123613901fd7b9aa6253706521c7d3ac58578e4d780d7075d3c571f148dc5f3f2465b1795c44309718d5a9bd031f8e7f18f507c52a3c3a389711db2cb2f5d18ff6f698520ba7d372ccb98160eeb682ed0e028d21451414319c1e4286cdc2beac50b2c67fb8b32d70ec9dfcd37516be2eb41bcdd569b2bdccb3d11d1a5a919e4d0d1c2e949246b177293fb8f0c02548a4044bccf7f9109932e48c3f35230efaa8826bb194371e5acd0a974a44e239167b4d7156faeda48df0a33e91b100087df775e31e294500a25813eb187ab26634d26be75e7485d035afe0741c3515505453cd263bb9aeda41e6bfd48488433bd40c7735e92e9842f158ca4169fe47dc14ae07a1bc133093f9d1722e42763fd9df1142359c55bdec957e3343ccacf2be71fe5c6d2c894973e573e73d6ec3118a07ee6ea05ec856748d73f79a677debd11321c3f4243f7672865da7dc24e6b2960fea3b9e0b43e6f04acc71567a06519b2b3509093c6d79faae228914158afe093febb2e7b3f9b2d8a8be3aaa7935f45f66b471ceb11eb9432ebfad196972def28cece4a61a84b7dbafd81f48b94ae2d267156e6e4496f2aaa969b5ee5370f02f4226203fb353d76f3b562b0292a6b6b153493435f41f710ec7f18396dce02ebeb80b9e60c964e1e35d27aa13883b7f71c79f9be87ae636b9df67310fd9690ea94359a93daf21f479b8f1484cca445a56de253e241c82f0949d320ecc80d1becdf296eba3440a74d4f1a4f174ce8ee5ae63c78970f3cee7774e719cfbdfc7cf64b8c0e7f61052d23e058da80bf60cc92036651c8d2aa7681b98cac6990e3e0fce29e4d8a38fd6678e97f0abf1b98424a45e2673c5f69190b9357c5d977357c6b9ec0d322d3dff42d9600cc6472e79b610139dc99cc794b9027f45080a1b06546800b4e6fc3443294c64cd9f3684885c9e85f575447c90a8cd65fb634d946d42296df0aa5ab6a9dd245cb67edc92fe6971a5755b682d1068241f56ccdc548f4714c648336261dd70dfbe13763f1bd645b25fca342109c9d0965063eb3441601ea10f9d1a5a62b6482f9609697dea2ba583c6757b085887ec832f11bc9458d2d773be3903736d5eeb80189b9326e6d8c48d5060f0b4e8d4d70674b3834fe98d1e8bbd7a197ec37b93db2da37cf9cee9fe9856ceef771ae7cb3ca7965b6ebbb4c7fe8bd4865c62753b62250e658629bbecdaadcd7b4627efd6a99e4dd7f19047cd5bdf773d47aa60fa837a76f05a16d6819e37e2fb2f51b2decb2492340bb4368ddac1e4f857e5fb9a8b3ff099cf679dbf1384b30cd6e360316f0df731f2591365ab4c8780046449dc314c0473a3d45320bf54c29629a93ce948308f18879b8c3849207a1b65a080158539369db1ffd0aec86cd0ec93ff29e8cd84a169b3b0d949698c8e070e2e895d5352c5370bde51f5120875c68e2ed7670970c15a0bf1970c9d1b62568ad8bb63892fe9b18a3f878885508734021b05b4b247630dd2ca065c5a0b28a45d8c2a637044738063fde659e72e848c3d7a7b82dadff4c4926583e513113b5e06c6fb913a1250c5f84b35faf067b8c8350413b16d0653bfb39141e455a7af801980aa863d8751fc65dcfaa3dc9c41353c156ecb1aef5c03c6d82ef801b494f5b1713f650e9c1a017fb4ff8f53762297101eed0e4a41dd69242426a766ebc698484334868e7c6d20485fef65379318b104029c311132fd5afae4affa658a18b64dc91afd1c8691eabd3ad1a596c81e00b686f72cfab8daa84f581057fa64bce6a44d9590b5c7cd0b1c79c65c440cb26b838605b363d8d9b07f299171710810019246391e3160c6a22955ecfc9fe71c45cef7af737c01aafa0743136eba6dac41c5a6956b46396ed1264644f511dd78405c7be13de6f61f5b13d373b12296ee709af85a338cbaccd6dee8de66c6087ef63075fb939ded6a7329e90f8f07289e396e2236720956ee80283324ecc15f97209050650dd690ad46c4347bb3d514f6405f67ec52155538f25c647656096d8ab06ace1880f53a3bf323686869118d323164b48ca973cf5d89012716b9a384155ba8a17255df58a2621c7af1dbcb20bcfa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h266f445adf7848f17aa25c5b40b190fb8db051465e61de82f9f27584be5f37f1270c9a969b6eb791973538fcf086ddd2462dd44d9de52294888f88f63a0af291795476f71de4b1981480fae60e14318daccf2bbe5e45232aa54088337bba88dcba1d00f993f17628868af82ff8110f9ee4c7909e203b07eee694ae9a1dd557c6069227ff25b166f14eec51f9199548cd4d9fe92b33063e61936a32a35dcf9307c77505dfc3e72b5102ccc6deb4751cc56edfd9a7e1fe4ac5163f3a5e970927d68ea354219a177879f663f2f126833e335dc422eea2168023e97bd779d0c8b7f905119a1f9dfd99ed8df10f1fa18307b136cbfe60a8944a11449199785639c07108a6437c56014b15a8c7a028bfb2215b0f889294d07e5f4c2d5c0a5434ae420d56ddb5cab68a860b0cd00f5b12f70c6c615b57a32edce6c459222602e939cd27a91736ec9515d462bde0eed1704b89107959d7242798bc23766799eaf0b52f7e07f9449e2c57bb925b1a19d958a7b110c7fa21b149c88df782170aaafacbe2f4ff5593fccc32bd012a1f5113ccb4f27008b9f9352afad9175054850e719926e620f20bc06220462b7aa305ec4bfbaf60a49ece0a6bddceaec0420c6c79b7c23084127daf89c49fa76f539976d3ac2692a73f0fe3c16c1b29f3bcfcea2326cc58a3bd1b8869977d64b8f68083123a7ca89a3c72c7999d1373fbc998bbe02dc1e31c24acfc964b22b3fedd814fde6ef4f0df2d2d297050e900ec634e2cd0c21645d710650bd92a97bbb99c21077a0cf32f7ca8cc92fe8c27c7c7c11343732f31aec58f74a45dea719df20d97e8075edd5137a35599b6cb5bd07e87461d15460c88b36d82c2ece4aaac4312eb73ae43375c0c144d8fd07ab7af0541fda000862a3928f117e7c9929f8492c6bd01a03f7b703d47154fe50d3cf3410a13eb2cdbdb4ba44f52d819a7fa8bf4417dedac4bbb661b4bc8271a08226a89c37433a83911123595d21a632d5a5a9084e3a00bc952296ba2ac6a305418aee95b7f253a2f259c702718c5bc3524a7942d6d6e81a19229cdb8ddba8d9a04068283eb4422ed79a05878d5afc0ff302eacc37d317ae52f516a0fbaf0482bf4c44313f92b01c8ce0f81fb0fd39d33d3ce3d96909d688352426d54131393b9edd11a592f721e7321d763124d7fa0b4beabd231f04f8b81d7583de124fa86de93ac873d27090a34b345d5b8c6274674189675136679e2d9b3c317bc76a609114993834df88bb2dbd6c2de7de48242e7785ef776de19c2f548ea27ecf8f9388b29abb0be6139cecb8d2bc341680d9b338b32a2641f684b13ed5d90af6459f55414df33892848093f55ccbfab740b4a28eb410848334352a2d7cf2a5c61cadff078435ec56a449f908c46b04ccaf8e40896e9f13d12d214cd2d11b72742df9dbccd261917fdb6e67806342abf867f7ac72811e851b910d793f8529857da15e6e2125a2881aceae9cb7d31d5e6a38d0e70a40dc5a059cbc64deb360f5f0e1f8d1b5d2c68f480c867e3c6e5f0f621060db92933a1fdcb6818de710b0322367d07e430e9e29af8c899cf096211c569bbde9a0ff4ed7b7050f5ddb47f8ef1e9445c1a236f226eaa6055a2f76666b02a32257f1db928c4f68c31baa5358a58efcd70fbeb15a86f999b31adca68cf7d85a37179eb63e053cfead062f8acbd056a1da9b3ec5ca6d71e8078ef57e1b74c4434c82a05513fb5bb33463ffbe759452147c92737f03266951176f7ded1b813975b9b662ac03347efa450a2c48120b2abbf1399bc5e0987502c972dccc3cbcb57992b8f43501573593aaa36434fd121418cce4c67fbcbf1521a0bcc2dc657c183f4c7d74dad03257702a829d09bd4d5cc4f30ba42adc37110c05eb26b159625f1257e4a3325a90d5798204484286f85d3a900e0af65e77b2aebb258bd6077ea974a0677e08b66042a8ccdb501f09e0ef7ec3a68671d6ce89bca168b8b7e7f5317fd7a6d66cd4a4f10eb3cffeaec1f8a30475cd27911c30c02a87fa8edb519645916baac9235946eb05f4c9d10d1511f1020a11ed4a295c41b4bfc338c97eaa7cc596aa345a59e0b9c1b016bba50a5f854d8360a71b0e479dd7ee2ea1e4b94c6dbee07fa253fc9bc1221c9343c8a34154b6a600d5c2eab8a366ad4fd32b1d00fdb6fca6e9a5632bed81355ade7d6a733f1aa90d94703ea5b04e47f60943255ec7adc58c809db930df4c57915706da36f44669f2e47ad9ba7ed04d4baf8d27a5ea126a3c8187360c639cc828ce9b3f128b968bcda9648b4d7a7d869389db4223ec1d2420cdb083c184927297fa432f8ebd80ad61cbb9db02e3e775ad65414b1804709a5167c06fcebc491ca0ea509acd82180d844d58d9ea2324f55daedf596c003ae089ae2e7d60a97a5bcf9bb87df2fb3a1b885cd74441ae48b645467afb39a80ed59e8a9641de71956949cfa79e993dbbb0c09fe3c328f4f740cd1d4e0a52313e044c8ffec1e465c1ffd39c57271189848eab07d2b66fa6c4ac436dc67e056cd51897771e08ea87ca83a23d8a2642bb91c910c21317779e0b47ebfe08b360d6df45f14bb132fab482acf6a6c25ad3c2a0361279ee7efac77fa3ab8bb8f8d24d5076a308351cf75cef203ea093d16da4ef21fad9f21483b071058f74e9a717df7a5b335b4008c31e22df634680ad77f89324f1100fb6277ac2434d5d4ca3666f2b8a18ec67d24e8dae684331565a2f40f2b869d016847c22d94b32306041867b966e7ad5475df5c8486c179257233bd7dff13aee12e611a0a81eeef16392838b79acd73473f543475f63a010b571193298c92c3befa5a6b3a8a8442592f0bf55b27b71dc5aa5736a2d6937f37b2114e4c437c7802fcdfffd11ee3848d2e00f693a02818a946c20c742424f702ea27bc83839c5a2f70870fc290cc60437b2d9c95b0b438f21ce550696b09f933ec218ef4a73cd0c37278ee1afcb903faf4ae40eecca5d445d4e3321098942df227d0ed044137b4c12e586964ca2fa1b6903e4249dc3fd905a6ddbfd00c356ffc4446a1eb73c8d0f1863d25f8be05f81b8807b0d4e8f4f490c173fa651146980d7129438033638b3c460455096bacd826102165746757d6981566ea39ba67662dc66f24664063b8ae8148b00d6f4b6d3d60d382d47f465347f892d2efdbbfbe5ae2d8e6071fdb169dbb8e07d72e89d90c52c330f8ce58465eb2ee2bec882eccb0021134c686d838dea6ceaaf1a2780c6abedd2f34018923fb40212b288d8e7742bf6c0a3c84d5b86eb3f05351cce55124c090bae484433bcd8b0a77ea4b82da344809313bb1ae039d9c86db1162b0c10c07a097cbbdb59102c68ed111fa1250b2ff68169bfcb6a5dd85d90f5b563b0386481f24dae2165f726612e51df3e47ee4d90a681cfd70810ac068a740d23e614acf64dfaa90eb311d2d7be7ed91f263c74b66af37bb00bc3b7272c71340ae579e800429a131c30c24473cd35938a987813c0a44ebe3c51aa7a9091b48ee1af59c821116d28d0ecfd054613ca1de02d6c941ab7429c14542bc4fb4d0611a9bf154772ecf91c3569f2443e1c76bc3cef5d6b6fe33e8069bf7f9536934a1da774d0bd8113907b7461d88f4acddae5f2cf69570c7e4a6cb6e888e33a5e173a7f54f0af8b02df69ce25c9f1fa091557758fbbbb593ae719890497cad5c9b83c98f08fe0b45f64c543a3c7dcf41fcc1299b13d75befb52345cabeda6c38398421af70b60009344e8d45aa81f676efe2e1c0a08332a6f4f7bfc9a3f2e2a01b6981018d539bd9314ccdb2504a7533db9a8dfeefe3b4ec48ba58beb01755dee7e7333c4af83511d5e5339dd81d62ad36788bb739b5e4694617059087a755df7f44c97157c649e2bdd5330bf9a908ffea9587a12914b3629d09f98486944e7087b5100461f299bc0ce0fa06094e3cbc83d37a7e05dbccdbc2cccbc873ce2d802df7f7cc02fc10d07509fe46cb8992c6b7c1aa3e4201acd11cb7f274aa046c3687cfed97d82477ac2d7eb1a1e164b7382594607bea4c67528e68edb14c73ea7f213f0982eaa37f058bbff08f49a7b8a275506a9a16c7ca7baebcb169a1036fa4f2782b441b0a5dcaf4479d06a4e9276643a0942caecf1073c70f894f291ace4aa0b0b79faf14cfbc0f3d2cf3dc1c884e053a8b7ce5aa8d0a6f839ea134f9eada2d41329d1edeb3fffe583049024621a8c7099de2987e1c1f83a708f893199b000204b26df0a530c0b2d1a5d193ccde88b5c02d40409b7913978bd2efc102257f4aa3226ad60546fcea8584ab02af580c93360869331a19ed6376700fbe4212a441fce811c6d1f824539d04ffc7484394cbd5eddfe64a784fc73b0a83e540913ea12c14168d9e1f635e2eb11415e0b0aa750906b435dc168352a06ee1314aa4325551dd5b28c915076468d5158ff1e8dc9707ad7be8ae01af206c67859059653a8596440b9529b1ae0fd03d52c72d94ff549166567e9a0c9221cb3a9c874b378a6e76d83e5fabdb8a7afdeb63f1fd904598f4981dbf7e0d798347ac9740a3b2a6ffa241960151c26820382f444e057f26f3f0c66629b0e13c1b7d0755fd0bb0d4baf3dc5b26053e708c2aecd61024ad0434c2920efa425efc600d2a93eb7f348a59c3b0c63557a5d0143d541d29b482c7c9212c4acf645863c5810bf5de89909548359ac57a2687e5e60e4a029c0a5d8d40c71c7d17b568ef29192d2c60a0ba2f60fe4796c2c6db244d9298493cd13bb7e3d17bd8c3a97662ce1507924231c85a264d76afddf18ac549d13187643da60726d1213c4752cf72f10a5337c26de23e792cad30f7436aae79c0fa7c9ec58ab653c205002e5a3faea554216722f3b4c8e9cf624a80946da2ec25b6af7563ebccfb66cc358ff3053008e69b7b89ec920917b7503e9d017f580b519c07c9bb24d81877a23d5d0b04675b3815c84d13da2a17a069e7521234082412e4da9059a070c12d948a46249b60344b243459cbbe7b49e4f6ec84878244f8de2f0fac18b5c4edc37e620e121782195d7aa36967779d3ed99064a2c071926779e014374da494c1d8fa692d6ecdd6bb4da86b0baa56a1fd126bb0d2f2fba2ca8ab7db5e730fd2fc826d885c6f797fbda08631c5571421b56cbef732845e792acaccd6c78786eec1c432101946f7dba21d10dad87d1316b3115540e49677a89527c4e66af6ea327c0c6a54b6bdee0c1d0ecc51a1505351d45de870de493354fdd96e6ffe72444446fb72e687477d43fd85066423e639179da56b3af8de3ee70e75d5716b7dc75dd360db34c2fd686f3a7837cff49e0d7d6d5d956d7d33b56b7e2e6c18c235351dea7c0287c032b5f0703e319869fe9712d8ab5d0556bdf158c12700862b02c289153b608d02ac50400954bb10209869c900ec7e72201dd9776b54ebd5f3b93620b46b016076df57445a04a8868f671d79a2638044bcf22da58d544bec1ece5e1b8ff6482f33906867328556b49a665782abe79c23e651eff53d31fca499d87fd260cc1cb216c9669d9c12eba2b2bfe37862228bb5bc8b0d210a829751a60ad921092f15c72f4af9d4caf2493741d5f3ed45697a7dc7e6d554983bdd5b2bd3b3c5a467c5858de13fbcf1f48f583a43bed2a470df036bbc7a4616c6488ea787e67099efcc324351f3f28f59b75c2deb4b0f13088979b56f817a5b4a2cc2b18e6e505ac59df99974932848e59c387bca60d3216d04387a1e78b214b921a951ad142ccfa12080434f95e5ac9d2497de1fe3bfe42e23abb407e6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hed2bde8da1b2ca67a0f86ab3d792fc8696846bc38a87f4f26f5a6e69cd7de4752fbd95558cbc6828da2f97817cf6e1f0beaf8ccdcb772755009d8fb68cba893da039cce4847d7127fa896c236a608e4ad2799a573c08ef7d8090a2d387398f2bc0f6fe3b7e49b02f7a69c7c83ff256c9645f0001ffac4dc0944cbdc429b4338c859e26d12a24eb1fca314314e516c25cc32a2a96ee1161567033cc81ab79aff84325f13d0fd56726c97a71c1060b44e812c4f8e55370bf02f61a19ad6e01624aa93e2156f335b3585572cb28558447d0af8e817380a0d503e4c2fce06d6b58593a2878779fe2152bfd4a1e2f26490c9a3d74e60ebe3bad64ab6828d3e7d04b71cafea307816b5bc5e68b5ab29f9d32ef8376ff1c7627d13d279ac8eb3a9980a9559f705eb27d20a704ce9637032dcb355c85cdd439ff450001ca65dd8f2b319f252a49d73b2a662eee6cfe530c9130ba2842b5fc9ef3fd5e0e0dfa8946c6514404273ade29119d49f96460619b5b784ba8988739f7d296cfd5f21189bb104f7414bf02807b30f4e4006c410b67fc603137b4d7d4d82e41f5a07967fb307ae302cfe8fff44fcbe54d170ef1d531c491eaf4166fa5ed28c8644190c59261bf872b093859c76c4cc0a185d7c29b5a90eb8f570cb526d64ec30f4cc29711ecc8f9bb74f39b7562fd1594f8ff47f0f0f44df4a1f6224d594ce851502e6879743f5a332aa475a7506a31dacdc4ad573901d309e856070302fbb662228cd444d3b3eef4fbc8e6cdb5e1fcefdc9735178581e54c0da1aae9163758d5563c5585816d0485aa646e866bc12bb9b56d406a5d9b87ac54d90bec6e090a8fa9ac882b5e90421569818017e3c0dedae58fad46960e0a5fb659336dcd5bd4e21fb891c476b7f368fa06bb742f5b877da64fbe8f360063848c5db3eabf6a4613a93beca91b714f01595d49b10ec3b573fa96a6e6cc301f9067b8b3a47cc4485389094265fc6d24a97d28e611fc62aec3975f357cadeb4406577c489c91184e71aca5a73a3a601c0dcfc9de73d9a30f2eedcd0b414dc31f52b70f2b508119c6b9e724f232ce01c9fb072fc34c863f5fce74148486d14aea635d733a5eac8b40422be2f388d76471fdc3d45d243cacd1b409470f6b3fccf058f68bc6fdf3d1db8b2e8c93a2c4525278530f5cc47708bec0f79a81ca6e8a6526191116606a9581c3f8fa8133482e5b300490333e72582927180d25ddd64f5818ac5286b16a8adac35fecb294206917cb48f139a6d8780aab7fcc5fd57a17dc803da7fdc562cea19db289b788d0d0f3271e3ec4f11d0a71cec8feb07d13744a5c390d8f83c65be720976038ab6b10d02d7c118ff10fc08f629435355c0c8f0aaec9ad8e471f9c84687ce07eddbb6eda0bafa0bf45c2daf4a5747e36c841cc171a90ecf41cb695a97f784126a70cdd9759016a390390aa7fc2dc2427de89235630891e4c283af4e22589514687775f2e3fa78d8ccd44f208c317908badaf5d55c35979563e73f8c9fb331d5a55dcf69a5901993443f2002279c60881fdb63256c36f151928362f0aaf959c57496c7ccebc113e5ecbe5926d391c75e25e997e1146c52017d7cc6fa31326f687ff8908be39b7904a3a931f5a68e3e7380909307756c71c1acb9bdb3967100a22d48ecbf50f9d9a8604524bf36f0507d93e3d2c068430379c7fb12524420213a0d831755fccf8b4136cd49483cae4eb0d84da5e18c46875ccdfd6e69e88480b2374f85fecfd9995b851eb65a3a9592f3fba721d6ab5df9a5d8270fb17bc2b05a9be68362cc8579049346df70d63f27f33382c3e04b77e86ebf49cf9cc4433dca21efc26b1c1fb8415080ab9b3768544b5f7d3c6edcb07955b67d257d65f1224b95c5a1e13f3bde9d829922de57c5a02fd62762029a4d3670b66d809e6c4ebfb2faa31a4de093ced4adf0495befb1a64e61c23493b1f4a53e12e3c616bc2e927858a15ff4c03a9fb5d59dc1083ba15051a49865fab82f763511fbfc30709e4200f687ddf9e170e7b4e5ea7364b7a316b2d6a814ac5cdb4c45739f9d8273476ce4ffa6c8764a4d5275d6bf35874f9daf9e36467a8a0ba8d0242c1be521723db7db589c9cad2caf23aa822e99ac87457408f36e923841ead8ea2d2adae4496481e9a759d55511a359203153ba4a92424a4a81ae4dc6028642a67961406126a573eda8d821e14a4681e76b7a841427a112ea3bde62ad1e649b786dca46cab445a052819890aaf090ea1bcaa6814bc4de61019d065893b3e925f61caf9435e6635106b28f9aa8089f7bf0ad607b167a57ebb10992a0a9279dba88eef004ae4034ab5fc9b8e0c178063ad203b90dd455a3e78c85c95a48bf522b87f13868d3e018d4e279edc62565a9d2a0ed84948d2bd8e3a22155f7888cb34eabb7afb1e71b0616fbfcdadcd4285668d6acee4ef2c001974778f5564cfc13e0434282316fdf7cd4bde9b48234af21a15a3997a9450a1b123c4a543fae19b043de95488f0cfb25bbfc48fcbd57d979f64745ec7b9a2a9389cdf38a01ad56acdf01a096269a70b8b4c586c465653c1fdfed4260bc83c774c9992140bf1391785695234c7d4953209421428625798338c692e96f34582420d685d0af337fc7d42fd6c45c36e9d9d50a4b40cf5cfbf85b80f3c0b56a7580e8da628164732ffc77f66e27a93ab891c14fe5bf60caf31cb07b2b2567c0e7101f400d4281361f1d917c702670e0a2c0b1eeeaef6984e34f45a6b66455a59d9f2b3706e617fa23f1f5ec2f6504994bd0a459675c496302640c5df365188fb95a0338101949fe80cc873f0ce5ebaed0fe7ad7f2438b0c4d27070e52c4ec3bc7cd48595970b6d06c1c65226803b04bd4da15716f798bf5cb956cd06d4758347e54f3c74f0be3fe1ded1e8975b6e3ca403bf60414a3fc355ef79b36e764876b0c8eed68e3a12e757dc27e68984902cd9fae2e9f336e6183ca6d753f9fdf750617ed4f18bcd31e2700d1c6520972e8f3a7685cc22c0195991316df062b242efae07656a46f16f7b00f0f14c8fcb57ec302ed88bb7db749e0258421fbdb2e80840a4b3f8f75ca9f603ec46f79c795132dd528aa5709694928ed495e0c49887fdc19ec4eb727f04a9c09fde3089d9b7a31c1507eb8ead5a11debfb85d73f04373222b7fba03a036ebe9004f9748564471972b36843be6aae80f251b6842ff14b89c288a8983cb886476293358bc28c4d2621fe796594485beb2b123731383765727cb01d4154add0b5a3e9a58bea5daa2da8055d04f915cca44356dfb4f150b0dd487f25fa4b6eadc6298be1b06bb96bc6df8caa983a65ba4482fdb23532fb59addee8cf445adfe60726fb85537d8176c7071568342547bd336490adf2b20744ba3a77ad46ca86b1b2bf5ac111c098594743521a4afb4b4e1133d92b7153dd12c34cd0f00140d0a6dfd35d8624b97cd622d695843059ffbfd6f35d24b3a907819f55d0f6e5ee079d9b1b36e4b38feef417ff57fccbc636d61a9f67ca41f485abd38981b513af8decc69d079f00ddc4a0f95d5111ae9a7f8a3fa501a4756a4486e904c5d30e412d7897799d18255d36ff89fd8b3a1ca7de5b22c76569dd5ef5d7c75b70154402fec89f20fcf56362e29e62737d3e0c900d74fbb6a300f8705476317484747b3337afdfa3e9df479ba68eee465d44ea510d66da355e740fd764c78cf24b28062b61e092d823043e6741267769aab971cd8982cb5d46ca8fe505904a8d58cb68791428e34b1ed314948257746baf4fd24feb1897a9073b6fe2cddd7fbd7df23ce524cd8427b7688303541907d0e84e6be56bda2fc4b778dcc43eb375cfd2e89861de6de3796ceb273d675226f30c475ce0818ea5c32411a2cb4ad64e38229eb00877c9a912f4f350c04ef8821fcfbe39f87143fb7471233cf7e673f0dbaddc3a9263cddf1453502bcf652b4fdcb3ede6a114c9dc2306d947e18c1dfec9388c338dd1ea8eb9125412d28f44bbea89a1a15b79ec0b0ca67b8585ed74d3402393b8b17a7f8a4b00ff1c8db36660374c4d8df1a0a1790864bf3e4f903bbb273aad3d739bb0f07b830b8656624a98e0c0a3942432484583b7ed805d7fad34da2f96cbe11b32cb31716e24ac9e9f859f486a3fb00a17a6383c1b5080fca07672c1b849e69ca7fa0fbe2663b077e80102c7be1c3177bdde6bfe363f9f45d7b5fd6ee95adb3fe630ed65ba0bf9b655a962c2e5483f65b89ba30ca0080112ef8f508837fff60ad3d250524077defe7b50101e059cdc823a1c7902288e56e0779ce5893b31be10cd659991f975a35220abfd0f6a119cacf42d442383c3d050d6a78339251d0abcd0ea6fe7e11444d0035c99cc5f69013986be0f33b9f26e37ee52f16fbf5acbba53c286e625cc4e629556d7686c0205d65404820d5441146eb2ce69b4565f87a60764aedbc4270e36e061d551cfcb22b690222868fa3da1e938b5f6dfc932a0043bd6783c9e75cea042e560f586c6fedc4453647d1227d2393c063ab311c1166b6393a0a1d57a3c6e7f5b0d0cbfff0a6b8f1ecac0ec6d5f0b285d92ab1aa9dfe8fa126dde8bc145bc90191c748f50a7fb1c91b12630012ebfc8e50edc5c2057df88d9198f721e71c0f50fa7c009591f68845de576db132a6f20f2e4ed0ca7d58f6a2e64779bfff155a383a4de8e5e5c5973449332c817059980a468aad9ea8ab23659d31c8f6dd5850d2615f8a9469b437470b6c3cb6761fdb8a188db4a4fc5e7b694aff4e1468a3c58f35048ef146085f0b363e32f1b3b4ff89fdee9034c9c6462e8f92d265e24e17582976547be150283a3fee24d037be5b1ef04bb684178a651541068f837bac2b0d7ba49ef4392dfd4adc73bc8f17ab947241f5be5f6bec0b27feae4b5d125459deb82dabf22be85524065e4d8b08e1a22a7fa7ddd43426cc92d2c1a8d78d5830355a913cc12bebd52b5fcae6bcc0edcc95760160745f16fc543f070c9b1ebe5a09a36606fdfe0c543d703e7c69781273918d273cc2a157d1d77979141a8d016453e1de61599f46c6e2749532467b52a9afaec9be23b2c83d488b437a7e32a22ad2f4d9165a89fbaa31a38f6eca10bbc8bd8a566aa695c3ac61700173b9baf8168e990f0d0c237faba215366b2ba3b63310271d573956f1bef340160257cbfe641fb2135603d7baed3a79742c740ae39c704264c76c2ac0a08a68e9ce4a2cb11dcaa53708cc68d78d855851d4f3d444e7fef5eec59dafdf6efc80f424a0e2896face5abda11b50556303d0e16c784b3e9b16d9602d48f01f478669755666965110375b0f7d8164f264dc678cfcfca3ea2724a25a6864a526113318c19b18110eb57f2d2c786a9a70b7f0fe04d9c7f4517c964618657f1e8e9ef9c53ef922b1d336be80f2d8ace94a5c1a02a365dccf1a2eeefb3d99f5b484775227f871817cc92b11272b60b62fd496b5c3b43fb938d8ef1a4320f113e7b72a4d1214d0a2effc917592f527157b28f033b1e0be4619f9d7bf27939abfd4d5838e0634eef2fff1bec5b3d590644a257864187dd243556cd2ca987e8beb25ce491ac9ce9ebe0e5be6e755d791458d2509a5bf889291bf12dbad0a2876e5ffb61ad9932f9adad9f6a5d98baee4974214c9a582302a99e66556590b54217a40bfad3bdcf21a869dfdb6e10f7e507e2b7f9fe5bcf29d30b94f57ef43d6e9ed0496cc56e48f020e17a0306d31955d4fe8037a13d49aaa4de89b2c84706aee44363cd4339a512a0228f1fc5a76bf33b29f5eefba304b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h52077a454bf317570955335746179dd29d21c17e9488c2c23ad7df75d23de27f9a9b884931b14c85c52d4619ff60a69d5b83336e519de0cce9e974439671220dbc2d63bbc46271e7d57c4b07d62e0c8449791e8e4191fe7db14d67289f6ea9961c68ebe503f5894e003cd55ee49a88231303aef907a63d0e095193be51066eca59ef84961869373397d257da3952a2e7a35c552286cebef955faa8a48e4575c7bd3782e84a243c9ed646ac724af94c4af8b06179360fd24166f06aac02db473ec6dfe7619197aa35d20627f9ea779e4642f4cc947f81a60f452d632dc99dcd89dbded0a14171eb6e18920065b5a824fb7f206a51b690608216f5030712621a947a30b5bb5901af0092143e6a29bc3697f670d39ab339b401b281727fdfde740619ace1bf59593766dc69672cc391191884f51957ce6b647330887c454d6fcdefd853987e46b7c61c958e0b87fad414f17b20b7dd5b1645f0ec547f0fd62984bcc90fd7c7de3c6919046993471cd4bae4ffdabe2b729846f20da31feead1c9ec246f8b1fb49402a84d6b8efb9aa4d8bd09df4f66d90ab9d01b373f8f062e43fd89ab0de62b7a53579d563c3e5f76cef06d5963ec1af1d27f33154859e7e15ec17f990c121edf37aa85bda7667efc05df486ed856dc52223ce610d3e4de9acbc2be3c8ac85f99501860a057abd2b760a682cbfbcb1eac80d2e12faf0c99293fac8a425416bd74199ccc77054a6a5741d74ea28d7267be4d654bc0947aaeb660743eec20e7dab4c8f5550e2ab7980a239d7b06f0abee1688a43e33b9c80aed3fd1a4caa2f266b0c9ed7fc54045d1ad3b19095141d09536144b7712ddb0b7244a15e04b2f72c82960c41cc6d58faaba1207536afba86ca147ef0da4ec43e1456c4c44745c76f8863e709335d637e9b77b368b049e174b6ac004f9edac1c119c516de49022b05767e3b014935b6f724a98331a761e73a5ed77ff8cd13873ad02202a472e68b339798d4e871e372be6d9bf252df24d4d452f5b561ca4d45d05f3e5694786ad2c81f12618364f90906ee65a8828eb2e3defd9efb87ae0f764384ece4ca1e2189f669a22af7c4e3be6b212f17c722ea420e2a604b2d69d8e42c42060f56dfd3e32109ef719927f277b048018c4db413f42276b716837a99fc855236be1be43b682a2d6d32420ad4b30c5ce1b93801e8e441ea3aafd3ba5d72eec27824bafed631e18ec1c20a969ab6e0c92403e35989cf190ef0e9e98e1f0910261536b1099bfd65cfb36ff457d5cf490e86ed9d5f9c96777a0984764d6629f20db75cf19ad37e9ddda0fc9c0f5e789d1db170fa6287465b36269f7e08644a1252b501ce40051524f01f5d0554a80282c91afb351591e9943af2cdc82b391bd386435bcf1091d7a0c7c44e2b400b852b5158f99bd639af52606a08979730e343c07fb3444c4b032f11c5c45e4263a160715825954f183a77074d85e03307f7badd9516a4cf2c453d6d9a7f60327e7401a19b44f46ffcebd59dfa35362485e95b57467db4564e7f0ccc576000d9d0383992259d4faeda003ee4c67152e3c3f1a433fdc8ca268822bac4592f5ca0def91b623ce53402ca937ba95778587ba2e65658bcff2978a56c4cc25704a41962aeabd8c1901e6e1d2d7e26bef7af22def57b232e92501279a4547e1567903a218dbcaf63411dfef0c50ce4e829bfde09768df3566d2b8c6b9d59d834038c2cd91ca8d3c3633538e088eec26354366f860bf071bf614353673f1792fc0f25606e30c45a30f51668c4fe75b5985c5669a4d3db56078c7f3f02b259da6c88eb9b6fe17f09203661025b53f31c52cb1779b16216202cbc4a1205cbbdb8f72dbb98242d1352be7966f157afa149b602c8219901cc622d9b0b0510fcf5dadd62721111f8a76d08f26cb386a4a4f58885b03f27be5337ca86a6de2dd40dff999746a0731ab62a3e162d14d58194fe8084e44c2cb471ed73696fc2c4eafe3ccf7682976b1281bae5e76044d3f33c49a94d396ed8e52632f70d8774a4fbd07466331a1a57f939d04b5c5a4fc4bbfc164d9e9e532834512f8f6f7409e4c298de6e4a109e0f3781991a43e35fc0956594c9c418720e08f9a65b500f9adb31b22882b723b8422c764a25fce0c83a9d24aa19661ccb27d2f4702806598e34ca066a6123b8a16381bbfccab9e91279cb8d36579763c11432d1873576afc14670b84137e7fc3cbaa3e80896c2a53e37d9c277c9f5a50e85aa7eeb18655bb23950257e6e779927eaae30ef035e38efe4e65799e903b68ec340119598a4495cf8dea1a20e3742583973b60073dd2d69f1a1ec205ad63d1183de0b9f178f256feec83797133637fd820b0c5bc852fd40f9eac8857a92698fc3b76c8177be6ddbc75a0f73f88431c1dfd7ec7dd5839fc713f5b1f517006756d8ca9432e3afb40eafd2684339895ca7979a5c738e4971668f42dad0a34b8d2b72fbed11ed6a8e3e48b8f46039f56f0eae9a12df78f526680765e6292e634ffba41b67c1fa1546f3a398ded1a3aee35b26e44e0db2cb2bc0a17fdb26d9e5ca37939cb5a0ebc5ea545621c3125e1bc22864212276d6b0b8cd0add8eb0021dbfa4133de9ec70c6db34a8dcd5c1d14fa7f5b99ea716925e320b2d1f7251c5e9742416e75123e102d634cd9a1576508286b0e24e614253225dc18637f4a80290a2dbe1ae8d995ced590524be6579349e0ae8f323218d8a1750cf12379d797190fec08d8f55f9955608a57cb0c7fb9c508fcf8699ee7897477a92554751ce8c7f4e11f30b1baea1c44f63d7d9a597d9d34934adc268cff85bc7b8d955eaff40b2a43ad8f8480914d41ce1879509b99e9d718c9ef43d5a23dabc2090b0f84638fab2e6539e0b56df730ebecd5317816bea23cab55eae9f8d13b56f4fd38fd46674db502fc0da3afd546f3b4fe54bee44077a9de40d10fab0645f1df392ac791a4c90c69486fc75a6ad089f8f9bbe569994020a820fb8e4138e9b7847e2886c97f6c42a2d328ab59cd1c195b752e042dc3183a0d02dbab39371fe54630252ba0aaa04c034a781593846855210e62a1835c4b5d69b056ea6f2f4198c9df5647785fd501d78bf1f47a758261c3405c2c0b0845b5ccb1a41c0b01f8707801522c7312635820ae192bdc45d7b56b201a3e0d43bd6894edc65008f3c77a2d4c1791b5036af216b9be4bb7fcdf3fe791c525dba4e9eb5a1eeaae14205671840ec15acebe1b5f6c4525a298ca83158ffcfd2ba886a27364656f8637d98eff18f4a6a67d478771415e21840b88906b71c8cabbb95926c271090a3355b8c9419c941d28c18d0c414c2f9e37248f48cb03ce9f2108a544952ba2886eb0a0d3af9aaafce9f64aef558ff2c63ca74633bce89cdcfb0810ea15c74b3d7924202891c0176f073e7ec3f36aa62eee07fb9837fc6cf3eb2ca0da9d116a8a58a7e52b72e5bdb03e3abc39364754d9856553f357aefada1c556655ca6594c2351d95c53737d6062b7c0f4b1e79e8bf5faa8a449ee1588f30f6cc5a5c5dba48e7243c5c401f855fff7ae3902dcadd65fd23e1c6e774dd16765449008f3a0b767ac3740c4d85f5f8a5ab190c9f46ea4696e0e3016cdba8363ef356995581c542325398c431cb86514d6411e40a77d1c85b9857d97fc16f2dba4f57a85b6892b2407ca31b75ff09448255f884fecfe3d4b51516808f3fe954e563003a569e27de8cac6bad9dd5e3f3cac3a23a5b74eb843542c47f71f8e618a3ef733ebaf83dcfc41c84e123b7bbde5b0aeed213171bd4487d0ef5593f3b7cd32f9421a3082dc3effe9745000c156deaa27b9c23cb090a865af24a20b2fcbaf7cc2ff29e74c131f5cb33512c62bef9eb04d2116875c543a803aa33c6eb13dde6258d95b1422d473b604dd3a1697973df452ba016cd8b8af04fce90e3a033901db37e7391c75c6692a364924e96f438e1e3e6e434863aacd88dffa6982db026b85239c4e54f3d30442a701db0eabeacebbd312e755b42c2d8224363438d3a9908aa86e6311b16cb9a19fd8b3bbdda8ec43eda796b5b10bbc2df94ba69196c2862dc037585721163b331417e6d8ea4914ca1337d092cde4d7676cd3c60342158ab6249a2b7f795ab1c88061fa491c93df6919aadb9e8cc84170eadb6dbf9cced6a3675b5fdf3261620adfbc21a388a9705484c1ef6772f99a1b6d46f0c54466c66ea0864b4f5f17490f96822d71af94cdbe2df686440370ef147f7de889c7cd4a42e9aefb9572eabc59d95ddb9a1349be1e14a1d3ea96efda4ac6a8bbce3d408aa2c14bbab3743e15b435f87a85243c3863cc89eba7a10cb0bfecb528effb546e4179c61b55226a66eb5ee8fc58fe736841ec277c24023c41c6b2e87e7a07d39c03f5d618ab2d5f8b0fc2401fc9cce09ce374c55540bf9158086920c3b9815b77d14866ff65e4f5a95e0e4019218b38eac9c8d3fe93e0d63939c9bc7923d4dbc555d786bc9278a316623dc1f02e3da3d15df3d784de7414422ff99d1a90ccddf2fdedc07c402114223aad9bdc5e5f67023eb45ca90a1f4bd342573340d3b6bfd1ed765768d77bb42d63385b6b1c1f62cd3bee211cc4d6a89dccf4354dbd3b521d9ea15cf275991bc7906f0d92a1e4b9ef96f4f916389fb6bf0f754b3108f81d030b84eebcd73c5c90b8cef0e6e6bde5754fa0d58a35dc94a8696ca1b61753c207bf00c8eb38f201dfe8b286a349ed8e9f2a5213b71b9267cda1a27aa29d45c26aecfceea8f5e356a244b649b8168719f5a955526dfe46f465319141ff271d26831e3caa0f29d21dae759a8567f47e20c9754aacae5350de9ac5d8982da19b39847468f97118ba3bd872f48055ab40a4c04642a620918480a79d5fca224339b1ab2967f6821deeea3507cb16cfaa38d0abfc19a818db100449e5293251593a2d51761f2a82c40a62f3cac843976ace076330504984e24b4e1e4128d3d5b9a9d48663e95f5deed8644e00b13806f0a82cfd6156c2606839c7926a290f4abb3f8058220293e7e8c7efc833c5197863e0c55a502c78004d561c0a7c89db7d69176145af4af7b35a05d3e2778ed452ea297b9c84c8973726588449d82fd05303f5dfd1551b12f41b39f1959fb8de1d033b178fef701d524d60fb412d715729866e5352faa95dc88c32bd73e5284899eaaa899a521056d90ee790dc2ed825564d9eea7fdec215e6aab709141c6cc3383750ef77b258e5d38a191ad8b40b8528455cf8f5db945a89911f58dc007fe7ec523a914988b382f478ac4deeb52b73f1fcbdf59cfec6dd102b7ef0f37c137d9b2c4f962fe5cb46f42a0b6aee9b7bbd3463b71819b170f3f70ce973ea5af68968ca72049635cf14e86bbd5a0a813e9172ebba546606bc5be80b6661f95bae4c85d1a5f4af4b06cf5380570a6a0eefe1f0270c99435b2c74e84d0115f2fc1e00d5a1ed044767a2c02f68941988ed4bb7b1e695fe7d65262b1041bf5cee70a3415c6b42f6036800c56c3c8324879f1b0b2b743fd9ed5ee6e30b9923d8523501b81327814e1f6f460662d213ddbfcd0446b6731b8f9384d453e9118936543c2d7f3e9b110837f5742c3c6a53f378998232c024237a56b6d935eaba42e862dc1c41f36316e54b1bf4100b2c2e01be4acee9896f81f106ca3b774f1674cdd4904ba86df89cb49e7f3edc90e5fb071815a0763dac95c94f5e694b3c07969ccbadffd398ddabef2032bbdb06f7dd68cbe032e194e27e45152f52e35ba5853d5648262351619f6c36acd1b6e4304779db2be85996;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h964be6b92cae53e9c09177dd315d9cb08f6a149cc2cdd5e7f7cdf29860f62e51ed2dd9494129733536d7516ab48d78f72b4fdedbf322bc717169355ea9dd33d4ec1a1a176c69301143939ff435c421b652455ee86c39fa7afd46edb029ae4143bdc128dbaf4b94c8a336a54745f2a6ddca60ce416603bc53988242ef6053b9680ace759c133bf6294f0004a527996381ef4300b0b5322b183edd81861bae7d86f66c351e5156ab7999a2c1673d99f1bfd0790c6d81417661bae421f7ca3f08376f58271ea25e13fdad91995ae9277106c062de1194381ad29f603ea90d76f64b927cee540e4fd081156cc3ea59b1da4282afbfc5a4ffc8ee28d0d60142e88b496c8b79541da48220ac8c0d479a72c2ac2c7502c06b16b266eff72ea57e9838a5034b5d080221b3956d716d57c70b44d9d881be91f76773760d4396261b8e185fc1bc34160615e71fe5128dd74c31c4fb5cf7c541812f6e4a65bc694358a3d75bcdcb3574d06251d3cc4fb6c65cb731322f125c2a407eb7a9303806c9ff96b218b6902167922ebefc16cf5d68353280b33432ac65640072ef0afab92864a82efe66550ca9bc23fb9297d85689e03838cf44e5ca78af1ae254ffb4b8fd7b43d801f111393a07937197bf37e2ac62443b8ca91c52981e1af24ae4366c99a00cfbe317c399331e8efe57756921b3b2720630c4a4fe9d46c43e45ac6b67a90968dd89a28ee7237ad3b58298afa25ec2b400a7ba67474dc4ae2eaaf5f9350177cd3534a4ab677d374c8ca570d0e127aab119dce3e0310ef1fc950d573940fbbd9cf50695f270e0151393495b0cb9f982ce9cc76b2888380e2491e3c5ebee14ff2bda49121b5be5f6bec1527c3d8043563cbf31e4fa947717f2027ebf0e61f3ebba525851019999ef07e4b63b020c6894ec26e5ae6aa09aece7abb9b107304ef7666269f5d37db9a9086d94dcb59ff0eb7c77e2afc1ad73787b6fcd5973b2734f673f1db03ef0810e33b0e85b9712b26b7f065444ab09993e7fa0e94ba7645aa4c53ea53774e901764e23e042dc35c7aab4af2cd5ac65de394241a3537533c9e1779624ec757d15d915747f21c2acd66060e5307888f915d728d4b6315be07f39b070f953b59cb1a877e34337b7756e5c2592cc0d77e0fbba85dec420136cc25ea9d642594c1e0c1e8f6a92daea1912a4a32aee4c3ef55b080e9650753cb2b6265919613217f01fb5b772d4113ca52f0e022630c7f774b638db8b81615db04917f4b9587f77219901ae383ed934687512a441a790ec7446b14db095bf3f6992d6eb81a6f0103e4efeafcc782ec3b33c3c13e26fb4bfaba073d9c38c31282a6f86d2862f4903288411a0b0f06717bdf70e7c71013ab587869f2f040947e65ea70506fa1c107e3a100b02bdee2d6979c0186e56cd9f1a4e4bc9122e75fb13c9c1825edb8b9f41ec94de4e2a4551c46e5010e4923dda8e12c7e3c1bea7cec1af0d9777763190d3c97951c07be8953d16249d332a45b2a852bb2526353eb968882db8763ad88bd85fdcd761217a196a7f80c973363e112ab87c96a5e13dc9518841ad750b5bd0de9fd6509c72f4780a4cde03c78be7da91b070c6e1423ef9d78acd7c7751bf0b4cdd9306cff4a297866bcd7f0433a183b85260fe1719ff1d51bb0c790ee1f01f56a58fbe2f4596d670ce5f3827b4e3f56611d7b14aa768531ea62da0552bc104281e9bcf6a9ee4bcfc6f1077125aebc11ede5abc3494eb2260b28477ff82e3805d042b065beb3db4bb547cf6f14eb4fafe8a63cfa93c7f7374a83187f02b4a2a69f63dd9876d58d6f60c7863df809bee98e2b1dc04a51eaf81ea3f900d85102803cf420899552f4130b86ae39da0fef3a4eaea022c78d124a6cd498c01c8c802e97b470fe82c0825156b0572e9dc9ae8b4d1642aeb2d07b9e0bb83ed1917635108bb39a0fd9d9be443676b54b8c6c6c8229f727868f0eb53579095f2bf9015bc4dfc6c41e2c611f94d264569ae9c4d158cb2d8d4433582ad99a330146f9d2968f03a0a827d51a1fcaa4514151d759fd78c26bbbed1df8afec810c03e3c7c140894e23891e69fd15b3fe2079a1445aef0ab9fbf8021136c5a536b0cfe4a29b304ce9a5b178815fdf3e5330b6bd7ba5fcae70fb99b234247621882f7e4261fe25819c217d6d5ae6b319e86a04c72029b508b61808a91ae2be1f7ebdba719d572285e85faa2c81e9f2f1bbbc738684b03f913edc1e401011c5c770477b3df78bd954d03766b5f5227f6c32b6768808bfc28f12a3758cea26628298802df15c4976410f75eb9e62f6982caea6d87ee3075511103bf9840053f3d89cd9454aec64323f77c4bed9cca719b38ffb6a81ce9ca93a15c04c474276d981274fcca893163c5e34b41e61d69ec42dba5ae866380370c3da150715338bccbc85dde83afdbb4cdfa6d645fa9720a150f6b9fa3a905b546522835f5b3e56bc1f9a400f080dc6a73ca5a614daf9f48b0bc309e1be087ce8334620621d44fa9d6deb14dcf9179d1868944523e23b14f8f1a3940a86aa15d86f1224c3a574445795b228bbfce7aec4a6054f705a913514d469b81be8ab197f8686e5607be766e01ec1cd650fd917e8ca65ee76d54f2fe71f0d6c0c5395fa453a4125f564c20fc4017395c521b23c3e49ad818c8bfcb04e81f0cf17d3f61228f6d512f0717c9c1c08588d41f2b10db671d9389f7a232461a2d5fc1d0e49510981166e048cfca1bf425c2919d7092a4132704475ff9f918f330ab4c63e365c6179ded9e8c5e49f18456e0d75c6e4137532043627e535d52dea823774335ddeda98dc01601d35cfdbc870c648606ce60b6e7e72bbc115084482c231dc9eb27bb963f4565a7253b9d14ba83188ea8f3fd03738cad4491512ce6470ce2186faf830b3c31c9a15f4cb35722fc1df4a95088e17d7062cdb67d91e3dc8745ee9c7cb301152568faf6a8efe13ba51a97db6b26b20706289e2aeadad8ef09638a10dc78ebca39723ef2d4298b167fbd072b58bc5705451f2f2cc844ed4007e8d7785ad683063a9575ba7f4a6896d9cee33645e02ace0938c1dcdcd0c68aed1a7f36548e768ed90ab2110d896cf3d1101487b45806da8c91fafc660bc489943e49c882751de872d963e9dda84cb97fc589a175dee78de4fbfe3e28061aae7923dca68e002cd4bb2c9329c8bc231242c0d016276e1f232f4ec017749bfc364a259e22767314a4fdaa0e5256acc5f01a963366bccaa40166040db58fa51d1d0904b61a71d35d7f827fcbbb19917a3542f8e3c071b74f22160e305412dadb9fa9ca7d534532ccf6337e077aa960caa09fa20c2c2f3ff9c9a076ca208f57839afd481784dae826318927b607448d00bf1eb48214510cc657048136f319c3782095369df70e240f595df818a5972ece6a946f2bfa4d4a3c216fdbb8b2c7e68523ea6b6c5d1fdfe5f717efa05ca4e1bec8657e6ba88565a780683b9be2d04f1ff141ab598c511f630c04d0e9281a61c111bc6d46fcdf6777fd541332c0625c65286dac99aa194c6936ade3e4bcf85ffd3fc20ec8f4c5efa7be719d0e8d25e916ea93584788e545a3bfa594369bae1fa361427bd9429acf0b2e0598faa8d69cc6f8ef0d97b767a588f204d9c772a1c3dbbcf70a16d652ce58d2cb09e1d72003142547d3161f281e75d5b048f56456ea900428297d5c15128fed8d7cc9912200896c76fcb0e316338cd80f17d3d7dea7b924bcc4bba6ad70237133a6e915f4b5fd4b471d9acfaeccd1ccf9450016dfdd22f8ecfb38dfb6f160f14e05ab126d11dd34ec6b9802520d5505843bcc790d49a7c3ac64800d992bde0d3d9d71edc5159309247c8fad48f24a651da877b90cb51747f56f05efec448928edd7a7cf505db11af417306ae9d5c6bb3ece7fb343f40f32195fdaedc85a76fe520bed641328a718b4373b69f9915877ed72b12e14dbd96298ff405ec4bb883353115a98f9cdf2efefffd0a3adfb4e587eecfdaa6af60626b3594db99061080c503e0f7a34cce5456fb7e7ccdb430d19477705873b8ec01e03e5bcb24e61576cf31b72702a0738c5d5e3cc972ac2bdbf5b352a8aab8f1637c869e7f2e1a510c21883e1288f002fe9a3b807d30af58b09ad9d836cf08d18fe3d8f2e5cb83866e676de69851758e83fb542f6e70d5ea3a6ae068ab7d24c021500b3e83c0fd85a02351da9e8f55983d4f63eec58f70a61a9eafd070dee77478fdfe873b54e33cf2603d31ca80ef76f90504f07630014694a56bdbd5f7fc62ba5b58978210b84d8785bd0793dce8716535c836914071ebfb9352306b0a604c2ae44780a7a5cf03b18fdf624516b295c901f6e23a4315c30317f9a6b1375265b7d333d4b71a4cf7b3fe435f5df8970d5017ccd620cce550d15b763a3fd6923d8f9035daeed4986f5f939d487f19eb2f39c870441752c2676eaca600dbc752b93f8a90ef095841f72b1e70a6de97b799a90498ba6b1c53e8d9d1d98e544d8fc881da632122accaf96bc8b6236816fa497dc7863bddd99b5bb75e717fed390e1bec55e275a03ae248f759bde7855aa39e20b267fa82e1723647dcd86ef62f64e89dd2ee783076a4bc64a963e14f8d181b436c13f2c92535a7047eb1abf1c76d1f9ecc3f3a2f96b4bac931f35d4526643ae2797daa39b03862cf2cfd1dc8174fe17696bb278fe543fe6596324cc19f7d9321af864d43623b003d9657691bfdac8253b30d10286537853005ca523b97d17b630468a136103b63fe06f652ad31d945cdc9be3786a940fbf1e798d3ddecea747fbd24b55027d84e7d7a5266a9db378e462888040ffd340a97176e3b1333bd70fcd22fe098acffe1b9ff38f5bb30371a3e251b60b99e3a9b3676204333bf7742844fe9f62d06dfa383773f567b0e7157c0eccc752c0f6f54862303ea774a57375820db45f1a727f0272b4f0277ab01a927251a27cb622f736f885da71fbd16c2c5923bcd146ecfbe5f20e5cd13968eb476092929fe3f41e292f6408a75a934d9a51f4029fc7ad98ce17de2c2dd3f39741576bf78df54969662fb7a4f323c6fc8ef9ad6219daf2d8cf754e4340458a3b51054572a9f8152d469ea4d5d9523f4407fe3bbf30f4a2bab424c2f4064e3b6120c0ae925d7e226ef1c6404c008e9db354c9afd9792a0812d3222b46fe18195cf7243ccbc2ffb0a2f06092f9d95f9f66f512c8b9c1a3cd46aa397aa8c9b5148b050cf05bfe8d1479a63bcef275e4f31e296d8e675a66f05c7b5ff026099d81d352a890f1251aaf2e341597fbb6f70a4280da4162b5f6ac0d68337ba2b229340f93af82f7d52cd9902b57a5f53a92f7b5a258cc165c10add825036c23d225edde4c25f385b202478b487b9ed86a86b049ab3f312bf38b0e88619273f3a5bde7bdb8ac25b8d37802655fe343afcdd87e09040056dac48080778e1a8671a66f6ad0d3c20feac8614f1824d353e81247b28537a3ff6d2640dac311c45509796fe4d9fda9039894127243d4a67a3a3300839351f573dbb4564bfebd8675c92e133fb6d42aa0343c66abb9c61d49ef25164f566d9a11d109781407830ac637db5d3a8d194e88ab82f32d06b7abbb7ea692b1bee0c510427863a2a10aa87e4a5445c6cc5bb8d4c34b93c786746630fae805766aaf479d7cbbbd0894ee5c6b2f8c5d9cf38b73314cfc05c7b35cca56384140ad32b00d3286b94c301a5f90be5fb37994efc473275bc535b1eea0e646c4bcce4674f514fc368cf1a3955bd805978fff39e048d2fbedc30c81c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h95d155484465c3315e45f70bae877e45c7890b8378d3f5cb2f7b3b289862bd24c1f872e9d8cad30c5d64bae8f1673062c68c30bf3b6db08b52572d8a4fba279ac1704c9654d6a61d525a1e0033da3df1639e592b9fa431c7f5a4119fb7af09593221e1bdb1e3b309889669282a0cc9f84fc85c59ea7e62f1199f6bf899f4809a923eb87acd2561f77a6e77203f6ff20c069e333e3bf9f912a86293aa138aa0f20f5d07fc112a0c2606b6b45ea8f704c4d0b446e2ad2dcba7e79978b5f9c3cb1cfa65e3ee6e24ba1ea91c2cbc354f493ea58c3acd6bec88a9b131efa7102542f4280fad441b59fb04ddb8a0b2af97ee11bf17cfa149a2226e1fb41406da23db3638e747d7d276a2d1fafdbeadf908cb2e780e92593483eecad0b663a5d9e4865a77cba6394dad8d06d02acc83b9b63bb1c91b90b8d3bc15db4d9111f2dc03aaf4edf65a02433c2f40bfc20245883ba6be6f250aeb821f8240fed07358e457b029445785ade0f7b99cd1fd37364d09a0651f7c59c0357fc862c3f8505bd9db5364bdd89b6e41e04c0f31f9f64e711dfb0ddf9e79f691449aa2d1547c92b42540fd675c2b6dd95d8a9a65d035d079b0860679fc2b99792bd073ff36855ecf550ec8048bbbb6e007bdf48889458531b9bfe0e2c2ac2e614ce84820183741e8529cf4d90a0faaf6af3565c7a13c3a8838691bd4830945b2acf084f691694427b9280a96c32448adbf6d05c129abccdd5c77c9c14a262bfdaabbf3131f38aaef9c044200392f0a0a754bbeeb4dd42a6d7642953b28d3eb3d38722c79cfdd192cdbe2821d075af012bed801b5ef4c86f7a99c6085a7686ba429b87a925dd6c274dc8da322046b4a43a487f45df49d92f4e99b02148324470fb2cb7021adec7a2afad064f7e908e6b9122bebc1b19ee3cd144668c0e1a2451842509445eaaaeb509d34f9e7f7c5234b5c1c9df90576d5e64e79e87bf3dd00433f78525f68b193863f7bd699efa78774147841379e917307936e57351baf92f2d9c2f7169caef27727fbec3a95f5c7c6fce5ba82a6b09924cca14a1337cdb02f00371ae075738d586c9aed6e40a1d73434e4d201385d419ac9d7b5f1eeb17ae055d4f2180729879c95d05c216d4dd34b357b148b004dcd088264a496b3a77760aa88978d24d1202f9cfbe619e910d883f5baf4d05636f0e4141c72ecf2d4ed2ed8113b7f93352b9e55d2ea848da3a312f8f98231a4a08c215afeac0fb20f951da3e7170e5849cc62b89559cf51ddc9c9fe98ca39bde59328d2557d6da3ffdc249a70ec09784a7c58bcc26b3eb65828f5e86b89bd6fdaa888d45bfb391bcf80aaa19f398d755a60d3d16870026431635c79184239099094ae1d3907eb9bfd58d0c2bb63c741279d9c9d110dcec96b6c354e39f874a253a85f985b90c51fef1c3a7aef4f5a72e80c2420124d5fd02f14c86461c320d21106d7a07431edd8de2f2e74a341764672cda2f598a2d57893d1dac51b2a314a79ea57abee8d62773eb1ff07e1279a057a5704f4de6f3e0788d55f7249799c471a89fc8b9cdb34e53b953abafcb534ce051b1a496f378e6d7bdd08830c5dbc393a4f604a213434df990d3c6496a45d2190f815e3f720a676d6a4c155fe066e2497793a3d1cbe5862e1d751191daed44b009550773543c5aa422c4b1db0361e1202979fae17af3ef58783738a0b9be760f59ad9050d1e2e1464439cbd1f81d85d68f1824070a507adf84305460e71ebaf8d2ebad4d09a913eab146f011c99bb77010ea07366f5269649308da1c0bfd61d4cb0136330f23ca37e6ae985e26c01cbc34fe0ebf9dce829f5b368522d3dad8cc698af8a976647ac91f0e5a0bb998731605164591ccf12fff3e4c8c66f4a0d6142d1d6064e28892f321d9ca8c47c5a87fd9e33e30ff559f30e13121829f6e49e6e8d8206f907a68cb4ba398b47cbb165e58b6b9f3a84428015772028e96c20a91bfd7fe565d6599d480a764d15d174762ee216d1b46c42e0c52ffd3bf8cfdcc3eee7722f13c3ce988c7562fededeb8ffe00835ab1ec5969c7e9661e5a2edbd919ba0bec8d40c9d08831d8b0def0e19a5183fe88bbba2621fd6f8b11f6f0a57049960c103bc684ed0d49ad21e72761cc173814440b3f0997f308d9e56055326328308fd80a4a095f892a795ba33f189fd0122080c1322c9b496e53cfcd07e91adbc467c473bf20688a25ff6105957b14a09ff0528044067079c59bee7d83a8407532545e10060bc895e960b2022987ca8b8e73e55856b4fc8437dc915e4dd7dd6f34c53968e0a97a94ce6cac33309ae547513ece4b658decb799a470860ccc425444f8749695aad9ff3a817bdcf0d97b90e473cd1c9dd2f39dc897e7fb0e93fb1adf319c0d88e1d76e0797db8ecafbd0d8c14ed45ede559dbc1f9c55c9853f0d137d6adbfe043c78af65a56d30c85d139e74b1299efc4d27c46afe7b6ca0c341eec0f22f932d9b1e650525670269bbe3284f0f0514b6a5dbec4efeb449143507b0b7d648da4632f4d2263d21d62611f72f5dde23601521ca20e751468ea2c9787393d7d47b137e37ae204c1eaff4616ef73ef526ce447b5a01894df01ae8a66a4b3a28fdadbd27a0fd298b175b4bde07f87d78b1bfc1865020f6c482446fe5c9f8a7ab9358e28c5fa4bca1732af3375173d027105e16311eab72b6f8c5c3bd6ce1fdbd72f6f24e87f4ce55bed948ed6d81b7be4957eedfa9c050dc1615718873138154a9372565559412a4a61c8d7a5d3c47c16623638fb696d44912bc9435ecff02dbdff56550b613799493b49691a0e6307819782de6c824d58e06890d228bc4f2c59321c6644f4c833e78ab68caafba9713da99aaa127349c20487b035c13fbec97387977279669b609344deb4f02e87fb3fd2b2a11cdda15066168d6a4d09864d316ba17118e75a2e53f896429e6281ef7a98a06ace9bf5d2c63e86eb2faf3abe6fc63cc3f86674f1a0474cbfe332c3953e84850ca5f35119a42d643892db714e68cd52e2de1e0d8e0f708d05afc887d6cd7895fb9054e2f64396a17e052f3b0a6b38e3a1ed1d8980e31c9b0b2c10ee91846877deb120cbcb84f92a1bf81104746fe4abb5a2b3c8d571659153a839f1f1dc5d12fcbd9095f138ee97aa1eecdd0b31f1d6af7ba1178557f87cc47cb2a4cc80544b88a079f7ab7651cfcd1ef4ef92096836b7598a9f7e10dd6a665b7984110a25ea022bf40a1f80d3fd26f3cad531a8839e54e4136ab6e749cf70cee0a2b447b5c3982272662b91b637332757a4f85c7effc84ce5b5d89b8c9182c76406532a980a3a77e5d55409df86554ec02bd97d04b9da8daafcd62de102599f0c2a00ccec1c7b32da0a0e02067baa6220b59b8029b5789f4acca017a4c5a0ae56c2d049fee5d9c39c01bcd5e4cf28ecd3416f3d940bb32a2645cec93673afe54b45f60d2e8586033cd8bd8a93e277a303d09632936db7d063520d6ddd839addf80f59654822eae12f5d7f0d00641210d315441fa2a8028fb4d654ceef511bb51fb7597f780187b6464cf756653b01e0e0ae27c2b49f9ea06dfa79f43d4e5c6952f2587bb23ddc94aef3edc3ba9fe981a2b43fdc57c29288fc5992afa561e2eb5c3e432e2006c5613916bdf7bfb7c78e28c56f13c1857664f6b1e82502e76ad9e1453c04da426b26624284fe12828f400e5dbab992dfae75ba72b3c1f751b3287a471b0a32e693adc06ab6ba97aff79ddd2ca6a372fd57e539465c36352935b6ed01f6062943b0ec2c4cfa87278fb7215969be5611010acd09a6b5d38e5e30e62103908f745c4aeeb4dc1796732cb084d35ddec10fed811d303c1d018b9eb3416cd4d3e943453b94330072c08b33d3cc20bb94929dab0a1b3da55bb687c4d4d2aebd6ed7d76ffd394f878ac4ef2248936e1da87245008f3736f26ba18264936ce33285b01a5d57bcb123db30c32353a7bfbd4ae812129049525e88511f237ebb6fdaa3eeac0f23439db0cc8685e459174c409f90d941158d24f2325d602ff61c8ee091f99e5b0d64438a6faf60911af13cb883ca5c23ea8b3aac41de38572e36154af47689e909f1e8a9aae2bb9ec20477d35d781bf0d3f8a158966f82a35e77d6aea110c9303e19743290d54ba44a98e3a87c78da17172ab3ab9833f0cad305cc8aa961909ad58ae6fabde1eb5cb59048c8f7fde407ee2921ea69206761f0a5705ad871c6dae5d661739d5a496e44d1508b6232054cc1eb2364b32df230f352048c00bdadcf1a5bad496c54ffe9a6fe022d36dc8e65750b37577bc7d870ad80a7f231802a76b536fd06c5605226db172c6b1cbbcd2710f0c24813e337aebe21a0f93e8c138350e7f8cf42d3449e8ab7cf443809572b8295396d51eb4ea013e09ed9de6eb54de3e02007031ef60b335c0a849e1032f5760cafe265a4b400309ef09e2e0c27f435edca4b9350a3e82d8d38daa814df269f945283227a63f337bc8bf38f86d2076f2757f115c2bec60f8c5b48bf68360e88e8f579b85afde9b498d5ab211753adb13ade8a3e5334ca06a4057bc6fef333a961e385a32e73f36135ae6f87a6ca38cae8db639d4ed363507bf6e8d1db18659a6d859dc3a123353b585bcbb4e582e51ff6730a8893b95f60f03abed3a8ea57519e0c6a3cda9650a4dc808fec75dafd19bcd4003f3634e0af723a5a076822429bc6ff584cd5a1d760cb682237445108f9f1fd3020ae2db389b8ef722e3c647df65ea4f25054a18b54c7fffb4ca3649039cc03eb1f4935f0a7a6b224c18c994ea24c22dfcb9fe0e4ed5b9de35f627d3ca90d1636f7982f32373d30387fb35dbbe4eb6e774464939a456cd69eac19e0973d7a726788581aefaf633196d5b3cbd23bef511aa6093c549fc9cd74c922e69c0fb997a62adc669fef017ba6169b56f6bfaee4bd5e340047b0953190e26cd2c1ce5226f24db29ab46c972fa5c86fb2cd3de9c09a905fa7fa9f9e85f433cc0d13552f6f529b0ee9fa1df57d776277bf9c301b5b18cff5133da708e721590056bc19c12fc405a0b856cc6a70de237e7d5c52e92c72f1670b6362c65506e083c8dbfebe8b8b1a899f6e6ae4bce469ae78510056955371bf3ed5f7b7cfe2321a3810dc74e7c7228d89ea5a007158de1d04eb1837878e1bc5ea9ac5cb84650f2d425e9824c1baddff3a89ab7b14da059b88546407f8c9f4654cedae8982b1c3adb81ee40f4ca970cf338a95728afdbd60db39e0fd02f5d6ea604cb30259211f8c9adb46ee08f851f0c25689f7f6126ad9a29f94305256f2ee6c2c993e904ef4c033b9795538a76efc3a92ebe669a1653357a2cac197a66a8edec815e6303f323699e05f262094bab8729efeedcc0e047c30c77e0cf770674454ca1e2cf35c6f8434f29cf06fe5a51b2707bc1b122c450c18bf1167b360b848ce02ff500de0c66750c2d015fa46b5748f7647fb85026089745b79e630601a9538cc4f79ab2d2a64023a555bf0c0476f8243190aa977ec101904b7a58a95096b307a8ed92f1d33a5bf707dcf7bf28ce44f35ed94f49638b54cfb5fe5c98f780c80068b3053fa8b2a0b5bd65d01968296053f4b17d6731ceae0d414926f4371d6ee06c011472d64bce010221655eeeb4558600793e56430f070d58dda9910e1f31fc186ed4ed236fa21791246f3a82c5d5be31b98b388e40f3b12f525c5fd2ac3f37de0145a47ebf095ac13c04f12bb9a478402b08db6391151f55faaec4af4710ae2bc3b4b3fb4d168123fe0e806cf4527d35248af06a682fdf576;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf60c2b29baedcd93e4d4dd35b41313e6e928b19a3b6a8956599b0a0b3bb02b6e72a14c323cd09a69f5994cf9acbf51f9924d37516beffa023b2411c41081e6718f69344e86805db6502660f2faefb6cc48c2208c9d2b37d82cc840caed58c55c9e82b8e88b548e2c075db63730cc70da86fe4771d47ec58c5a9ea9317a6135d3474bee956b7ce8bef452a036f76a231264e50e73f404b02a8c50e42c98dfccdf55f7ee6224f229ab8fb42854d5d2060b6236492a512add5d2dea1a54304eccb46f01445da2028a2eaaac8fbbc967a796cfde28d803314fc83d3c737cdd81b42a210430cc5f10926993fa48180222f367c1b5a8549e0f445e919518f5fd4a535f660ee0aedf765608e33f264798c9a125238b024b92f59a8db57b0dc1135713937576cf512c5caa050e2e55102c9532138be87790d40771edb2fdb869ccd631f4baf9a2a97c041dc5e97489b4bd25def6edbadbab6921a95f5aa08965a3973577dd4c9bb392b02d33ba3bbbcfdd22e843d42eb2051900e20144d1c05d5ce77bb074b03a6756d0006de18a3258af68ffb9b7a3ccdf60633d05c661c4072e9f8d66a1b558c079dd55768a5e674813be09bbd8d27bf1d1f969906caf90cd94c1cd46a74d260ffe5adbaebcce44bb9376112da06ff1291390691704817de98b982605cb47a4ff0ff1134731ee23e07823441b51bd56b5b4dfcf15c2e5f614635b023efd80ae96aa73d7b3762b0ae3cd3cdd3305ef39971d02dfae244a3d1a4662f5f047728ca1a7c65e6be91ffd2fb7dc8517807162c12468b42ad788ff6da1298f6e70960869684eb74c7fe9bf7c2d603583153d8f811b418fff3121b27fceb7c59ae920a0fa15a9119494f90b906c128d52baeb57d62a56130a61e9412c8ee29b498eba82bddfc8a80650356ef5d8d7d9dc33802d3dc352c9436cc55a51f81aeffe6208d06e3d305ba73c716dec466c3bd4115717948520a81d7428527f7a4dc00ec78bc2dbbd7953729710ce6fc5aaf300da38f6c85051a56e3be60cbbeb8118fef59a557096720200e89b9454e18e9ba3a3667fc2444aa26d67e8f35b622fb56f8bab5811fe06f654f0d2261f2864424790bb71d537f8179b2b4dcf8ea74c88b521a08a5febbbf9da422a3b245c975769af2cfcfa6b4c030b37480d2eeba97b842056db6689bbe774c40d7611195845b2c0b328e1bc793e083b07e7dbba8cd78e5684b5790a0b1c8beed45bea8ca807c8e9e9451187d364123441be073d66574ddba5e34091fc7c4ffbbcc2088abc27014777b1970cb6d901e1a4d80c53a181e866d7812b2fa1b403113f7467693d868e0ddc7827b5a1e8eb4db8181167b19bf361363a9c4f37e67c337e19a47cc6102359fa184a380cdda6473d92a03863a094c239318bc8b6bfe2b06a7728587f4db84f0b9569e67361a181c7d0549b24202bc4d2515b84e1455788444b82beed7baa4203a7bfcf14bdf35c204bdd33e1e5f2cd13318703c12f81425be5ca45634ae9974aff1b429d776942672b60c5497411dd295ce37febfbd21645be7ff3fd8faae7591b1d3b3d282d524182fe71b526c154d772438bf041c73f0998b13dd8c689b2ea8c37853da0173f63bb3550fd24a4bb47236789721c7edba1a468f17e38d54370b091ee6282fd58da6bca60efe1c637d143040d66a629347f8c2a8e8f9a6651adc6a4cdaf4d8eb0df9bd80ad3276a18aecd2bbbd7cee0053af667be9d54c184b59b978156d182e7a43c5a7353f42c23da6b8116af71097cf97136411a6355edc559980c0be030c9117247a4533fec450a944699cad3c6d6fa440c79b2cb62b9f90065fcba819c22a22d29d82e78fa56e1358929a7d009f5f86c377dedfedc21fd1781646e8a96c9e10dbd8985e4d7bbc80f08a68297723a713f5e4285b3abaca617bbf876e7cbdbc1393d81c5a8fdb2f7cdfbf6c1e01f3824dd371b54641e158cbcc1441254edb9f0fdcaf6fc5e44d28f7fbef4c7ad13252bd1ba46de4533baa1e79aab8ff2c1fae5b07592e8e2fae947ee583220a36159865a8890b82211afa2609fe3c16a846c5366fcb14795954eb5ca5e36e08d2c1ae9d3fe1ce4771bb6c9554e1034393ee7ed6e964730b3df85f41d2c080f6c5b76e73b66d2bc9d325ccb54e839ce2c9b349001bd5d118bf796ecf2d8025a2e188d462abeaee7670bd2c28f7f9e5fefbcdd6e8b6cee025362c673c276a9d21c5bca6156db04824501619f540a255b5d3ab92763e8e701f816fea7b2d40a184cbe34d2cb7cdf8902eb2d32ff240e73332e7c70a9c69544473c24c2b5620669ad54075d9decc48a1f203b0fc4441e64be493c933d847a70db05b893695102495495613efc8d1c41b13cb79b59a9ebf8451929a36b6eea638a0593ca8442e70ee8392f145e6c3679558ca90809baaf09334abd02767d2a0b419d859abba0884b4ab9fb37c2be1b9bbb0b6a21eada9567204fed470db38fcd3209f4757257d3b7fe8aa99368bdab9cbe986be96ec156aa7fdd4d4ace90708c26df019c22d3eb216e52985256367360fb338a39ad568551b37195229239886645eedc737decc755b83d7c42bc4df04a9728bca67f5232985da41571cab41489827721f48cf3b3bf96b1c5593aa5fa9a6eaea49ba6f5aba3b765824a8d0bdff44c60a9d58602cfc1b4f95a8d31818e14d6a2a892ff981753c69c1232e0d4acf0963f72d3a7def7614ee20e9f73878b98d49c5fdae399dccea8ce0b4cdd244b5687f4c935299eb768a7ce19de938249c4ce5f900bf06c7802ce9eb6c870377a52f39df2774d4ad7ba34f6af86e749d618b7b6b69a97384793032c9666d8f4cdf204e710b4d4e91973250f3e1b03204e84df6ea15c2af39ed2bd1c298857ad8ae1241fe13fcee049de7789b639f5081c776e1d71ae6eb284eae494127ecdb4ba52230070daf285fb59dfcb691ebbbeaaf660f8e3aa5174c01f81769faeb69d08b7349a1ac014d199d903919c808d9f3f9187c18110f88312147202f88c3b67234eec4ef462964fc8d1587af06953f4dca0c9623376453dbee84d42247e6637aed69ab2c53e55085e83285d3f8e10ffc08e5db6f0acaa91b0c3c7f554191dd1f01cb5b3c8546ec1c40639324d24455d27078a7aaa41ef768271d93effdf56f9d07a08ec49a738971ca266f7e8aa1573117d1fbf27c95aa68bb7746d79711f1a687c3581b45c03b1301d3fe20cb0b58290b53031e4f404177c3c537a8398f0399dc079c5c7cbbd417abfb59312e20fcc42e9cd41cf83a791c41e3df34f7faf398f05183baa46adfef72cd0452ac2a50588d8baaa0cf48d0ab8de72b7ecffc2cbc5eb72b5a0bbf770243b83971684b6c460914e5d8ce4793443a1e32076e6aafd7224534a0042879d5a0a588a5ac5b4c8c9a6e437ec232af2a19caeeff2096d271d90aa7671b44a2dba3147bcdfa7485079b7c21a9a7cc2384bc92db751a868816c55a640edf9f23f0bff1924f3e8cee96ae628d9fb09e12e410d737d96f3004443203641f866da5cc4ac65f2395ed3cb22b1861f81cb6f450fb0a5f303140191dc5417b08a06148898ae3581ddf2fd2ef78224493cffa36f0d4b6eabf985fa35bdbbff718d96e5217bd869d875e813cbd6f05ecf25115a792d7b3430301d7ef6a1d6a9b80acc04174852f7bd25f8bb74b96fa510ddb28d068f23edbbaba1144bd8c8510cfef4ef01ea9c0c8f94ef5b939e3d9b0f3967f90850386e0e45fbfd056ce09377f80f903ef4a416c765388a42b10d861952de88d8be65c795111d5847db7644df4377f196e361cdbd188c20e074833eb48cee015ef5900b743f3ffd2f04db915353771d8ecf0231afd863d90fefb3c829877a1608752bc93d703fe81513f0bf20f64126219d43018a3e999170924ef128b6690c9b5c5614d83797d282f21ea294e01e863c093c28329cea009b59b12496fe4bc84a01a2aa6fe7f13aadf68a41534daa7a85dbfdeb11ae2bcb1378f9d4d626f7c97d58a12b77e9f24748299ca59274d8b9da9d9638839d9872e496e9f456f0e43fb339697df364a098dfc2e515330a60b71cc0aeb228c2405247352d90c76d1c391fd4d172d94330544ea3586350896d93b66d27e56c031e74e5e06ddd7c6346f07881c9190923210b212610e13b54f70e69320f323fe0d2f5cf38fd745069fc5106efe31b34d1f1c2c619938eaedff09f5c62cabe568490707d058581b189e8a817f729f8c70e5afc34fb0ca534710cedf870742a19868250c0d737609540ab0976ba5578d6359e3ef710d770b1a8d7597d81b512550817a094ba7622bcfbabd77f25e9655fc547d60351ceb6af896ec90e4ec87a4afd8f3d1cafb623d689f65113ad2403848a1a08c42271a6d18ad0ac7d588f2fbc8e2c3e87c65fa1293d7d6a26bc5e182618777e214bf88bafd9bec5982dd05e40512c69f77eca364ded8ed618d6c4102ffe1d6f70e1cd68e96babcaf5c23cc5b7b6fc0863392f396572b15fef941b8d0eae59282f1a51baf405d751fd47ec5dda8b77182ffb47d106662e2bdb3080baaa09fabc27c2d3cf8f90b60689bbf8a33b0ddc22a4c53f96ca6989f8f73d65d0942a87d97f0a03c8af4311f1715ccb7738821549a75c30dcd3fcc51b1a884028df234baacdf8332b4666ac7320c2347440105da467b0b25de258f30a81b8534ea9f195dfde15a04254d7eb7479a294acad7c48f71edd99f51b8a40c6a9112bd82255e8f10043613904e601bcf750474b523f12be97bc4cb7bca2b8b40a1c29c110cbad33154f4f5644406434da1dbc18eba283169f371cd82ff420a7a36a4ec0080cc9d59b7a1ad94fcfcc1f4143d71bb22ef3677ccbe82862edc153f8a1188896ab9dd1bea903f56044dde4e0715e9c29d0e77aae9ab4e47e7f8432c496ae4f6784c398ed26caa06411da4711d88a1fc50cd664d8b27d905dc8544429a264d63553b7587ae64184ba852701c892c8c1fc0ff69522b4d4738817974f2fc4a2beb9c663d0759ac091f8d0dc3a9b9633cf1bc6520dfca0b3e4bfb9abf84bba5a3a54f701459733dfc644665375eb80383351ec3e9ffec6124b244d65dd156c2aab630a81072611ec099b7851a5b86d7c5be9b8f536dcd89a3361fb15c138930e7677276540628fe13b877ac59fd5842bc6c4eac580f3d65a54b6ec91259b789346678615f29e9d6d7c223ec37c6c52e034b1a6a04b4f984d9662ed5d014ccee67c3beb33c50ea9096e9a8ffc80dae9e4f0b79844f855336013961228310b5d42b1aaadd4544aaa2da9f15f842fe44126f9a919b5e608748e336df708a1baf8f958d174eaee730bb9c24d77e2d165b05688e86668983b1d216397ee48fe4d2ec9814496c4757b0e54ad13dc6de9856bad20bcaae912e8c6627f01277188bb1e2bc22ccab18af347e31cdfe456038bccbabfaad3225b4399e808e38a21bce9ef806bb082dc7ef3fd58ec70038bc0e85f4c81d78d0e347875c823ce810a8be5f4e046ad4365a9d4558bda2f39a9b6dfd57f9dd61f61b51c9f350a5dfc5a488cb147cb477653dc6de2eab0901021fea71a2ccf5948d2c530bb69e4b9a9bf1abae282445142a147f99fa4d1ee4cd5bf077a0fb80957b49a327f20cab6d374983308e9b2e3bfb4453977fc2173916e791fe4f2c981fae0955a4dcf06e3c03b12ccb4aacf7820e4a7bf53b612c5d86668585b34d118812299fa1b349178680272d4464bb6cba7f20e8c1d650ecc0b4592d6f840c9eaad0eb170a44e1c5a4560bb98c6bd18cd045310937d22d2d4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha62aa8590b6657404b30a8a6590f94cfb5d1bca458d640f344114584a8570b76b6ef47541126996b057cd6e1fa1172882ab757f48b3704ebdf2dd51b3659e9c36bd3ccb1013104abc9bdc4f62cd9e897ca186c03cf7dfb14e98ec5aee003bb51a422c03a070183dc3fccd111150bba61736f34b4f885a5177cf130ef1297bec1c6634e1e67e90fc5bfa65be04a1e28b3e5d455084d86ce13707e7a62de8c30a793177b85cef201d749af2b726bc66fe20796895ebf6b8d2659ce36062adc5d81e1ff234c115fcc2ec25eb12d745924757401cb07160983e67f3a16c625eca944b3a6026db6d6cde0c4aea99df6211cbfaedbf994456966d713f5f66e3cf6bff71db71e2e6463ac7c2d8c7fdd98ad29a0a6afc89ab4fae08d7e9c4aa059370f67801f0652b79df06683ae54d7ba42d10b2ce2c601b35fbd1a271234b2ee4d55bc5049d99b672d7a681e6ef547ddc8f303c083c2f1807cb92ff84f3a86c770d835a9b4ed6a1f6fa362f98936dd9464bc13a05e0b4000af11f01619330f65a3c63d332064763aedd07e94f63ef37ed23a3a7f42d68e9c112ed0d071b631f534c51d41bddf7eb86b6be5ff2ab27d5bd10597bdaa13310e8faa204d33acb7100459025e36ddee4835a8ee50956b784759ae39063e72be074f25016dd7656247066115ec27e787c958051a064d40f80e4bd20b7aed40b3c527682ac2b55f761e970c9a294561c241e4813b0185a0ff1008dc3faae18fd7f999002a8f5a88297cd979f74c647bd6a883e344d13e5560377ec019502ad422af6534aca74c814e922bbe1a466a19a7b1b1cef9c2e47176ff79c4b0ca76f8bc4560bf741d6ebcf1e4be006efc40979dc6bf1c513f96a642c02b925ab6f2c19aab320a59223e3ff56b66f8f9cd4d9824faf4a92b849ff5d0b469228c3b7d448aff30c9f6d132c83bd9ba8ef6a241d65552dc6fc81e40585d9047f365869d2bac871b03f93176531c17d0492f9df73dd92e55a7e838624934112b283245d3cf6c0b58dff288556819419e57f5b95acb336254bee02cfd7da88dfd883fccd892d2d656be60ed241157b6c6803ab7440e129ef5db117b7e94a7b422d957d08fa9a3e6ba0f91b63faec4cded930d815129bcd9b29d5b98e765303ee922f9c2e206e163ddc75795e883f953da406cababd125e1c0710c444db98f40f3b42261cc7520a07e4abaee1307516456056e9b7d3b48fc88407832aa4d89182b3ba575ce751e064e3b2a5bd1d1647f3c6d996cae809c08e348822e0438b28271ee1efbc6d29b0485f3d43dd4393b94241dbb4a11351a73f2692494d379c93926810cf35ad59bba1c2333af16617b3aa11e2af606cbed34eab6f7a2a0246b2ca64ab574aa6e6bef0b4aa0f8ff9aaaf424c1b120ad72ddb2dc676bce43e397bdb546247ee2e062220ef6b3643039053994e9044481b8d19aaf045142db1ba8cf8a0ff64aaab4a5aed58a54e335d7fefb07c4a2c6fff0e2d8cd02139161e9314ed9d569bcc4b0f1174cbe95c0f23eaa04b68ccbdc4f48bf5235d067cf16a3766ee891ad74a194d49e4850a1a180b18baed5e7be601138e646b8c3a75fdbd36876e2e5da33c30fe4c3048a1df314dc14ea21db96d6b200c925414ed0a03e0c77e23fb375fa1c6217eb2709bc4def0bbf7e8c4b457362ac815bbdfa330b51c7db9c837c664087d3189dc651ca005ff810e1ebc194f7c4470ccf114a9aab6411ee1f3c4c5c1322944f19c3719171ef7bd168851976db15852e484b7d980ba23d157cc672a3902ee1381171a2af0ac7cc5d850c14f31c7cddd2cc531f41e070c6d24f19283d60fcd2a79b4947fe6fba276aa3ae8dd3c59548a9b70e079f324d1485119ee041689c0c4a29c58009269c51ac06d357e3e5f8761df4423e5f4443394acb9c919ce10712b3738001c472a603bdb6b1f0f36f80c81e1f1acf2c3f5dd38b3500f8623d1d4a686858e7c4175838edf0215066dbd97d962d5f8eb442b9acae22c590028c71281ed7d104520a09b11d3e97bf62c9c13c39702ffaf28f6928502b27f67fb53a1ea5d528c8e714df4977c8914cdd695d78f5189d56c2008023acd01972bb65737a82781e5ad8c992f167ba8a5e7b61058297ff0a81767939dc88b8be431230a64e6fb13aa693cbec4c21b912f768fc2b782bc9c413310816d736b3d62e9e4752631fd4eb0a246c1d50be67c72311826beb7b6ae4f4dd8b9e54ab5ea8dafa441a77a1fd5139a9c01fc15178f4bd890fc7e1e52d4c6ffdefdc6579f067f0389bb5d31e6f85fe30dab960cf5a8c0c6f13b112f919c8ec04cac59a1e0eba9dd5c60f7bd087260807b2ce122c38cf481ce7c98cbee3ae6e9e29e0b159e28c28eed6f5b5152baa39b30bd19757e7a513c3ca0e26a0252b2cd35edd2c4754e586238af6c5a20c5f7c14547aa851ebfb2553cfd670b9d45ba5b6e9383259e58108b3e350d2ad5206d51c5c71252dd7a610630a49c8df0586b7d91a3f4fc00d3517dfcb5aa201b75787122450bf6e97640f9f79a2b2f672f0194058d1532e42eb592af9be477e26db2c552679420ceb3822401e479ca160f65e646eba116aa9c6464998c77985dc6e3b8b54d66f81b344a28cd06e7350cccf2e1f93532c8d33b4e858484a9ecb90255ac5e4736644962e6f2fb3dcd32c0eafed22a0ac7aa8852e715baa2c02f323233aca007c6b5eb8adcbe8d93e8526f04ee053f9b23b4bebc70d3faf74faa69c5834aed3f588b36d10dc850602d4d198a45a86ed354f6ae91a901a14e4406f60de879687fb027e2a64f7f167df5fa791adf9cc5f4f099ff0d70f67df11a272ee6894dee6b608a4e56b6e1bbca4fefffe3bd1952802e000b7af42203942887d77026469421732b9d1261365015205586af1afc22ecda46bd528772dd8e347e2d021540e6028d85d4880d39b073d63aec0d6a62b798a5120a606178ddb2bada899ba71a55b4ba234be1b1bb01dbeee16ac04cdb7858baf9c1eecda7ab7c2e4a0a0ea8cdb2ffe2e5c60db11b788c4f125cbd39428a25478ceff3c2b30735ab89df85452993a283efd222951e9d4758607705fb8d1aa6bc18eb84f4f6e6abb9a345063dc5b6047f4ecb5fcf07aaea29a4b9d68efd0f792ae1c68c459dbb3cc3606c712626f1bf3e8e4ddcba7549ea79e2752d4351b63dc7663d4c8fca158af57408f3f387dd303b34b26b5855bcbfc27f2470741a3953d52059963f3b0a4deff1fb94cc1eafe8ef96e7ddb56c3a5a2e482f30a76890c723c4cba835d01749427c99366d00011af01eb098a780b0e60b247817e3f4c15dbf17094bedb54d694ca9875dfdce8d326c814f6e5d02847d0212c4f4e8211200a8ad2548c474fe56be80dc5a9baa41ecb795ce01107a8cbe7f324eb10bfc6ce9e5d9a77be794605834b7e26c6239dbf9b3a0a0e74a2d1bd1dbfd8fbc910411d9693221239b61c663d3fdfa0b08e3c13ba67b80d65a21716ee7573555b388782d784306d8b1c6f10409114f4c5dda2929d6324a5950555565476e11743ec7cb3918760ebc90ab792a29e18ce1d4a248885200e7d0e1d04b3522f8be168e5dcc4588e72a9418974ca3dd89a8cf56b956d263bf711d4115599f708a342f764ca2458b7ff12c5f94a8d5dfe2dec51c236c7d2c5d9ff16a72087b0186058f68518543d01da91bdb073e54d7ccea6349a5eb5a7351cf1274aff63002bb37b583e9428764000a5bd1f53c828a154020d1e2a5c076adba243002fed20288c5509ca7de498cf2cecc8e888f4aab418370ddffde9f6d76489884339458bf07b2685ed32e0689219255356de2747c6dd27325dddd3dadc35759f522a47db1674ae8d6664cede31e91b6f3bb0c60d3fc198cfdf944a60eaef657a66be5ddf341eafdcef61f1e9ba7680a11886524a0546f6bd15195c590e5c40ce7994182c83fa9702234f9b32b17508b4380284a0a4daf1b9ffac130ab6f2b00659a77d3fd9864224c0e0f6a1211e2f8809fd108b698789410cfc21f1b4542cb22c94745b3790fd6e4851e7b717327b2250879db5a3c0e888d79aa95872e129450e49effacac5654c0e161d795c59b2be96e2a5c3b25387e8e30b8cd1a1b8c4a4d447dfbc024a23e32ff4f131a18f5379ab543b2c401885d7e89c77762e6f07dfa8550a12d0b509315c2cc7a6680c6bd24f3b4ca7d5f0f0c44bd8b79ffc7651d58cbf36df6962e7241aa856f60d6b805d45c8ea2e9d8d71e9f08bcf0085ad8f31e50da26b5c1aba525776d0304148fea4bcf9b8b7acb5f4fca5b282ca31a597e8979a05ddffe8f1cce4648fb6c1f28e830f021386acce4838f9ed386b6422c3f22dfcea0bf3145ff00ddc328df6ebb322c2aa9e57d772e39228592bbdfe60e54e612003ad0488b83612f9c73261cb0c1d0081cd564cbc6cbe0dda3f56f272d2fc1d159ff534c622b2d5ec5f2234170194d00feefb781b002eb7acee0d762b6a326c2775739d7e7985ff930b710f0a70ca175fd6c07d748f3d5c02ac6fbd236b52d5cd96697f9588847dc8e1c855c153bb4dc75c0330e325b2500afb0f59b9d8eeda86c4d1cb782ac90e136eed6b84c6d5b5a2d8967257404960d769069d15fa49b09d0cc3982b7919cd859c2d7fe09f9881a15f544bed49a8eeddf133894050ccb0c48437f2cfbead3e2dcecc783937f5cd87854ff00a71c0d3b7e3bbebe71aeee911cf91f46f432643cbca28d646ca08fab115b4df2f16109b4defc6a1184200830be31dee5ce27c6cc5f5777b76ac7d675a2af8e662f90fd21af0f21a2508ae667656545942cc0dadb0c2f2490ed5993cae9974b456e11128f8685e0cfb87bc14a37fa1402346b65877c1a2c9188648ffb2738d918f15535be2ce9d3a0299a85ad8e37446f5915328d8caaecf23d7e8273030904b45c04bdf39660c9d67af749c9073907b2d98216383fade32267f52b2e63ae84d895a4527820d7f85d325a0ed847807f8824904818c36b157182cbd61a0247d33ed8c7f9c272a86353a1c8d33b300d7f3cabe952126f3ff2dc0ed7c560f77e696c67d3f082d6d4af5943cdd0fd82ea39282fb1a322821d364c915aae282e32d1401c4122ee44314d75245b426bee547d28b0f55cabb59029b6e48b262dd7c3ed3bc2500891e48392e9116e58aaec86e042e66d388daa755f49c1614f741ea93eb1e7679da2a761c8a4ec00dfd287c064a7dd660b303e9422682003406007db7e268cf623f3b72538126d03942f7cb6e3b55c61bdc2a67e0f5985b16455b2d1c503fdb6bc636a6fe87a749c02f4b7954ab45b96c7938bd18f50dd5ac3e593ec04d62faf9a3f9a57c5704b707eaa1ea7b2881533913c763fbb4f230983a1cdb09dcdd76389c00feabf1b86e272ed631df27b7cb729ca63c6342772ec2afb4b541dbaf7c97aefd525b45030a35ffec569ab1ee4033fc4e561aac6685f60e66bad3f4744514fd288f1e857fcf774ee2a439b5999fc2213a80154f49e031d8aa8b6f19b8f837c3feca5fcdf8d4440593e58aafeea022e0bab953a7b3f1083594d008ae627520af4350bbbfbf0e2ab2fd3866fd911dad02c0388ce5f595e5e30ce33553276b65235cac28194b032bc8453e08ddf524c67827ea4699b63725a4bf45527a430fd00e77323cd147d1dd33088d29601ed7366d0a17faa55cf6dbf1a208fb1728bf31050da2653a5c47c3c99676f6039d8c1905d28e6458e301bfa665e61c74aa5653d2d69ca5fae3936e3691e7cfcc20c4ca249f1a5e23a3e38cbe4cd10595c17fa6d41d352d4eb9b46a3bab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h433df362c9af02742ce23d374cd023430dfb6cd2da1bbf9f8da7b3964254cc4b2938e15ab5818bb6b86386761027d1c5ff5d817a4654978eebe3c03a9df732236178e70dd7fa0f57a99b6ed1eca43555deaf4c48732018b7dbc7bfc334acc9f482310fb943fa05ebf39e193c63155a0eaca185b8ab9af5bfd7b2750bcfee052f9c3f42bfcf77530d6d2ec3f9bb24f8d9eb5d7806e4c7047bd7fe9b40aee2f40f977003b32d5b4a40b681d05805d3e722954928b6d41347b1b6bd2062b480ada01f683992de9c22b9804c304e5b73f0bf350dce3596db31b1971192891fc2290af7bfb403584e33e9f14cfa0825873c9c28873a085b986c79d92a0848566a74bdf01e0a4e17fbbbb8b0c260ae9358c75794f1226924a3fd62693ba2b0451d7697d721f1b76f8cbe1f7e71f62a217acfc577b082e25d81f480bf4b3d6bcc9ee9c56f6e29ea8068cb935cd7ef2157e87060413c4d46198b43f8506e1058b053c941c29e8743beab8327e5b33386408674f264c9e627161b4da2fd4cd0a65cc9d65c6cb5d6ba988df07655890919cfd79c50816c466c9e3684b9f3d885dc00839f092f0ef69f74e4d9a1458327aee3826afd5ea128fa37017bf2dc7ea8c4a3bff174c95c67a290647de0000ea49fc7e1a5a6f4dc3d15c052528495d564c50ffe8316f89889509b4444964d36afbce65a321a19ad03daa4bb92de9af83766054dc6814f739cb3a724c97a60716acccd259e2c91cd5a1d9f03f078d434d1e36f866c87b3d076b0426235761f22f1aa345b9d6d8ffa2fecd987c50c0a3bbc9022bde4c73842171cefd098774b9b2c29e533cac80d7aaf85b7281007a08c4b72781ef18a2ae7c3b8ca5d226486f36e77e88b26cd56caab54128c0d4e3da8632c0a1ae3e60ed333ea7978b78e8918901c848fef12951aa147896cb51719c9956199b854992e98d822361e26f51cb7e7c6697bd9a0559da230f9335afa0f409f9899aa5d154912f1a3f9d537b5a7cd63444470758eae94b41f9737227a13eb0d8109b297c87cd22a40a0c5451bd0baa0b0e77c63f77ee7429fa9a383bee614f293d1755afb8c90a21e0bfe7c4466b25bb67fa69e227754658af3d9fd18ea09ad7fe1bf83d390ee32572164314fddeac043e8d745973bd5d9f5e8eff3cd6115c85124ce266427818be15ca44eaaa8b04352c14e09963ae231f86f3b9556071c4a01bae2c5983906f79b85987a669e584f37bd38192a04ebff62b31ab00df3a38839a509a9462d0d61120325f56ac66cff3057e65462f870e00a59dddfd75205e70e401f7df0420734778e9cce3154fd0fc5b10dafc47761df7481a16dddc3b27f3823c427bfd470614fdb48aa6518e51f7997bfda58f3a8999ed3e5d5183b9b2c3e238f29f7bd8023f3fc4d4603d1575f1b0a251c0add0734dbfd1ca3c4d07a3034e25da449743e99576f1d2ba05ae8f3c6ae7f8f5d6dd5bf4cb5154c419a8fdf41b5207d79e7541353450eedb710efe2a9f5977be08bc1b10d1b5dc8a57abc4285ae309e491c82f6408e74a119b9343ac60f1d81f5d5c4c49bdf1d28cdbe9888b550ca1eb5b56943e789c278fbf3b399600ed1c7cd1564b13ee840d12558a0fdf5364c5c77be49e211c996af6bee12a3e5795e04980670bbb15a1923fd700861bb8a1f64546da8702689a6dbacee36f23a934d34b8acad563ec37fc523be58cc797d64d07c05d8ff06fd66b54d2d2470a1731a48c463b69d58beb492df81260fb66264e196f2ffa9cfabaab78725366aa066e78a53bacb884f96a0cddc8589b9fec43f8c250379e7959ca23bac00c6fd248aa37f9d8dc5c2a3a365f5236f04603735765a3416338de04b4c9c0ec00711d2a5c1126efa2b84c3f79a8db150eaffb2fa246c1b5906d83a922fd81c6cc9ed31b599857fe160e87f53215437c86bb70c15b9952b04613bd5e61a9b4048962172aeba5c60c26b2cb3f468b5b2415a738ea406e84f38688f9e855e445ce4f67101ffec5efdb70167d3cd58c7cf3fc9f70e49cf47d64f57a63c016df483708eb2797fd393acc9f6c4d7307b0dc7c3efce5a188fbf3864f8956a369f490a859dae89161dc9182198e485990f6c7d2436f20f8db3f2afedc60c47fe512d8a7b8bc6b6152980cccdddbe5651c3cca2285d71df396e9e2ad35e3b39b6b7ae9511cebb192cc51ab675e4c863d2bf0768fd4b7ee9d0c006161bd35739764e69f6d6deeebdac496434a95ab70e12a7235aa061f8358aa0978168846472bec315f59579c422247d1114d643425492b984a998b6ca2b6eb9e89cb062df4875038fe9d730ca453d8bfad399ad1b7a0f658880a5695d3a818b493c247586f910073252c28ce7f5f45e302e9cdc35a1a8bdbb89d889a82179b339f8ddb4dc2fd966c25fc6574d8134b78a8382e2c8e1001b14c9f563b5d19090d6f684072f792a234b937880fb3386ea5e0d45d4f15e1fa9571674e7206866619355fdb940dfc4aef78b093cf253294c4c38f2a7c1a893df00ab247923d313f039ec440aed5069fb531fe5c9e3ffe3d43c794b1aa51c888b828407603a9097ccaba7e4db266533ab5e0c6f8800e487ea3cf0b94eeae688120be445f98721b0922d8f903c5a3b321ccdefa6bba4f4c70b22bda49c7865a4eae51e3e17a60b926a84c0de475f6b7ce558fdef92e9aecf357c6a45a514f0be584a063a9c6416cd12f841fa2f59bd7618d491afffa0ca10f9197109e475b2dce7745ff7f47a598022a824b7a2849326c9742040ce074efe7c4a340e0d47b67b9531b8533ed96f38a68563f5b7bf8ce691e88a6a866981ae3144490564df375ade077f2d9c4ca11b28335471297b863dfda9e421ecf27ab65fcdc74fced43ab97583cd1c3bb0220bb5bcf6579ccb46f124f0eced54ab831f899f0286333e09fe4ac83ec8394ba42a8a95a304bb39c45cda59f1e9ccf7b23134cd7ab5bedee2b5c1cc75752c18a2ec894712f60b3d73d99f16050f564b389c5842c77abb5bdf8c2d694ff2c59cb6d4acc66f8c0e82e67c2d37f45f8d31dcd5e5c4e268ad68f73d366a0617d2554074e2ff144df6588185055831bf24442a543c2a0f07df960054caccd2edf035f70f3d44f38ca127df3af00cbcf5db32cdc559c384815ffe4fe4add22579108d772b723c5b7c1659b2b105ddfe2df59784686aac7353940f3633eeb09cf44c7104cb49cd9a00f40b6705725056afcc34eba6800ec736f7c9341c364c24874098ef5dfe472deb7f0154d95aec6dc8e7c42a0ebdadb04c78564383bc0fcac3bb068fb7a3f16c19ddafc4ab8bfe905f69d27f00d15d504c50b73afe1424e760a5d0635e615a95afad880c8723b4d239ef3f161a61b10a9ce49f69598367a4bd94bc9ab3016ad18cc2fa50232031c661bd21ba8d37ba65b68cb29094ebf5cada5f8a72d42905b9b189d2c3fbc469493b196af44f1abf714c236d2388080a72c4d4e2c0517658ac19a6eec7c780db8ec7cdca286850c141d35968ff1ec2d6bee5bde69d88e82f7dda84938265a1f7173a77c055fff3d27b90d717e7286829f69d778305609a20289aa9d65ab77dcf54161b98895b9655224a3f87357f792b2c536494e4f61ca56b7722f26e68b7408e24a3c94d24a4c4d0e09938d13601bcf05b46e0d070f07e6ca60835b87206763ab77e801e218adddd9b4058cad1d8dd653eeac8fc71d91fa757e1f428dad475d3dbb5111b556869be5dd381d95cd2c289ac72b95ef918eebf6ed55e7aa349f6f24ccd6efa169a5df300d9eebfd1df6af4035f99e446bb606151289485add35cfad1fc8e8fb328c730c3b04ca84e2b480c3ab4197d74296f03b69b5e89680299eca5120439dc51b499bb9fa1f8790a61690b8d0947d1492d5c55323d8eb558768fa1b35539732f6ef6f8293135e626f2c7077ebd17a7d2d1d1bedac7575851668d085983d3d7ce7dac0005920a1fc42786db00c5ffd187001ee1a86d2efe93ac423687085d17b505f9793d6eb80c97a053fe14f3d892c2d598d0e010d5baa83b8a812261e486f7acfa7ce9e9e9b2810b7d443c11f10dc9ca25ae15048a4c1818109398ad72977e5770117b7bdf75f6b3adb8eda3d4f49d31a27358796278fc0b0e0854e92b81b402cf3e443f196ee79d3b632d1ffc6311fa23a2f8d23c9c097efa3a13a41cbb9b170d5522fdfff2c1b37fb37bbbb752eee5d5a031bcd688f3528c0f32f2570f8ec321d7c6b90eb4c3dc88c29f8f640350f40a17a478b2b367197b491669697dbab9d930d329a7e299e0d2cc0600513a38c3924e1a0c25d25da3eaf1aa79d5daac94b3109b0a4f6b9da6a583b11ec88437123ec3883709cd87229507c1d8e5a7e332e42d3aa6b14cfbb9a738e031953e175e91c8b0e8bb3d1bc050c68957f6338e49d616a489a7976cba0ccfd736d138a21595afb3126471b7366fd831502461a1ed0af8cd0a18c913fd9dea1a285faa384aee6eafd7e2062b9fa6858e27f5b713d92c21c71dba8c71de248dea97782743e7318c211718c609d4e83109057521959975803990e6851206ed861face01f03bf68cbfb2a8ce6443f359e5302340ac5eb6b10c1304bdf2b8d4101243a8b3594d56db35dadbf47f5469b24a2cf819b00d943ed310e027c3668e0d400236cbd7084ca0f3a1861704f23e6b27c53e97b468574936092fb616cfa5adfd42b6f39320d3dbf7b8da5d48ebf0d439fc9ce13b056c85b566dbdc20fc25dc0ef476456406bc7d839321467ac381f606b4151da30781ab1adfd403a52c5fb000bfd18e372f57bd853c2f2ba8372a920f814bc244c90b4a9928eacfa0865631ff7a33bfc4d0dc9c6babac93ce2803d356676f3b9e6e06ff1bf937658b93b41dec09abf07d7e7ae3d78958a0a78085a0509a40651e1362d33404ef89f8444ea8b45e54fca46cced901b9d071feefb64652f780850d92c3723c08783f4e4df438ce1ecf787ce43dc6c553c422c66ee1b4332b60b0e9cb2a9cd09dbb906a2794106ad7603477cc780318c7de4ef4b917e164d0afff11ccc1c75541c6ef1671f7e898f0fa6808c357f9bbd4604eda108c7baeb5d4480b698ca25d349cc204d0b122ffb5bc387c4d425c76372705ecc9f8f42ac973e97c40117a17013712b66bc2d526957ca1993358f91bdd058143c5294d89f69c3bcd7857e53831fc4b4cafbd71ba0c8d7911988b54a3d4e14b57ef5156e41788cf36f1683f3dc27cbc80ef5091ad0f8064c9f3556af959d343c85f545798b8751849b3cc534845d20fb55b8c783b466942e946a795becb18a0b921680fe23a138d19da5d7e22abf835d88059ec3f51d72e2f2b11653aa833512f3b5426b78bc8fe96726ae5ec325b9e14d33a665e809e9df30b2a9a2a6413006978c1956bc94d4953a34d9cfcf0f0656ca20ed88c8d6efc8dc9a007d0260f36f216f08bfdd5edb823a165c6640aedc680a931c849c1eb61b5824bc209ec4a1b422a5f53727511fd40addecbb0868822e9d69537bfa11689e5b5980db436671c79c2fc7dc8df1f281fc2c6bfe22e5c3067ba1b5223d59b45ec0c6be90d7b5d5fb2b9d8103a7d8c1aa8335f95af21bfe977d42b272938d72a58867cade51f66b1466a867653ac78e8cd346dc03913643db29f2c9901b2c3053d1e1f3ffe1f4836d2d621e71b6f787635c02cad289797a0b546a3452a9f432d285e209aa6a88a8d7f53aead078b9d96fcdc8391b6b6124981269be96fa0e466fc31edcfa216e050677dd82e116b8d4945ea40a9acebb014ff40e6ac306e70d3425faa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf07c13637fac349f1e823eaf888321c8f6bfe8259e8467a2bda2a5d2cd4f53ffb8da1f278985491ea32cc82b1552f9d0265e450349e14934e8c07a89d5d11d86947421743265a683fbba6b1480eb855f6d0c7b7329a6c758a621d0dc3aaee3052009ca443898a99463d045136c926a7b28083c182c279788b2e6512645d52794496c6119dca1b135caf9bb4fca65d6e232b0a0ad7c0be6c414aba912857b413facc6fe6af4fd166af030b6914bcdf43a1bde594d3f67df4575431aab5130b906715ee419b39a54a8ddd3ed200ac5d0cf99bfd52b2ed3f8074cd67a9535fa1d0c1c1651ac505e7a91e59b8e5df682cc7f87637ef3974e068ebaa9f4fa3111f8dca7f50e0ed974e3b89e0f55a82337c2e3d0ed0f61e974f78d0b9185e7b6de2c9a9122fbd9b51381a2ad34ffe4a5a77610ccddb5f4615360c171ea72fbc8a1660ab87d05077714437de2782bb5a5471778456e8d6d816c51135d33eb7bbefc96492bc5f1b1a61ab2834fc8754ad7dd482c435a29870a89a01519d9682c9f5549d044b38a27b56341311384f7cffb4c7e8bfd635fbe4a8942e5339eb083512f722511225b7677472a7052d2cabe6d26ac4f841e462ad606120159051da8fba515878f5eb59dfd1a800f0129fa1f40e730346fde85dc100dc0d0ce8896124e5809683d8645dfd2a0b99c797891be7757f74ce8fb9d27a7d7dbf4d8a01446daca0ca47d8f8b79127fdbfdb97fdb08d51eb73c2bcab33563bb25f78ede5b835b126958c76c5ead14bc8f0e31d962694b66683ffb219c16676954183f3ac09ad41839d25811ceb800f7d156a5045fe6d2085c20f31edd7f1e2d09659eb07925fa9de2a6d30aa08ca1c55f2125d5038a81ef72da1738f4942945fd72489ae340fa0966a08c0ba088e962ca29ef109dc84285081285dc718a1f5c0fb7cf074995549ad27b51073516b68254f5539871433894b06fd5d9d99a80039f6800fccb2c7ebeb3ed2b5cefb599ccbd46067658c6837df19138fdb82f3acf4d163813fabcd9ee202ec4dff23a43ea3da3687c1a4b2c6db36017cfd134e7929d1618d0085231ac75b15d048031f2714718976218a619e4651ae4ccb6104228afd49ef8d6891dac3005cf4d692cd202cc7c31a3a4c26f025ff2761ca98a656feb01985dd8f84974a3a0ce8b95d59dddd68af742575ae7169d504c476ef78236338b8c341bb10c1023d31d321a7de4946cfef062f98c2f012cdfbd5bfd2fd05e3ca11f6c930c81a4eb1eaff5d223abf62581aa91e1b2d120d2a9ea2c246dd6150d1394aa9e43bbca009ea531bfb5f727b38394992aa4363d1000f24e23b4ae7761dbf5422f7e3171b073b73aad7817a1904bed86d9ca42f4dccd9947b8baadde8a6bd723382b2a1086ed02266e021ff1cd5d56ed40d0488b3e7ccca8b0572828915566fca57f0df180686bdc0731e4558f1e145a53347fc1e670150eb46faabd06c7602316f034373e64d272da8680bb0da8a35044a75f3658cbad31f9a07820df9a2f5d0ee9e4ac03f3f791c7adda821bb003fa36ef6f4fcb37126fdadcb84fc8f14ba57f9486c2f1c9f89d3b016e2a28e2fb23a5bf91182c1be205e2dd8fbdad05f6c02575405f6f8b9d097e103e092cbf8e20eab2cd59c3d2c689c4aebea6b36bbdc308c527df5d719599f752bcbb1b2a0bc0dbf1713ad76d16933bf954ed3e509fda9cd534dd8426454db42c739ad9ae2e1088e408b96bd8f33cd34d2b18f5f87e2799bcbe4478ac4d7d999a8508ae9659d676df3fc15a26400f89acf4ee2ec293e0b01aa14e75f91a85e159cc9d7a423a3c8988719741c64ff9b3536e17dce3e2a16fed505491ffa1be899556ead42aa29c003592a0c6616d24704d84ff74f025a3952fe301f62571d351b8b4ac42f985f30fd9baf958eb8062580e0e14c6d5fa8ed2ddd7dd1870f8fb1af240e454338ec23e65c91821c830f202308177050b5bcaefe252518e6f1fb1e1864d43a0f92a7211ff8b10dacb947a7d829a580553d38b29875c564c188ea8ff025a5148190c70300663ffb5704de9924a9d02f1e3ee421dc5aa33d3b1dca5a387dbf5d364c5bf125bd156c78a018b77088f50a4e9a71c9d7300b23a902669814d4b01dce0c8951f9bd186e357c7f3b462caed4b4d195cf6f906fa1024141572656e82fbe1ce2931f9fc3cae8f5fadd63f612a24c92808608c8d31920f90c8101262809bfc47441a912b3209a07da2b01d38fa749ec75005dd29db8960d9a4c0a910d5da1d7cd9b3111d71ee41d1c463b4baebc692f31c9cad27dfa2ab89f2d8df538aa231a9eb24451b31089a75cf9259250b151dfb3f1c2c3d89549ff517e07b1298f57143d69aa54fafe327a4130950aed9c753e681100e2cd87fa2249c3c20b561bdb078d28424da67b42c0ae20752da4c31756a6b94d51144ff36de868fe526b935a903ffbd276f2740e2448ed01d5b91f375f4b547be5f45361d83cdc5599fdd69e1ff54873185c8e1c55930d4248eb98587373c6a05cd02e4dbc37e104acc521a7330792a6f7b76ccf72313e035a57863cbd586298a2455f5db7882dd665260a4f973c5cae4c14ec86ad33e2453b46759a4dfefe228616020e946359b1eabe10462c2a90405175f257d2c67e14aaece814b33325ffacad09fb1918e71c03ccdeb8a08da4e540b83d319c3a97c60f0f02c6ea65e241f9b74fe20e8591755e0f24f71685f8d804c1153283636ee68b4c0941b500d1f337f8a75efb44f8d5548e08adf2bde807eb86bf66987586e9975912918ae44aae32f679d6b8c8029ddf07817340b47ab15f20c8f41c7442c9d0a62bff48eaffb186152dbc71c7c4cd5394389a263603896eef6105c205bc4d763d24808df0153b86e68c244b735f9712df0549437f05dbd61fa68fc8316e740c5f00f7cc54e592cd06b7e9482d03f3ce2ca04e3d8dc5419bc03b6f8bbdd5a32677f08fefa7a4957d3f12285bd6f99802d98a6fbb8ad2ceb19847fbbb82b242e1a8c37b17b8b08a035e72aaaf13b2dbd9709f432c928a890ecfc80d1006c4135c89656e536b77b71b66338e6d44dcbe212680c9959b407e447283bbb41ec236e0e038e93418bc8455f5285b68dce62a91d87bd4095791c83fccb750c765dffee593973635a89cb82b90f882d950ce714dca410eaf091e7bfacc49d16fa3aa4e2399c9f043057a6f7fb1abd6814b4b85bc946170c0d6569a0e30e428124fe5e46792c5dbc9cd5f3e16924a6ad5db067848e115d12e78b70708252929cf501a2b8d45239967c1cfe76d601d704ab4892642c3a2773b06175024b26b57de78c29b70a3fefff16d04b307b59a7d09eb7e3007c7b24cb331341a0486a33082cbe436a441811ec157ef5c410ecb64e6ac5cf9b67aa5b5963668f739d5f43cf50cde0e15a7cf564f1e7457661e961224b1c54d2b094b19c4121389e6042df3bf07121c1717d73e4352a93cadc193398fea3a3685634bc018b863dd42060bd8507f6ff0b72214ca13a28c9f660659223fa66c7bd9c455eb1a7143a55e0d92d7ba9c61e17d2a9ae59b296d8787db4dc514e49c0b0d432a1d22d0b7c161256bd710ba94f9fec2ee82c19842841636a727ae617427451187c9968b3c9a14c6671b8966fd8efe1502ebe47c042695f2dd37a43da12e9f7b9081f1507857fd33e37416765d857c02737a0075be0c28d59f4d2664da563e4316b3e5588a0f6b4f018ff2ffafc464b6faba7ea4030b4193deb7421c2a1115d5969dae2d38cdb7f35d49b394c0a78532c2a9cfa0bd334f2eba4fd2e13ce96105ecf7bff67c25ed146cbaab069d0301f131947fa33a907e8af14511c6ad73ce44b7822055caa700b3d1333ec604487f7bd263588e398ee8a9f7f499a060e534cfba7ec9eb4848888fb46140029bc50151083594a718ac433c1f487547868fa2f9536e07a76ef3a3d06c2e531c03eb72aba772fff92b0f20c210f4693d81f91dec21d89224a03b911db19600fdffdedaac4ae77fa19d4bfeb7ff5f322c3c4f7821f6816cb703abdeb75ebb9c57513d0ed22ceb76406aa160e11265513963eff6af9593de4128e3efda09e636964a3b1b89c25cf2a7e6fe61aa30ec723e5f3212fdb5dfd78fa893d2fb4f36e6631e607110f14a7d1d117f1a7e172c633dc3adbedcec4f8b01547e32bdca6bc1ee43f94d3402eb76819dcc2d33cb62e4c5e4ef5329a88584ce63daa223291c90746c20739f20d60abc0991a04da489dc251c5e9385931329d86604ea20727945197e6868eb657df41756842c2bbcc5cd19dd0d784dbe84edbdebc103741ba84ef228203c2854fa9e82a854b7acbc8e6ee4df610a9d753c0596fbc77f5098b4a1eb6d14d18486d53fd58843b0ba39f0b33a440660c6b0f1b5b7eba53e1e539f9b1d48c61bd15cd99be6729a9d4d77832d02e7641a1fb1660a04116f85fe56e85070c39c2c063ca0865827b4998d4d9c284e2ceea8a409d1b3cecbb2f35d94b915ae54efafa3fcceaebe9b82306c0e24efc0556608dc9b21553a2d6a0a8fb3b347c196f8bbd1b23025ab32feaf6f01f98a8e99ddc4283c0a558e9bb0a57873195fe2604908ad28fc5bfdb42e26c2e6cf2fac45990e35ee37357b1aae4092ca5b7af1285e4f72bc667e9707932951bdf5306e7e914f6f72ba4cd1f5ebd4beae6affb7bd370318561b1fa75e4c4d3d6f55ea0540a93372d887c39e6d3e7991eb492d03812c4f51f19819f0ba42546444b8ecc784c6bf44ac36897eaf5502203825741158010d6ee9d49e9cde27f4ec1d7ca3623cb923f110f43ba73d009bf68a0188e4f0433016f7dd9c9145825a93d54dc9c92ab9b1af528d05fa9df5241cdaecd52f2a78442c5ba4b8ba1b3694d40287b2f0f67b1e9f51ac85a8b6aafd1a7daa6e9bc8b83de14dca384fc49bba19a4791513bb39981a2131ab16fde65ffa808ea138b705b24c1972a7cca3534b7c07c24fcdc7e6aad2a1f4ba3b97d8e872e559a10af36f6a91d9df86af3897ca5daac25043a8d1d79fb46f2cc16bc7f835191fa242817c7b7c902c96edb258e2bf492eb2d07506b5f0a9b2ba6f589009799addc45a800a846c4ac3d12a7574608301c82290bdc1037caf276fbc6473ade3fd198ee42ddbddca810f14c4176383c71efaf15077431069bd553a2b162db5af3eb39ffa3737c6952cd1d2799af24bf2870d3284cca915a2fa6cbebfba9ab8eb45364afe6c38a1d8e909e1c71413f8647b9db3acc9b78f6fc48483a4041f860d03a853b58f95f642f9413c51fc908995b8c134174143b8bca40261f7528da6eaa301bee3fe99fb79575a616623ede32839eb207c28510413e14e684dac92d19b828f0a61cff6d7e39a5c7f0fdf7d059cb017bec2576c87580bd1eaf4d5e930cea90fdf0af8b1bab2fdd421c6a57e68236df48e007697daa0ef49d066ce867a2cd67c30895b37a20a45a7c14dd92d84da024f59be6f39e7cda81f3a5769e7bcf36dd0e6d940a1943e19df491296b190190ca211e208e2ae49477e7dfa11c86996c297837f3c89b6ce902191e1bf3bb19d78b5e7a62daab1c72b25aa4e1642e78b53fd3b1740241f16687d8e2e9890874b7ced40158e07c4f208ef508f72727ce05223e9f0f73fedccb583ceccf739e9fd734ea46ea96df6a07470b2d3bee3c93b47cf3bf143303b6c1070c129a3ebf1601ae16e88f599a36d01e249878389f2263c80c5546f5457b9cf9f02d0925ae4bcd2889198657b4b9a112a98061b838d774b4c2698efef99fa2953be98d99eed557fbce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7eba33f72da66e4ce72e2171becf06d5ca57a110b5fa459981319d4066de3d2499730a3243f0b4b73d9b68377f475d2abce1872a77f32d3f0951391ad051437d2415038360b92e10156736ed2c5da97a96e12d93ec53674dc1abf87dbc0494e8fbfd7561e70f41fb27cacd08362420e62714d6040437fca5b6a09af68cc14f563ffaccbcadfadfc64f4e3b684bc27089178e760abd377669d3a24d45b89df19fd249099519a420c9243188c92d3d479804528e0d8656f63f8aee51c4db16606e0661f71f48484f9a6bbc8f1cac5470378fdfe6b9b9df94c588c586bc47f28741d3fe2fb360c244ae99cdafb88a9ab8eed8a3732002453157cf7e36b4927a9cdbffb9cfadf609faf6d42e8882a685be034068a7b81e2dc2c894f1d7a2293073acf9f21e8596985c625fb0eb1f6ee35e1e010d47ed8f0b59001fd94a8299aaba17c56207c895507f89f86c04941d8baeab4260b383d4ae9f126418c1596733e2084fcd9b2546556b449eb0afb1c8a62a08e11775af33f213971e574ffc07cf0814f9f0927ef3895137e9a64b24b6a6b1254a4c4a9be9260592258366a446af1650a4ae548c20081c748adea50168a84957217e996af30265a6067f1893db484a903adb3e1a2a81220132e06264ee3eaa371de216f9f29b3b4392cf6bf9aa9cef054850bc9c870ada67e0661506d51cdbf50ec6874d8bc2d98525720c14c1b9239f6af4282e58347bde464bf6b518c3eaa67b35c6359f0c924fad9905d3ad770d61112fb806b382864f0757a732f37d3fad4c38f6fdf55fa692b365d86c2ecc1ada59d3a2b846f25d7f0f039248b71eb0e1373fa729e097efe8c8fa97b642c9dde73dae36ca82fa8cb0d85c4e43f60f4bb53f09382841e510a5712da39ec87d7466fa0e2d0faabf8f212fb8cfc1e996409f28165f911512b702c39c0ab3e931a8eaf5f0d5de8338a1b13f7b3821239e41a8a74f728c498db49c53162ed0767bfedddf95ae2bb16623f1d236aa750e0f2bb25b1d53b5da14da50d32e47bb51bd185f4f9681c36a8ea880abe73da44fd9db74017b3be9b2cdbfd8432222ffae8943e2eee455c9e78e956e8896e0efa2d87d108b50ded3420c659308a935991c41fb452dd916cf379e11fd47054e630e3177f61106dbb1aa64e62a4ebb6706e3658b432ecb2709dd15b9d45c51aa3883761e82568457f11aa99f5ea9da897b460cebd803dbd90c5aabec5b481859381d399a871290820383230605bc7d48a9f9b2a01790fa0fd54a34292232887c2ae71fb7145fab6aba09d1fd5f44cb6410897425a20fa85223a097925b7098b6f4caf4657261981b01828f96ad904ab9f1e6976e72dabd679cc96ce9d7ea2f30744f53edc7649a30ddf540c02889290d5bb58749da7d3f26357777900f0ecebcb9756834c7d39b99cb24f64be5d4a10dee2fb5650a9de9c44d92bcad98cf40f1af67b0ed56bb13ceb6459eba4e22f8526b4057da27714f9357df10fad04e8550dc29483db69ba36f3de0143bb83350401f30132d2e4c439240a69b8e1a1ece788ec3f7fc728604b68b6ddfe1dcda0a0eb1ea8e4801da5efe4a5d1153d4791e178c275d38e310cfc5a7f7e48d4ff5a4208772e43cde764de53a53bb978f7d9716863bbb42406808f4995ce84658f05ac9db2e11d4334471eea607d0662943b6384c2ab333e67bd7adc19ce0107bd89f78f907db57682af27aeab3205a096486b2a8725f82487d836c97292cb443d571a41b0248a18d74ebb4cf534843afb3ca6c5c6ed797fb726970b2a13a61a0f297c06040ada38c88c6e2982668f50f2b253eebd7f4e585287864c0dbc9b43ecb455df2a25f37a4131b0ed419968a9b4971f924e3418bf55954a586e6dde756ec8679911251bd3ec952f0a857a7cadd26d04898b3ad8f9f8f7379ac02fb001725a4ab01e5dafc5ed2ba8fb403f60e8553a0acace1b51d7e529fc03aefae502ba7da18eb919bd6b3083edb611803265ed8d671593b00f5349784c1411cca16fa6bc152b943d08e5389dfb0cfcd64577d25496215f6e1cbe3ccfeb82fcdb0537999edea470fc83466aa37db108ced62fec0e9eb822dc9556c418bc4a7ba341e8cab2ddbb51045acdbc3007760b5002185cc42e2bb1becdd145bee25549a2c84644cf11a87ecb234652cb1125258aedb3813e66abb4eafc88c2e97a5a913722bb75e0185e350d285fbd3a678146ce77f8327a45d525a4b0cd1aedc269a227046f8d06b5328efb0ed5231c37d2f58b2ea7f899c772e055f41261134afc987c76b956e085ea28b8e51da60a1aced605dd1b206a07e65584fb7406ecf1db3f62fc90af6efddb248bdefe31b3bb6bb366f196dfb1ece394056abdf1999a147859ed22d0efd11e3b4ff25b59b911acadc156d7f381208e798936a944e77f3df6274003ce544d06ad2e1953b5b9145dc95a8ffd27a53911cc1477b5d90baca50ae43a9155bca7f514810875f1609e5b1a4e295afd80da17a3edb98ab2dd8e2a09ce206514bcf6144453a8b225c019a2dabd9f6c57abe49a0990e9241656ccd81c32e423ab2c00f696459d48bf22a94cdfd96e4d9f1957a762dfa09b8f7fc2c22ea974cc66383b8ab923a6f3fafef463109b06609902bb46ec25fd6fd5be73110cb970dc89f36aa93d0879d70423417f6a5f3a691d58a8d48657669c7fa17c78e503adc34b45142604b733358855712dcbb9e43ee02dfedfea396547eea58ca720fe956874e8fa05fc92ea66ecc0cb6d0ac36c1a854304a47578e03ab19a29b4123e46f43f13404fdd2c747e61e1e915c38f46f2530f65d0c7aff9f84d47a1a0dd1d7d8c84a2399c659bd534ccf03eb85731e7857c368337dc661448e472a817ec43e9fae299ba892497803f60f29e87656ff0ebec95f6fcc1d8e5258ecf6ff61baf8f988887725addfe2369da8d584f6b52d745961572bb55de679908f42b82692c6345b849773a57d1bb7ab9ae61a22f6705bfefc0975adf43beb489f634d0d6fa2cb2227a77b2e49283c9b512c010d3f8ad91d2c631851fd08f5a30963427a31c18c54799165d0091f81dfb655e62e2988f0d257b12cba2dc7587934ffd223c4245008ba4c0ae293696c374a79ba14cc710f8aa1b73755feb1ee3b76583ffe2cd2ea69a7b2f0db19015d2386e7533c2042bfbe45b6323ce4b6686f34d9b8e1118b780586034ad2b951f48d57b8124f4faedf8d43698de6c5d47d19c311a03b07859846d26c7c0e7dce062dcd53404367082a0a190edd1013d86f9f0c201947cd9af75dcadf44dced343f931ffa100e23170980a95fc581f08500f8bd93fef22e12e27b202ea673436dbd0d1594fbcca6d4c9a4a2c1ce8988016ce787912a5b4551f89558508219d064736f18967f8b33be7a4f292595444c635b519afd2604f8fdbaf99193bf2a6b1b1648b9718eee347d0e755c0d8985bc10a7b72afd57ee508da5746c010e1584aaacc66df358356008aa69521963c6dcc0c8678ddd72ee5cf078429e990fa95f75d848bfdaee9d7a4bc0316e0ce30b9eea16dc4b7d2911c6ad2e5ce619e404b4aefbe8c6a957730b0018ecef139d75aeaef6b31e5b5765e4593a13adca425e40ce8b0a9d9259ee0bf034f6c25631ff84f8681ee76e509d6b3cd045c6025bc7733f38da355a55ee236f269fd082367203214005a8816f0db267dad9c01c96a7c2eca7cadf6fb75c7e04e9372cefb1f13b1d26f088f5aefc812a13aa52b56ca65ac06076cf1d7fbf0fa01c0b13d61ccdac65c47f62d72c52e68ab0b64e25b137395072c5558b02660959e7f58a0c75a1b1dbab2f9dbc283047e22b50ee8f774f463a3d7e72a64fae8baea990b37b8113907405c385383b02bf264ace21a9c926165a765f300b574e3a67bcce6900351f9312656f26a366c85c229d1c296b0acbb0b74f58b3682a29c0067472e4a457d9991b57350e05e5ba4612576fac2cb4622c95903a7d6f049da3e04164666d8115a2102c0d0f96cc7d63e7243c9f3a5809283c9bbefe4708f1fcd7cf5217172c0d3d7a59562d8815f5a7e0db13e53003c665629b2d7f7c924859989377c9ce9dbf92ac11dd41c23263f455c1619c5bfd10e5c92676defa3a6626730b219e272e006ef051828b58ecf183b9941feefd4870ecb1c41d5944a2f32d82260b6554ae74e21edbc6f6f93fc1a887f95603b97a317b4512e7821246f496fd90935eb0e0604b12579660e1a49c7a7325a32f06bbfbe07b4951f2f3dd5a8d5ec61b655868fb35f7395104d27fddc02ab42853f6758a6439fcb07146642fd3894b06d26be087ded413e93aac829aed824212f76c9a6aa7572e713a065f1fedc37162bf5eaf676ee837e21ab3cf76bdbed767c15cf32a6f0cf64c204a75c213d8e9124504e75bb9847ca6a11dda9181d364ebf1d8d700eddd81a0450284445f52e2cee4c3f102945376a23483cb560afc55e252a30192ce70d44d58383fb9a64fa2b62ef5cd541a3b7c4c26d90677b2a881b46b121f4202ecebd6623a1bc5521c462da3fa635d53dcb3e0642ab92ad34710fa11969a9fdc42a07b5ac2bee5f31a40ecfb7507d8f6e0295dd4750a32ed995476db71bda0ae3f3a7a97c5f9bac887b2b31ee711df42b7f0b799648e252367f95834854a4dbaef663b6eebbb0a20d36621ad88b3727f8f73165b21225f13f42b4fa3ed21cc58feea511fa0adb7d83b034f65c72d1be2047e840c55d088c72a94feb874d659f721a0153c83e97d4456163a2670cc73b0de5e20f0658bd93f1e1a5f06fe80c50361568b1ab24ad40d90fe178b3211cbc5be7ae6c6fef767b2268827b29e477f97dd6b7b28257ece0d7ce82e87db4efe2a4649bc066615836687682ce248e766e36d8f69f0b3256718a1dc1edf2618530c65a84db5ac39ffb189959afb68f5eb5f75070e0278b02c836b9d28a3eacc281fbe542f38555e25e2f4d8239bcb8b2fadb7bc35e87a9ab8b3e263ef7c8fb03d129c3f09744eba660bed121bd747e6237a9f64beff5f45be72937539b00b01b9e3bacfea4fb438b3b41946b357c30dd588a6c97e435d2a896f23bc499d9b8af74eff1eed2831c6c363ee82bd8d8b23fa02d530a2afc4c02b51cc53354bddf5f6a673b165c363efdfee7c5d4180e940501356aee23bb55a84b70bc1e94cd69f090048467c5b78ab0ea2452aae5d9c7f5b6f5a89e2e68f6af5f71e86d0353610d9bfb322ccc600fe303e55857f0bc7e88016503a26cf657863e7fa0cf98d2e8068f7e7c627772f01d636be3a5e64652f34b2b6fa85c4dcc489ccee5bbd7b5068333e7e03ec41f8a6c7fbaac30006e96558db8330a200652d990c6369cc092e00cb3ed4f0d38442371d1a1ff3fe4ce9fbbe4532c45516fbca920c31d555ad338e7beb3c38bce40101c886b3d111350143b60660ff764ff9c62b9aebf4bee8a8eb75c46e7a5a298e0c735b89a36c5826b6213bab928733fe51e20e5f40c303733a425235cc0b577877f1a1747cf751afa6f54a2ff58555119375e7fc8fc3e9925949f4a8e4442e383f7f39f09464004970e396a6fb789fc9fe17f5fb800ef5ab4d3f7710924860b6fe46933db68661cf9229ff473ba4b7b6c398592be82aad064f741fba701a427dcb537bcaa8dcc3917f7913e911ba5f5716bbb6410dd89999e537104edbd00936dff75b7f316e75a175f6b82827835ee5753df1f47044465bbf7393ede0287bd387a35fd93c740d2dc5d46354b613bb65840deeef6e2219982a7f825f1de77c38e90342061131005e6e7bbd79753f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h60cc7dc36c099e687cef2fe2a675fdc2191a960604a63969f95a48f95122c38aba0138164ca7351da9464653b57f536527528646e0181bc2d37e4fc30905ce3af0c5d229bfafdbb8b1ebe277f31c9d0cb795835588d0b723b7fdb1dfab08aaf7d89c7748f4db20ac2ce6c5ccfaaef8340656f4e60e165605cac9aed03081e05afb2b043a2562ee5f10654bee0d1b59295301ec7089c55778d0984828ffeb5f4f24291fe5c8165972c91913505b1c9341372c091909597ed233dd59dd2f637ffbce231f7f154dec2ecbc04ba03189964ec6788e0bb0c74b5dfe6b44fbea78e5a3cddbafbab4f63f16951c6b38e7cc6c4ca69a4983b8f1960305c5f7a433fb946225af532471d499044e58903836cdd4f8f64677fc4a164d64b18618ca5e761515d7732f84fb7843a3b908564cec2a80ad839122b7abf16ce215e798a5ba913801e64cc7eb04e652058d8e89018da29db3232dcc2f61d4cc306d804d16f28e228dd99aefafe1a84374de771f0f8e7cd4e9d7ea008d75988089ee547899b77f65f4111afd17f9f3887a6c35eaba064b800ba4edf35e72e7a99d849fba72ca4babe7a1206b5b803d514b544f52c2622474e2f04cc02a58872444182c7a8b7820e9fe06b3d809b228a9d606a37b551ee7080957740956bbd14679ad3f2c330d52e2e56c545733e6388f82c277e9e86d1e569c6223661dc1ef5bb6e833498558b862c4881547fb81ec7fb3eb04969782c9d82fce7e4628367ed2d2a45d4ab99d52915bfb9d7ce64dd17603115a5edd037e7de44d4ef9a26a0a613b5f224ae22344750adb54bb498e3c2a960edffb018d74e32ae4b0492dca1596d6ac1941938b711f5fb4a0188a92981c3c9cee0d837bbbf7e4bb380e8b7bcb83fac3a2e7a14ed70816e32d84b715f7b1e708eb8cfa7b21d6bba902ad43ae96b540c79c99a87e8a1482666f81af543c29304de98b68d37686f8263d52810fa9dd9f5d90a41a88d99d9591261191b56ae57fcafd10634336ae8f8d28dd87da28c4b6d68b834dd0899e0716904cdcfcd282f50966a7027ca6e333829dc7e4a0df4e34c742095d8b0fc6293e00ea469c51301d18e2d4b73ed465d8412eb78df575a9e73026f976cec392bd7ae9c06b9eb76d0d850db5e793493398a13d9113452597f5cf7e57ad743820fab5417e3ad996fc5edf19b848a1859b8caa867f1a3088cd3a3eea48bab1fe02a9ac26813fb81d24cca850180f4979f99ae19c67c963f3ebcacacbc1da1ee1a8a3f796535e1ec569e66d47375c85b2fb33a25c97da48ecc3c606b19e02b417bf5d3925e4bec2335eca67d43568aaba06a5536f7a80dc2c94ead4f94e6bf797ac94603d35626ff8a1bc50555d48ea210b13c11112030ddc988b68c99050c07c2043ee2a26756ccf08738cd992112fe7ca5736a5ab1eade1e0bce717f8527cb95d779ec97cbbd2287663f3c2c6cd648fd04b5d06578728ba6a728a04443c1897f67e952cc6aabbc140e73e3bfa7e9b289eb42c5651d6442415014e868394fb2bdc5737436156e05d0691d4515316a00ebaa599802f78ba746a20e27af97f891209ee3e5b871497e92d4a067c2b3b48191a465a3ed16daf6061078a954b3c719c687ea4ebfdd6b4d0b26b540378f012048f661da832fd1b319d09a87b6d1dd1a7a051586faeb025eb0b80968741d83274590f47045ade19117c5a80850ef5c82c0d1cb2b1983264690ec34fed695d5fc765155366305055ffbbafdd738c661deb817156450c1b54ace349d9cd9e89adf915c225ba74821bb9c0aaa3082f1ed5fc139d850ea936851e707a0343bdb5b45f4f4555108b1bbc24203cbd41ccc439bccc1460b4f66bb34d2c02309f17524dbe5c7c99185d4c89a3553b65ccaadf68c2cfbabeeaec77586118c8745cb1d698c1fe4296eed186426953f7bdc71ea3e36fa6322957a18105b70859f87e47be2953572f8b4fc738ffeca020a58e515f0ec9e5f6bc604e949e080f87e005c907681487b3939663bc8120125a4650e4d0759f9d46510dbd20f89accc8452f148016fe9a50fa4c2e24d736616bcdf651e3e5a35df5a1fa58b387a97c3ef2a49e5183cf030cd7fd30689f7ade90d5e4210c24e8f0ad57302f30b1576d1566bf3122996d5b8010662db1c13767b4b64b68c793b7c2676431c7c62b61ab38c4f5f9421b4ea2030b08efac9f512873fa0026052ded925f1e64937f023f52f852e3566d0065bef5882dd832576ab9243f06032d19a47a69ec4d30e9047605df3fa319aa18c40a918f0273d45db6e0b71e1f5564f53b1fdcb495edd93656683684e472099494e7d7e686b670fa4f103661e9ed866ddd23a8a28063b35d642850e419e27702c460ccc621d3251dd2776c8169738da2835b9eb83966fe48ecc0f40494e9a5140de91cb4b2bc52353adb3ec8cb8e0309cd7e7c03fc65a24b481fe998b494da6cf16e2bdd94647a667b589e4518646697a704d7426d363f39c0d2be2b4e785d2fa77fd4ef1cae676978ecd81d85190fd2bc2e9b27db4d5472d1094eed9eb7b3ba474d374facc98c0836b52c67e22b4b7337f81a1224e5a3d9d266dfed55754f45ba4dc525a148e3817e6b32d16c17b87dd1d7484397bf41b836acf0e17f457f6987e5896927364209a37fa9299cb2aca77b8426bce7b07570f2127a80bdd21c17556f454ecee2a82d0dffeaa1782f4f67e78755eb7e01d1847dce1de22337a40bc0da2b8cefb39b32c59ff4acf4717cf9eadca34463fbbbe2474575a95ce61a1d5e88d69915a95acdf5387a11295a088f2c8b3e40b9ffc21956bc0c42b68765d620badb7e79c93f40d35e3d3bf8f443e523da9dff8f0a3b8c09e9bca99e3b30a486c2c1a5f103d1aca697067c43d1a0a0b657e363616b7c2c6d57b928bf4a2acdf20f9b1adb652eb126b4ad19ebbdb30e93b1cd20fbb8fd229b406d2073d7fc619f60c2d1d1f958b23aaf2b98d229fc9c92a510be275fee48f346752f664683d92c1e742a90e6d4f254c684f6414936b1ef70979ae426521c7c3e48615d28f7d870319dbf49699b16b0b175d54efcb9046bb71440304a4f8657c3dcf2380c39cbe90a63ac4d051dc99aa4869114b7696f1fbbbca1048dccfc8057be751e7c9bff782d7f52e056f85782698e5e98d06e3b648a1636a48bc22514c2bee1b2da2e9e68d32e1d4a5d607edc023c3fa7895477294b32eed7dfa5f50e4452b524fb10105c13ffeb493e32f451e690c13125e42e2986710864d1effee7c9d91dd2545740b142e12817b030841c2f4103e62a2103bb71410cfc8baf5a643dc01bf2571d52d08138e68107d339c66ea869c039e7e3bddb9e8e32f4efbd3755b32918e1df8b9bed53129f3479d47daeea6270343729a0d91a59237bb9d60cd212257c6b43a5f8d87106e51ecbf1eb8a2c760602dff86ac63b147576b2bf1fd28119050c901a57a2b875036cc061512e7d81a4609321449a0492e110cdbb13f4a304690d71807b6db0042643f5855eba73ddfaf5aad1a003a44618c6496380993ac148d63157560964c122c5b4eb0e621116b44b0034da610cd80e4d5cc7b4aeb98471a3509bbb1bba23355f0d76a4a606b9e706b426f8d62a63cec7494d1daa3716567b4638fb9be6a11eb205303172cc77906dc0ed777b5e7451c2cfedda8014908d41a169023d86a2363c9f2d09bd54d610da0ae9c22653568a7833d9b321297408b6a6bca2557fc8dbf7e625d9d757d392bc7ddbf77a5e12a0d7411c0057bd30f214db56527119e5917873496c6d82a4a4ac6b0dbfae4cdccc75ead1c0262b923ada95c5b8c1035ce441f66343cde046168025738dbd7acfeeb2fb30eca5faee730242b2043cf91535ecf808f338baddd9b5ae1efc6ffc8d7cc380560cced425c21e72901749afa4d9ada27789c3d21ab1d9dca2f31e3bc58e3fa7c38547d2a799f081a6a9703142b175ac8b8db768234e53d514a8e7803f53b2adf8f485d80a810bf0fab5b3606b4ea9df7c394fa7a504f7fa89231da2c195ac92401c7c390d602b1f9a1b73bf1626b43c26a3ff58ff439f4cba199b01948dcf035ee20b2e9c4f099b24fc23823853b94293a59360f9b93a6ed3682c5bb8147099c6bad2aab2b0b3b092be44c919f74d2d35fab95f6b2a1f253fd13cc895db45a7d503b5f2718161b7c2755659c1360c6d7d484bc2d2091423df82cc5ae4db9eebb98b6a2d0a960aea45e21248b0cef930196a39429cd4a7fe7d2fa7db90936794c61d4d0f2cea49882df57251743bb84106cf633367cbbe7a847a1350b0b9643ccca7e56001637d80d2c340e999f040157908e5bed4e04b6ddd36eb98572fe5454cb18b4e0077aa196fb39a410a2677453a6c0831469631b93a1667f63abe1e4a6616228656ecf5165dc5d16e7e513982ca3ef65ccc194cbea5cab0ab665939ecc6f7d0735841457ddbffca232c91ff31bedc8055f742df3a2e6c9eaa12758a914ed9f1fcec590f055d18535a5aa4d5a4cfa5e491cae263e82f0f6220a001a9621476ce0217f7fd3e064a013f805a85965eb7f935732b7f616d5786410a3f15bc82baaec0facccffe0099271eafda6157f048b39b67311ee974132d72646231430324357505f3ab9a90e4165b0174915b33f0f39c356297420ab6adb024a207062fc93dc8520cda661a803c152453af57ea802132b8dfb331f1c889889c0535499d3853c0c6e3f5a3c341bb4820041ceb731be1db8bdfa1545b8921f4786ea85f022ef3a2fc937ef105bd73c97265e33019f43acb42101c1a7e9dff0f33e754997def0123829d19fe5e6f59bca4d57888d3532bdea593d3e064472da9c96b47d32d9757963f439b92123cc8d3d8158c1daaf3716d49251beb83a584e350d09234c523a3638cdc0205ebb87d022962b3b913c44faa419a5c2a8e4426ce0cad1c1c0605638eb302f92cfd7ad468d3111fd142605cb253071cb96a41cfb548b41c2da12282b8cb6bbd09a4d09598758a100e0dbd8fcedd473eef1690bde5c9d5f8655c9cfada972bd133f5208837c0fc64e4a32b7780a49e120c4b678473f7ab4e2566fac2a876f535987cab833172461fda3028c13553a418929b7fe1892edcd68dc488742702a17dc9cb6d6a02ecbcb2d936bdbfca232e78723ecd5424e0b182a2fd6fc5f283f06aa0cccaa5dddaa662a571c8cbe289030e62f0efb6a6ad2366e424f47d17ecb5b60b7e44455524b0e45f2040e4ab149f4b2fceef2b78a85ff4c459b124837c1a5103105576ccd22ab06ec783dc3a6e875d76c607e584a9d282b0ccdbcbe26509a56f25561f824362c8c54f4bc9f893bbba57c214dacfac4066f73a02588af2b9a452cd6a6f93de6dda6a856a5edc1200035c8e98da7b4e9a8784a8271c2c2d8341d65cbaca36e163e228d4f57580c07ff49c3bec9988dab71e7a043f291a7df18af1466f15119dd5908f9fe796ede38619814f3f53b73f0fa7f97daffa21ff46fd77620bbbb12b2f588231cb484b5e819e6e02e5c4a9733f08aff51783c5e6cf3dee7e3c80e2c82ca69d42b135170b6c02c91fe776341318e76e5b43ad664c451360c9c1177d166e20025665264abed452ae61fb1e0f8ba191ef1a4efd89422a5e22632fd4011c8e764e7756798f12f7382a6053fc73f062b2fd15d400d0ff36fbc76662d0992bb210c1c1acb0dffacf3d8467d9ec2b8c6280cb582fb82696afc7ffaf950d804652b430e0755fd98cc3c22f259490e61e4b4e161c4ca6e2a806eaf0ba28a77376b3395cb05b04fb405bc7d02e5b8d92;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4df8442a5be310fed1c8ae6b344c837e534d8d61d139dffa1a900053b5f060a485c8cde9dec715f18d0e1c33e422bbb95f8cd7da70ab19719a1aae654677938324665fd2771039080e33cf5d6866bd49654f7b1435f8649213b53ae76b706e900c8be21884b1006de139fc8fb5610c5488d3161658ad2695e7e581462e6dfd3dfbec83230e14b8bc7721df684f8337b9df370c6e78c09c729b57b5293dd2f0439afc9b65a748789fdcd3d49b3144c10da6eded950b14c2c68616ba7c1e3998d62870c47fda6bf098dd42ed49caa96142997a3d7671d49062b0c583022dcc092a43201c9d0119331db290f3cbced6ac599243fd7f0e99a30b986efe681cff386603c1a4c4d1f42e64b8f9327013ede966b8eff887097f0f6f9af9abab6043502356b213461be3307b1c834183cca419feeb050425d321a45ebef234b864be5d8bb3f5bce8e64c8d9d38b35d56e708438f7be246707e32a3fd91a03779ed897b538899defa56633e32397c603caf6bfe5e46cb09eab9c98d55819bd9351ad5837b8ebf7640da3d19f13b8352e87b79e43d273e8999eb932cddb4bd4613c9f79b1eb22b5ca1c3e49bb4fdd717cd86b6a5a9cef5b5b4868df64309d1123786d0c3e55c592c010a1eeae14f88245967bdf4ee2b46ce8ad1bf980cc17db7163e72db07fea1e80baa078afb6ee7b3bdafc0a3fea4de24e05a69fe1c5786d64c77b03809bfdeeef4a6ad1dfb68e13766688a2197be9e0cb858a45978491abb07555e6e3b4b6822126abad46a4e9c9ebec9d89f23a476006a403782e2819e9ae474687f5be7d5339209609229a28bcdb49fcc4ca933a688480d2a85c6965587c34e146cae40e4f625c84aa42fe61bf42e5abec05f7b43cfe65fec402817ab740c3ad11943fabc43bc78504224837f97335fb29b11f20fef1d52efa4e227492c951c390cb43efa101673da1405ada768cc52f44ac2e25a1d7547b1460019f031d7fb01d52ebc364124cec41c044166ab4049f2011236cf0f787d4f862a73e84fbfdacd9ceced10eceee16c84858abf2c9358e74921403a79281fcfffae14e0af53b1c1bfe699e709011a8ec19e115dd10565fac9f85468c0875a2919e39919ed029ff84fc1408393d42ed49ecc4e765f54c6e6b940a9ca7b0b49f6fdb944543a90a9ee112b5e7763b8357b975e98ca93bfa2622a68de49cb03dbac84eac0b37bf4dff8e01da7a54306db59a8406b64a8845bb98bf8d9b1b22dfa153de65d0fd609d8f10be5ea7dda3a18c5b2cccdf53a5702cdad252b395277c2dabc68380e983395a8b656929ddc4480f85de9ec95cba9529260d59865c9caee75889e5959c67718b41f8da04c52a88587d9cba2a250c7c10579cd50a922d8c74e4c472b9db872bd247090d73c84b3516ded663e8c4f33fb55e687623cbe487e8a993698ded9d28603d7cc32c788f289d6a5f4a00582c8e357ece0cc1edad945a46146d8b8acf0baa9495692219d7fc64db74c01f2a79e6789f79545fc4817deb3b980e76ee34a14aebf020a77f0c9b2ab2d8ef43057f8ef59db3eaf1c2085fd7a583c5409c268f6f34cbdf53bd3d93b8a55bbbde3c2a357c182c9cd367b7746b2c7f89dd93cdd9e2f4ab5972aecafa3c2a301f22c48ac2997edaaeca94f12ad9932d8853a8b69605791862f47e3a26ed090b4ef112c88e8c38c11b1dff30d879d809b06c6427447c404d6f9e69118ad02e9d4bbc22030833e067f6555ae3a3d324c9b8761dcbeaa9d19ec461a15c8d7d2caf0e933b6193c82326a50486032c95803e3ee9882ad24b18ad927dc17d0a989a876541db067b06ac6942d7ab621ae9e95597838c29e55e2e077884ac627744eeac82591c16f7772253b5cccc471f223f2542291b6a81b115177f19240020055098da8caaf4be626de9135d920ba1bd2185a715ee8dc340f479ec4f583d3bda0763bf3de6a4b1b1a5830d2f314acd64ed360447e6da2a59a91cc4d229198f3151e5b4a4035996eeeb3fcfdb49fb48dd3ae49625406cb6dbe3309a13a19c23aeb37a900f281cd27569b71bb43123bfc1fdb6800073cf362e0984f4adcaa3c13d8e00842b05723cea2bb7d4f0cf63eecbd20635c95342efd15952386483fc97d45856476fcd6cc6e409d8094d434e67d4c0164381acbd013ff6b94d0804eb8aaeaea378cae812854b2dfd3730007f5616ba149bc3a9f81e6c89c4ba6dbfe7245ab2b0ebd586604050e1448e70faf77b017b083235c8853a1cda646a58312df893d3101cbe2aa405c64c4973548ecf0d7230193e2b3e8f8b55fa28c85990f18a274f975517446cc352af5a1ea79f1106a0db7624ba347622290d785ca84ab1382d2b87a3933c0afcf7c99c753e67eb4a88ba70bb132823f10f2ffa593630c148d438b38e28cf0602546650a30d1af46644cb9d3bd85249464f5f8ba865ff78bb88b573d25d1214aba27bf735b8401125bfe33428bf02a235e3eab50985fd0458f1c9f29b97db34135586566ce69b0066f4c54cba9be4839d1e896e7757834c299dff1276084c486f56f3ce830c659520f8605fdefe988876eecefca4e1d3b9cf396f0e252e31b1259bcb85502e3e6b1a8fd86b979704a355b2c0729697557f2cc620699a8c22b7c601f00128278225f5ea997e65b5728c6088060fd5fe472f926ab24816a29c314bbcc4c8cae338f89b8bb0837637a13b62c3bdd9e3f0896f04c2139f63a412486fb48774cdc8fbef7542bdd681fb1076858cf9f4f5e435c628154890af9b1811c6c5d3e1ed75dcf95c364053b79c62df5d2832a2bdcf4b1407c35aa89ae0279a6ce27961234f9e13cf77f7417fdf0f11d292f3080ba378f13c6a7e3843c62943c6f0b14b125391830d17278ee2b834e5e6485d58f74b9dce216dee29f5df4c113ecba8bce5331c10221e55c3cf354dc3fa7bf251d8c6b6edf00f90cd1514b29b42526dd0517ecb0d3ce55b4e385598ec0cbbd958c979a5002d0d824a2291162579c1122017fccc6dae091ed67ed213977c58999906542128621be46e1081513f686c80cc708fa98dfc6f9b620bb76e1510ef985da92ebea7b6b8b12e093e8413a2fe15b059cf48825bd0ff4f6d0ae451c6aeb2dd7e67df966f1a073ff903569d062a9bb0e972b4e862f7306084c47e2d79379a03f55d6d49703a670d1dc64bca989a9b17763420c3e93db03818401ca4e679c5c6a4147938883cab38d03198a845abd91dcce6ec0cec8dd4dca16f803e660267607c2c03e2e876d5bc4e755aeab889c81a0dd6c6f25f0577b4e5599b0b33fa3fc53c6d07f9fedf00ce3fd5dd669da7410c4fc6473352d28ed7d8a2c5cc74e346fb50eed2127c30722a5abb1718d09ad50d62c0e42128e461d3939ebcbd0ad8aa0b41ccf2d6b1e517e704182d4fdc76e9344c84b9436595a70dcb70f61c57ae29af13a543f7844ac4a6428b991acb914e871befbd747f54eee634fb52d69f65ba79af6177d66dc0c8d4c38c9b5d4c9d1a9f630c482421bfe6dfaf1e2355064ee4d2d5e99f24a9fa249e74418f8bcc7d4ae68726d8a2608a0d46883086979730ca4040874e9a9229680d18b117476985aefb65aba096e629631b69afc404eb600d08f7d6c0127454bb2d81e326d064cacf2171f3e45fcce670e76fdd08ecc7727648b234d85dff6e6689260e7cceb9ebfc973646d0960c81c76fac34a638dbe3df6c71dc6c13e59421bdc3ac170beb8512eb9ca22746349f29b3a447792a46fc1f63807b8b0a42976d2dab4dc4b2c12d71829d0c3e08df00033a9259c292c02a8563d4b0cabd115cb848476f0f52ab05932d646ae542aa8e5a86ce279659ab43810c56bfe0dbc27daa0016a89d12cac3d13addc1a2c96020a2507d31fbb285322e83e91f93aae48238a7a63b42d99c41d47cbad9722e3a3d6b55ee1c91e9fc40d1b955632dcec1160f3743ba6cecd5fc760644d281f25591656f79ce8d3f2d07378d74ff2f4bf12796f560009a55422fbff2b854889be48515b3e2531f105a0353921f8ab68ac39b900d1270cdbdd72de61fe054f7bd2877177415c499f5d0c0f9cc19bb8e07e66ee4d446c93c7d131503fe6dcdfdb2f15215f86d6a09ff9edbe62766b4902df9b3ae994d36248c8d6c72cc5a4aa9fb4a021232cde0cd1528c351092b3226e8f6414daaef3c88567f085e3adb61c199d41a1b6dd5c8bb06c2c40aba974b777f9df84d98ee26c816f74718e670053e52a21321a399b1ba88c26e7f8222fbb2bfc0360c00d98f165f9483b9e6ec173f774f7e14fdd9b52a97c76b65266fbea12b74974b2300d8a603fcf0de042b0e618705c4452eb846dc31594ad924fd017348f0f47a565e9d518c4b33751500b5760faa3c2bbb7c9e9024bf9c395fa76d09bfa0261bca6f20a384f83d1854edf72a64a888ac8e7b19bb70fa875ad44d6c35928ed553eb85a361ce8753812014427a4209242b9578b8e4f33d63a0349732de3454ee70effd6cbf34465faff4023920342a489627a79f4aad1fff404213cdf00988e2a1c9cfedd83c30b6508782c4be61c25e525a2691d21dbfc27c319a9b9f7dde98924d84f8a9447be54a309088fc9eeb49469eec797191c8e2349c9b41264f7029528c11593ea9da7e71663b8d723edaa6fa7d0b495945cc931c69368b0fdbb103a368e556c78504ca6eb47c089f80027e0364d8e970c6a634b88edd7295d2cba293e6bb6fa92e024a0c3354f872b54a1de978944319ee523245677158d56e5fc026799df2b894af16dca71be93624998aa101e7422c6663db0bcd232de3619a24767ee41752519e2d3a9a5143b0d0548b21542f066f42627cafd40529e9a089d8a957655f84d4efb77733ef0396956e94351101207becbe27f3451fd1120928c121351ad1edff84a88117defa3f9d34b3797b1ea3a961322844e354613f066a396ecf7264195654a4b422ff642a0dcd58267c4efcfd9c6987087346d26d6e345559c91ef59a335c990512084856c882f386d4d587d2f8687f3e2003c98ef9d998a61712e09c3648a8fadf74f4ed2f0db52797f3ee754a791cda37f03649b86a94537bba0ba7cbd156d0c5ae1c34d88ca2d9897729369ee5e4134d951a423a63228c44bc3a0f77498c4dc8b9da9f3c88ce9d93c9a60632b6980e8eb979b410aad576a825ee5dbe0c5120a51107e5768ea48dc901c9d9ecde238fbf06a004e51d5704cba4c01707d20cf02127f172ef5d85b22a7c6cefbdb68784d44354003ab8825968efa331f81598753485c30068f3a938174057cfc2f464af8e4b613e4dc7abd21ab70cb3b3f2cf4cca620b4e55751cbff608ff03d04d060732d63252943ec37f4b4dbe25b1889964752cd604c5660a3bda7f9cd9d5656528b37744d373db45ffda997bb162d8becae3c67175e2b49dcdd8dfcda6723947a637af63875e3544d5b8e46bf38106fdd696667bdd001a9bb7614e91483e80e3871b446bf47a31b51f6c4647d6150cfa0b55561b121376ec7d7e6ecbab486c6dea019a1c23d31d0fbc508365fe7219a7ce2da3ca2f8963fe81df9082cbb294a086ca9f1b46d13928229ad3e6a5dd8c46ce3bd4c948e514176df714e1655baa891cc487cf04cf142b92272004861ecac013f45f2232d321606db5f5bc4b086588ecc39ba5fa4a6fde51d0a128d820e0337b1f9eb4abfe7cba5165ac875b24e8911f39d37420d38a88518d5e2524871e16b8328d6d936d7a26cfd1bc298971951a5adf61e79fc3180eeb7953af9f66ae7911e21ee32a35850a0a12d47b7b6616ac97077;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1fd7c881c39d218baa6d77500ca909aa2ef78b43e83e5cf3c3d3598510268cf7200a13d7bc21de937d074e1aacefe3d9cb66fe05a133014cc723350f8c83addce035e641779858f7be571a07413c0709aca9a7f0cf68bbc30470ac74ff9ef31389c88541317278303d7bd8da1385bede9424938cf19301efb3cc1775d8ff0f0996dddc5c219df927549e8972cdaa60a1c7d5fbb9d1f7751d2347e124e5cfd994415801da3ab961e667b32ff93cdb26ad2d0d35d62c1766cc4c411a6f598a77be5ced5880935050d28a9a3246829abfb2419303314972c84d1a4e5d86ac0d4d590c2eecca1bd90cf1c202a0c4b9e956210d0e0db2f9bdd1935eca5b252bac46180ba297a2b7c828c1f2bcbdfeae56a1764f58148e0a464bc8aa2dd5b8a594b53c40cc4c8b6282cfa5ce335275b5a03b56f438b3f84342a3717569e1a2cf583bd2cbdf6f72d72bb930192bc3f0f45497be4a11312d5e1ebf8ce333ed882af2a34651d13f6acc0ed9623f3b90f53e2488ded658cf66ff1ad54915ce35870f5efe61eef799bb1e55d07134986025b252ef25fb1269cd0082df88baf3f15df16205a315b1b570f16c60e95e3b835cbf5896fbff74b62bc73a9987876263be3fed51d6fb3b429f5b88be75caaa26416cc9cea6593fda08fe22f7e7b71595a4cc51201f5de65df5942b8a90ae638554960f6c703c818aa68e4497dfb8aa2562772ce427117aea916eeae78ffdbb44acb0ac5fb8372a836709aba4dc134f6438e4c0775cf6a301cfcd8acf2c4fda0459cfc987d415386d98a0a1ccad386287ec26c858fd355fb40eccfd45b435607a4d6aeabb03cebbba47fb22dbae5465a2979e13671ea900b5139b7cb63307dd82951318b4703d8fc72bc1d47c24e5de66658cedbcbd08a037c96ec770531ebcc0a06291e73721892004a7ceab46174692ff7f16160802a428594090e291348016b4c7a367058b5abaf94c1d80c8a51f13951583fbdf80d3e910f27278a085894e6ee19921c05a1584eef46be733944064169e8a03000e258d6feaf5cb4ab6d3efd919251067663e5d86817018e1ef2a853c368eae8bc741baa144b1340518194bfcee6ff28f7ba54c9ae614bd6476678e584b33676e62e586e4ccab4db1b2a3911d762b3912e1b8145296e9d2125d4c5c3e25c125d9f1c9ed39cb949cfa5c858aaf31c13fa655aa7bc4648099b8c1d17f0e9c7fc7a96e721b7062b42a7aa48af2be02c866409d4c3cba55a2ebf123e78be5ae3b027cfe9434894b9ed70f2c72d4b9b76540ab0afcc2f8dc475b3fdbc809e0aca651fab56405c4f89d77269ca46d3081eb15e01198c2ef8ed38fc15f6b0704c683ebab5003c74de5b691a217afecc965f1e239205b9d73ba4f1a93c4b31dee02ce1dbcf5229112ed54a591f521e71fff6d1a0ab8ff4d9802fbccb150eb9047584cf677404000c11d73a9c67a9a4577b5e4118ad0a06fc628f346441a53ee69407458d078b8a79e43a1d1a7a1e23251798d19ee8a0738ceb96dd65ac689bf55c0838fd0264d6535b91f98e5cbba4722743409604072813fef4a748daefa91a35bd668100587d46bfbe7367006104e7f1fccd16eac138f7a92d15b3ef28b97edbaca7ac063d496461ad8c47d6e91b1e4ba67ec210f9f280adfd2ca63742bacd74bffbc3104897558ef0cc2ddcae06b39b06f662d94a035bd25726d468fe411e9ebaa4f08a4549f1a8520e2b67092dc7619a366a92b6566a9890a639c5b20de690d6b83d10707de600bf17b0e70ab8151be66559a83b1f34f39991379d209f2002a87f1df29aca97ddc1e0b907d1ecf45cb01da9b9f6cfc9843dc779b1cecb00e8dd6fb6fb274d54a2ddcb7813bed5b49a27ead0b240c7cfbce509f8d755ec963cc996ff2ec34dc017793d0a893d8196cf7f7c4cc6a752cfcb2009d0bbb74d37234088125259fb2349a793fc607a9aca94c104b1da75dd593bb551f9c75b144a191a219134aac615aff4e2ce0bcbd372935b35b3f3840799542c7f571e986830645d8150e44fdd152aac22121c37d3b590bb34a51e19d19794b6ad751a06d39d9229143bb97eb4a16fee694deaf89559f4a7c3c46f37b45c69dfc4c95314cd404a05cd040e7a173216af812b7cc6b8d2de2b70e1d32b683065e007995b50347712f10ac6883bf4d46cf4279edafaa1952014f2f6de49a6e74258709e9a3d7f137caf464407a0ddbb41353c3f77bba17c564f540e89daae8a669bd4e04060ad054f9e47018ccb77acdceb079eec7d5bb931f01d671f276b5ba8c76f634f63cb10c4fc5a3e2c29db107124f52e100ac85215bce12ff995c29bed34044198e997d92f3ae15b0033c6b581dcbfccc74bdc245d2152528afc0f0f60b9edad5e253cc32b510b911c9a380d05fc07dfc39238df8cffc04b2a8b2ee78f1edbb464a06fe8d2041f5dfb70b9f75f6b747c3b32dc4df043082412bc96a812537877ee72a1bbad832ffc20a30c1753006023efc692beb2bf16f601d50f4a72b6e1abfcfdf62db4204739f7b7612b5c260e904c52ac5432b62f6c5d4494a436e21ff8b1364a8d5fe9bc731dfaee64f8994c3f019322f81e19957c4918e017b20ecea0bfc2dd556b0cd63b5fe1eee1c7bf3791f79fcd86f1024f376bf3ecc8c30d041aa058a60939005d5023e32275a15a785b579e3089364f5b3554c08cb5fdd512f976b8a87598612c0d862b00d284b7f8fda4385a2fb717618b0226541da1cf130d8c063add6486785e3d3904e76300a9ed8af1987768da32139846d69848928b3e2e029a3c2c2fa6c027a5ed3418a2455b0df8e4ffdcfc1d46f9aefd0bf6dbd6d12f8580710120cf8e906a5973d79a9348cda44d91bee7d8b79114f536e0b5b57c93e881beeacfaac1e0cbb67e4f96c95c6e11ad9f622870ceb712483d9cad51130c3182d41a594874e3ad87204dea0e0318f3bf38d9b1ef1f3f38e79f81c24c23682ea9df9025b865725a90891fd62c88647d388588cc6a9646141e1287835a46855be62f5acb1d6040633b0124cc072f5dfc796b499750cffd6c052b73932083fed0576e967a5da899b6fe5113ad6a247d75c3554a49c76cd25e145f86ae6a7bde70cf6c837c4b43b3a4704a994eadb7d75a3dd2c78827fcd8936969c9ccbf6172c2daa092034018b871462cdd98cdcc2babc30e61a1532e54d0005e8bcb27c9979dbd1eb76813f612ef2ac8723d1e9a9505bee45af3cc78f7c6e5ce697349ccd75e69e05098366080d206eb7d6336b392db64965944d0da27081462a0a92ebe026db6c34568ed1a9a991bcaefc622317e452a26d8692e84e5709267ee0bc535c7d4ddfbd1f2666c32fa0b72b7fc7016e9b39ff6d844a19c5c028bb010158f96cac8b6ae289acf96885ce253c4e04ed46fe81d4f512a7e6f6a76cf82e08c38a2bdca57783f5f847594b9dee71081b1501ac18776cbd7f6940927aee718f405d8391c7cadcc1b8bc556df714373ae5699b3c7414577d82d263331ca64f90b8d8a82f869a475817508860ea727fd4e43772dc43ada6734f410856970bf5f0fc0cdf10c7e27e87cfd57e43446cf57e34ac43d7f2de97851c5fe9949d18bde6a40aaa516201654f20d05b36c7ddd8e132a9e95a2ee102494f60781595edf0ac74e4c4a15f45020959e59227c06d666ade2620b70d7054a814e646e5dc39c3e83708b4ca689454472b83fa82e2bc768f572a8f3b26293726930d2709ef23dba045a0f7f88262af847e8c1dbe7d258215f9895674dd3bef9fcdc4b8d52adc94f8f27b9596c37e83a5572fea66f172f6f68dda4f3038cf1c57491d205930937a32f950957d9a6d24910f6de8097da72c6ddd0eeb0e95b58d54adc0bf5c8b7daf2eda2c1d2c7a96ea1f8c5a869273c0b2a11d70d8a6c465cdeb9a98d9c768e89c418ab5381046343333bbc8e104e67d0a74b316785115150aab05cc682b36ab1056e46934f2d7fe98168c3f2b17e34e6d21b003b77961b3de8730261a40bf36681e548fea87e12a682845523847fbc36927a24e32fd6d8ee29df0ae60a7e0a34b5636ee4ba043a06b0b304f7624e43377afb1b7218bef28e00ef8ed8ba8569debe2bc6d0054516795b0b6cfbc87be397b148f5ca6f6b47e9f73dd94323e8850a94f0e4405f698c9c8b59d472699bde902d1867db2456399bc77c99e2102e1bd523cd297d4216e5f599f3c1364bbb2535012e93ab07a7204e0ed1c50ae80acf74674a1b54cd5ba7f281effee876b15bda54d484e45765578fce3d21fccb7e1d8dcd33498390b60638d2b4a3966c33bda6e9b21a280112daf02c4095c83aaaeb66a20aa5e0c36e4615c2d53a4d5fe7d502beaf27842c4854bee0b5738ba1dbd7331c57a2ec21a09d2d83f6a5c8e8cb5bdb073ba56927a02cb1cec1a044fc7ba8a9f2015eac966a579d589a72fc44ddeda17f456d289ec28a6a8ee00ddb67377724bd7e61c6264fd99e0b7126e8eee6bdb7b10e0e0c64399a590dad0b33b7ccb006c829932149a5496a62b242ae34193115268a8ac73f278d4462b8c36927f70a14f3bad33915261ff49c599ce335929f07690b082f6a676a32806068925b1d6a0214cdad1a692109e81fa02b02b82ae146772f09cbe694ed3b61b7da81280d69587caa388b3fff0a2cbf5b41c5edc2a6a06d647ab92131b056fb9d69d80a0b95a822504e8472b11babef317f9da4bf3e6a543f80e84fd94be2991b2693e174701810cd923af1d8b2c6da295f1567189be2a553219af6654aca80bc5e38d6bfeed8f9aa970b9c2f9f0c9f549623086e40e595084c1ec48aa89c53949cce173a9edfe1f7fb9d15476a921c587678d37392fefb6dab7f7620be40c28759303b3f03d20bb8879982424aa3f06687bfef35c234e2387f99915a78001cf3dfa10f81bb63803b421c29d5ad09eaf5f7621e487ce81b2b1390511167d82f10542b7fe59878085930806ad9cf59bd49346ced262c1b80bd5088c2ee3f0c210db8c1e2e5bef5120b73c70b1631d23f7604809c7d9f2d7df0521c34b2a88d23d2cf12cb42776b463352151505171c8b962e239a4b20ae1c39e068553d5c63044f3613c6911e25394297f7ddabbff70b7cc0eaa21e364034d71a506c659e5b5291b75e920731d0e737bac694c20d99fad3b473d8cc52115ea496818089264c81c01ce8ca2958b6e7e85f03a199791ed3b0102ddedf1c276de93b4593808727a3e14103eaa1280468047618d5c7ee690ccf9729936a0faa441bc5780ccf0c60b33b576dc85f4e2ee09f13035e236b190ef5352d22f11243d84c87cb0bc3c6bd8774d1c46fd39d3657acebad24e0b9d7866ee7bd1a5bb39d280c6f8bcd53e2b6ef1fcf0ec56029f28134ee4b6e81333aba6f323c806b1d1f1ebdb20d8dcd0ec189dedc6947a6d5138e55055ffe161c7f0d71ffb9e887775d5933e5310e0879e6aedecb2ba6957e4a7c90cf9267992828ce7c004d6ff09c81a7dbcf4e9ab7d7d9447466a1b144b6d6d6d5c6da7a18e25048a75b70edc521ce7f8cafda5167033bf62d41739c9c2de648546601335c1b272241c1988a4cd937aeed5e8cd8cc88387fc26af21751fc4c4596bb2f3a95db7ae5d2f61aff9a016319735e8438606663239e6b25c1e679a413ee4d299a9a80e6e2b3fc9626b92328e199f21adef0ecd767aa57db1bd0e6a56e7f19283597323d0baa2cb4559c4a6c66cf98afb0a34f139163e394eff1181d264018441c2d698db0e1e23efc224c05e46add37052c214c4604ca882a8331f43b94190eb7f89e5cd2e2a98fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1c63ca14e37b63d543fab32f2ff4b91086e6ee690f973c6aa676e4978f3cf2f21ac4e1164701411d4c4956263b684221fb3b67326c8ccdd5b7840040011ee12122dd5b01e57fccc922d44b4ac4321814e1dc85dac4c398d7d1926bbe3a6aede6155b206563b8befd6337e9a2ed850d304a2ee7477f26e77587c1c4d5a4bb55456988c665a730b689ee100cdad5f64d5084891164519ab1e04525c96616cf5950f7e50c01af648c1e7a9cd1b5b3d1b5ee51453d2cb087ccc3df26755d2976ae643a6ac1de78f9a555801c137a656914505459bd7c5bc290dfe78714fdd70eb143e1b8fce635ea7c2dbe6add1b6b5b3db4db173c4dd260d0cc47865f622f18c5f001ecf0a29c60d83fac4ba0f3df0796891d665f24bf44d74c11da176bbd2572ee84f332305a369d333ac3a6b4806103f22765315b04db269bdd75adccc6f6f5788a028a3304c4083cd19a248945eead896df43057260787cd34e90037f236348ea4b0575b84d124beae1efcf95e89dc9634318dde65ab73816964d85c174d8e9751b87f907a8dcffe6aba463d529a74b20c493f34049fd7477cc5adb98914c684107700abad90bde4032ba0667f64789ebba255ba693c0bf3807d6e21f7774ee7f311df34234c4dffec388e20c4a18091bce8160e9e2d43b2129859163eb329df7afb5c73464377b919be8b2daf1085c2376cc7f1c1ea0a636e11d57e058758e99c67b9491fa8891d4a493a437a2ba6e168a650e61a2f50738b063763f5a1dece2d861e0c193b3d2541cf740b7f04a47cd7f9248d77a1c3f1e9242c7e224c35a8ef18cffdb6e6b426db95aa4763b999e852038ebea9ad3554612405f4991923df5201ba4fe87093a30fc06868008fad6402c14e097933d1773f12262271073e52cfcb0b1c87ccdd6c73a6aa39eeef0c014640136e96fdc71307f292a783de21d8c3ec6665eac0d527b9e45cda1233da0dd572276944b98a5696b705bb6a132206a4d047e976aacb679ca8318f3bc1b46994ab9c320a438ff7b0411ea81d1678be27ba350b8bb82acdfda4655978d5fd844591eae45bafc1b7031eeb071eb0a4a036d6fe993c08bcdd9aa5f327400ca621befb3245f96141ba5ddb1c5d5218286a52570b75ad17178dda26747276588210543e17e54aef4d849a0efa0606b49ea6bdd490c77607173edb3fb630a3646c3e8b38755b9409e5f6fb4f29eff34a2d929ef02968c77a4ea5b233774ea92d9a52f131b4c3374bda35ae41df4a8de34a8b6d10c8014536a2118a634533a49ff9951a1bb79cb2e2a867ab631c2a8e8cce94d2c347d139d7f03e55de3300c02aac4fd6d0f29c0de24285c73b6cc282879969d073db9becfaf192419566feb126d853bdca149241671e842d6ab441f9098c835ca3f01cbe5ccb8435296c81d0c1d7303e928a100869efba08d6f2cc1422da5bff3142f6467a74520c64f18aaeb48e540bd33edf5ac398e69adeed2e44a5586e2e84c5b363a42da7a1df4274b758c003427a6f6f45283e90832fdb30aa5022de76c07e7fadae7ef655936bc4273e8f948b9093ff211361cad5d671dc6857349232245f68b7cd73049ec2e3abdc0b458e1b19ee7df3bbe83f2097cd914777a304f25a45a9cf65c59ea8e60b96d93c55a1bbf9edee5b274d2b5bbc6e87e3ed4dc8eccf86fe681a0fcdd520d22dedd67494a6668143a07266f1b6cbd89df3f65c19f17942ec47739852aa303d5dea6e5c19124a9dc61b49bc5742afa01aa4e6adec9cbb0d528b8a5b2838ae70a6ecb8ce72708f98858657c4a3cac86d69382d378a3c075b4bb52fb59f60918f3dff7d12a8d9e4ddd6e2041d97bcd2149a2fa437996eab7a2134fd11ebbff68ea9cf030e25c21fff985f26568c233b0fc6f109e0cd3c9739d6596c8e49edd7c3f6abca36a10ec44bf8f609053f32787affe1be6941b97c9bafa74188ac63179bcd4971f72513df336dca042257ce0de47486c620fadcba9503f8945969c4b3d9b092674d90468aa7f98606923bba0b56f841bf4d34e44a79582e694ecc7fdc33cbc0de67ed73915d8f4c88f27e49945488f4f7bba2251db58117c74d8a3b3b5f959b3b38465201e1661cf281b015d0f551bbe36dd33cdbf7c1750c59724fd41c5d22b8855b437c3e66b07d2aae60fc02fdd335ebd025e3369c6a17ef74aedf8921f08535250eac816fdaef483dea5fa49415395ddcf239e1a0732cb3adc06e659f2e78039fe61649c29f69e70ae7299adbdd7ac8a8b71f9d47c0cec010a239549f634e941f673a64451ae30546ffbc6996bb243779f553d621e85d270a7b11b7d825c667786123dc6ebbaf9985870108c8bc721f874db96ebe17eea7ad0b04ba9239e73a2b431331197ef4abfbec6dd5665f5feac05c8a006605e8bdd3822305ef8466a3124da0c5804f8dc1f0c0eedb34858b7be63ccbd4b1a9b73cf6be64960d50ef9becee911d594cff703ce8c380f013a80f83aa4e0b4701bf298b7ec565c261e922b2fb5f8cc311c8e855195cbf96fbc382572c0894924340880cec8f741b61ce9cdd73be524c5b54713a206a77a603991d43a7fad972a536495a1996e05c74784a9c428f9cf100825201a1b5af73baf4e22c35bd6f58b3d77072395eb1a6ef45a3dbed7b70994796ec321ccbfd8083cfe61f9f03ca8e3bc0820a29cd7c3a69c8edcfbc56319fb2b58cd6243e527fd6e6a0aa55a6b8ee3b951792c43d9197fd398ca575ace34a91a9ee443f2f4b2a3e41732f15f79dfb9b4fd1fdd099604f12dc8233c3c5f914323bfb45ea294a9d545977b956002babe2c0e76a0d26934fa572dd5eb44923b14bc1cdf7435453ddebbef61517a6e95b0ce4067d09d99eddc0ae9f71ec4c2f6e30040e0c713eed65810cb1b8591709cc7135bf0b92358abc2fdc0c03d2aa288da58986a1d489910bb7b97961244589e9c8be5f3ce894c1a1796ea1884ead6ecd7409d35e88a4e5771345ba1989335ba988f7a033db23347fc51626718ed231ff41fa74e6bd4109cd5cd78cafa60a80a8780428cbf8560480d06d5b157c1bc79e244c8448ac2018d9379b06a9ca589b8599783fa874fe746112dbbd2ca38eba3051f0872dcb529f50ef575ec386f74e910bbe9a327a690832d4852344a35f9da128282f8def455c940849aa4f614f7c0b6815ac838eab31f57ed7ec5a9314483ae28dc23285f6fa3fb11d236169427c26b396c5f6fd6e19811dca9ff7ce32122d752120b290f7a647c49db3b6cda34cb84d3b3209e68a66ed7662c4158f2c6bc697b3d9e4d9c03f0a7a788b1cbb9cd54083feb559433834cb901dfcae35758dfda48f6c4063da1a9f54805d4619fb7934c2cc58bc2b4517ece8c970e38be15ee871b841be3ae6847bdf4e3dd3c444a75d2b870a119ca7a85ca0dd286f31f258ace876ebe2f95395e70e99139bcd2961504bb528ce5fda4523c45e0ab31c527a7ee3fecc9de3f15a41ac2b49c7975a276553c829a0bdf8d93feb18cccd33b8c7de673125af84180bf7f72bcf8bf1b7897bf0713a0ed524ad648432ccd6d9430786d773626b9fb2b049a37437040c0914fb05d0c8f27978b4925a50e6f4f49bffc768ca2d1b118d6abfec22ad6db90fc2a98d3a683c84b30d24fab0b943fa027b3010654ab96c1cd7402e6e0ed9a3813e970c41c3b2ce059ecb1da83b6151ecdf7c2ba31a1dbf194a3ceeebc17064d2c6d191db2f5f4ec93dfacc627834a2bb6f897d2d258b4f849636e1142815fe2bceda05dd79d38c6a37e9b906143edbae90a36711ffdf3c795b0ae6eb3b9c79f6328e3aba835e69a29811228bd45d3c3a5da53c03b1ecf72195c325139475dc0becd54cdb36b7bb10b372b483459e801f3ac7b83aa6a2367cc2b2f889a05f025408fbcadbd2b6476d32ab9c1ebd86a02a0b88da4dab3074c2e0a902a5d178998340a85fb1430980e5fc89480b4ad784054b3ad4303211beb7e0abd689e0ea2b648350708868e0ad8933ef17f69b2971649507d1722cece984e65c694b1539c7ace29ddda0aacc7117acafa77c0b7728c32e54ba663a04788a8fac757c21609d34e2a5a1f01b7de843445da3a34163bdbe919f0d778ff0c7482af0e4afd39c39ed1c604abc797fa78e185f599f01d6e9137cd1760751c8e4d2af65192fa837c0087bf6a6929ba3937b736f26e8099e17101775730e94708e17685879f9e909e3906b8af3c626e5a89f21d8df49b02cdfb18ea0f4ead64215554e56dd7df8c482e979e780c1c7c5ee0cebad4dba645841278d2a7d473797c14c465c3d2d8b1c735d68dde5da6a1b1524a7f19a8ed04bffb72a4c10fd81945af7d75a95a1481e55ecf5845393398cf385478179c47c523b2c414d0c98f0251bcc53ab885a9c6a171e8bc7df5485841954d073804ceb4e2c184b9da5094976ee733a94e24b4a6bdcc09b9e11e7b5e14ff489be62d98c72e3307eecc9accb3ecfb4838ea9983674ca18ac143472d9f95ec50da9349d1eb178ef39dfabaecbbbf89f670d7946335b932bba500cec08ae206648fecabbd3eba529b56bdba0308555df698dab2c5e3aec4e922527120b7a5a7982c9f5f6c27211d0e850d725bef45b190943397b499d6937765193571663bdf276f47dddcf87bc3d1e4a6bd24cdbd5ba466dedcf60b14930173bfaf3ff7d1fea2efd2603d15a55e6a400b105114583198cd6b56454b96b11bb6afd1d71844950ff2c5e801e49c79eaa8b071295492f0b9c96cd49fa416a23e85780122fcc5013269b5cb6a6404ce4b3db3579ac7de86886aa7f19981b17b086199c5cd6ae3aa358be2da3e209fe4f3e10f84ebbc7b93ef848e3e2e00529bd3e4b3ec78623fc7d59b166adfec9867fa61b202bf226be9d93c521db9e51d85465e3ac4975852833ff53fd078d5e970772e657c5630d624bd19b2126d876a4a17d3385d552178deb12aed93a8e2faef84bfee00feb037fc0914b6e93de122b71a4304e08e3d33e791dbb18dfee34a9d1a6e227f6f1a16362fbba24720024f46e6c434c33d1a72f6ff84c65473be1d5ccdfb7d8c82f439be0de6974e07aa3c9edfc07d170ae3006d9130c50b6c7fb4741e3a93487e6fabe0b5af6d2814cfdb5cff061bbb0c3fd7ac871e2e950f1f29958a0f0f8abc3c1311be4b79e879a21cef08f6b48b266fe21da36c2f93d305d38b451215d284dad562541c62f7b2ec801b14800fb735cbc21472938000bbc25d4811b20f16dcb326ee7470ae020da3f7abbd00819e559d1e92553482df886e2aa21adc0683eaefe435a5d675ab0556b576b0f69f34f036516b148a886f7275e230109ade970e72f676d687622784b2a4c090f1e608218bf9cc26ff98087cd4023c62c9233f1f209445e94bd0acbb45473995e915374cd771225d1cb4ddfacc87be8fdfd31dc2f719bf7da6420bfab223c25ffe82f8ba6ed2137d667d8d358f4702b98a331c873a4f83cd0d3c749932fcf286262ccbdcff65d7be077ed80997b4430b62aab867787ace7e60ad55a6a03940a8abb6c89e20c2651c842652a4ee16036582da828a1a9aa0d082a09029381b5e16fba49a5d8d13396e6b9305e6f2992a7c091b05b99c6f6fb13d06a96dfafef6abb09d2c9e5ac1a8f9f1d810386a223eea164ef16fb5248bb23aa0796698f0d184284697387c798e01b8cd277f0b1123cfcf44e02c3725f538c5e394a37eca20f29a3ee9fdf6be239aed3ac3b122b3108042420576f8bf9453be9ec5cbc673f23976a4622537d275f8519d17f7840297de9ca11807f57c0061680e81998b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h96c28e732e8d6c13757c189b3ddbafd9ed2d31a95bd4f5392948942d997dcafd5bdae464e82d6c03bd40c3e2a4d901dba5e255e4a14569690d2786dd5031ed7d28daff48aa7805efbb24907bf910c7b86a86071b74abb77212fe84b6788162e291125f776962b106e49ad5155070e2aab89ff5b8289eebe81293b4c1eb158d2284b6e1d3491737087697e2d0ab8213335071e80fcc0bb762d30cb34d953c4dc93164c41b5e4fb674f2870e85567bfa810ab61e7d4587bb2bb28e1fa3148c9639fbfc61898b3869c80a7bf38c603ecb401aa2a0e7397dfafd2a1759d3185a3c27d4f2834a6ef6d2d18b3de3279e8309b250d6824eafdccb903b7617a230b5cb6eeab198a8eea80ebae6aa096a13d7e0998d7c5cc2ec65c68240b2a3c45224633f3b32cee0f3b26e7692a02e5f690c60b30402ff282194992a0939c58609cf66e86c5c5205297b69c311be831c5dd5594cc15ceec221a10f2f13edd2ed285934eae93ac9ada8c7a5f03d17ec93c4c37c95a8d00b76ef287796491dbe7f00380b68671dc025b0dfb249ea06dc521908cf2f657d96faaca8bdcccf718eedd6c151fcb9361318b32b484fabfa65400dd38bc60fc207211461ad189ac2da512bf2ce5ddfe417fd1c4623dea177110e0e7f9e17b01f5d5735c494507dc4156e24f0e08c07bd2ac0afb658fb8f036390936cb1d1a232bf6aacc4d6b038e0b7231b05ca6fb50541c5ef1b011f40fa404d157ddf97ba952dddfa858078d407127b1cac34d519ea19b06462b0fa38c26abe5c3fa08d40b35ed5c2347973d348488be855a8843072d15bd3e37bd7376dea32b22073e5d9eb2036de9812d24d617b35456d535d92d52ac3c463b33992340980144796c048ad949f27fd0758005f090ea09176934f2ef70e0b3ca9f38f13208dae75e69be1a2da7507cbc6ea3f40ad99609322167acb49f04ddb3c42fe13bd6954c013ea5f25814acb040ff0def08b263a271551f9e7c789cc6fc4b4e60603c8e08ea751e10818c6f2b532e9e96d0ad598e1ff475bff51f40e311b885e1c39a00b19a78bec9f115c8743faa603b8cbfe5ebca167c0185d0d2c9ad71fd823218f7be12aa2afa09cc0b00c3a39514347b5278bee4847aeaeb9549a6e2179df3da6b030629b11d8da32535a631fd34d3e62fc2bd78a6eaea0d0ce7ec681c99f57863cb7ff0acd1e5d69f10594b92439bc472ea6a435a785c6223160e8773d01654e26aee2af5333cd99b725721b3954935bae3997abce115682ede98988172eaa49229153ecf4c8432ea30f6619fbd7158cb23d8fd77f3b02804d0d5ab9e4289ac801de1ea467afbd776fab5a4984372c260edb1aa950389b130053805bc75cf34610ce6fc1b54149477fb2fb5ad9b2c76ab410738e2d550bf4027c02ec4b18e1260248a466d747b9b41794d7196e96b9da72857e38f52ba5eb35c5027f1efe1790e9de8719b95148cd283463efa8192c23f04206bb08933e07de0d4b7fc111d49d84788c28bdb53dc645b264c8b1fab494fe8b251f816f494844c0f74e334f36dc9a2021f88ed37fbcc908b8a52948ef80c1f88898efb544d008ecbb94527960cf0fa1fc7977964fc3e73d38f373165715ae94538641039fb68eda2843677f6b34c253ae394aecbeb87232e7f6f678e5fa87bcf3846c349e1e591f2a77dff6ec45dcb274309d1aa6393cf2ad2fbf874fbc29db83aa54762d6151e1d350030e9ecea4d1af4849818afb8debc8c4df501e323d6635c12bebd262c2e55fc192eb4eb47ec1c5b27fd327583287b95259d0e5cd14f995f1e0f110036791dcea116c530a5b506f5ea21f16759798e732e4c4b00a6fa572bfeeb7367a930fa060837b0eab4bd5b2b022d7ca24a814f81bc761d248808a4ef651fb22e9549ceef75e201ec9b7da5d75eec41a2d7b2c42107286a7dd44e49eaa604561c0357ad8c5bc4b9d4b4c463f14048d0a97e71df261dc498dad6f3c1d3cb18743c4d761548e8b6f65d14a1fee9a031a18eac674a827cbd133edc875735b12e442d343dfc4d9800f8c226adb18448242dd1f6c36e05123dd7d47b139b57d15696db60cb6d3e700677f7928489f228406f9eaca0db77084451caa98d42e9e3369e47a242f08a9407a10b6ec6cd0b96aa528ffd22ac472a2193a4d34aa49e04f76fc529fe4565a940844a13dc75bb7adfc1daa030d75c4d31d8af73eca2736d0dd6cc290d2e52d1e12ed121c7dff2dd781cb4641e0ff0cb47fe4e69654fd9070209ca007a62381833212f45d09e100df15dc9848ab234f1f54845bb1e27289b6fc1043d745e7c1d75f394e4346359ef33fedbfc0f74e1f0330294a16b096bde34bf2cdfe4657b241ee3f1a39c00d039450f21f479006897d01d3a01da0a826df843009a9a501a6ebb3f8080ef7104e261234f58e3cf59c83b8e9274f31517f935f008fb1985c117290c732f2d0d9b9f1de0b76e3ec677885f4f3b62834eb9144b66fffb467a0851a12f9a5cadbcb23036a546f9a0476ced5345665c754b6a0ced8eef91779f593fbe892e04f20e5881839c6404abdd31a8e8028914fa0b806f640e99afac08eb6e84c26b1083a2e5c55ca23269816e343b7004d28342e51f80d1cdbcc1c617171ab5888b383900d813889348e03ab2d63fdff596fe0ad286773ab721217a779ab7b51370d55b67c86a120321c5afe8d3f09f369f9eaa87d28aeee2eee644c2119dd3d9ccdd8b5bac8cfab88aee93d8b33d7d8c4f76016774f89634d39e32f8dcc8a5b675bf24ebd50a01df43e6ae0e02a545d1c4c730c166395fe01d37f3a772dd5fca29e3ba44b42e93c3891f5f65d5c957656b47dfe271b1141ef87702f43cb7a1b975b935240681bda2434d7e6de6563c4af21d59e7b50d957a9aa0204e438ef841e6c3ed4af4f0ca67d9c8668ce5bc56465675662e95abcd0dbfb73990207e06c595f22edba426704910bc93f749c89eab2393e5ef2a50a40f8931ea4524a2d81cafb6754514e6d794ba94157be04ee6b79b37c12c50484d6f3c5f0c9dfd12cc75b2ff41aee777e1ee942408c557ece0b3b6f4e582b18db0984273764ba11b900a7e5d6de13f5353c13cb5971202859cc4dc1c3efd53e72f49e6c4300dbb53266b8d27f568de2c0ceb93af4e554921920bae0e9adc8e4bfeaafdc1ad0262d34f67212ff2f11273a07749784240750847dc8fa65310ad651e197bdf24e71e0e9932a3d150a116578ff6095ca04de59253dd5464c06416392270a79789c2e93c972fb567f8a288b7eeaee1473b3a511a72d03c86dced2d51a4e12015386f4457b66829127fee5ed3ef56d87aaa9fc00a3bdfd2f8d8d63edd6d8666d520bd4e529022b8c341ae28c1d8bca44646ed4c6840c52e1675d874e432a6fb49c6b8d8424928cc4dfeae2a2c43d2bfc69cedaa297a47c61de31b66d879182e573132d7b4de670b41899c35bf21d5624ec1e9087a50d3ebca4b06832f87eaaa73955ccac2b57ed7642aaa3b570753394a2bab1de63c1690178fe973acd71cb17aa5fc53945fcb741f9e8b41d994e3a447df8d267791983957cbd062ce5922f5fc8d49a8504ba88237c63b48c0bd85caf1dd53451fffaa83e8a2197111070f0d0b12c98c2acbda349919bf1941ba64908020b7ef7e9d265a2399491f89217b2e0f54168ddc9f3b1fdabb039f32114901837f0fbb8aa58ce15044309230ccc549b8dc11d5ef1a7d296a32f1d3a7e64cf8da4c6ce474ac1d10e4ebbca557d3e52c48b6e2ddbf601c0798fe2c622490d4df1fb608db68a37e12670aaaea7392b49c49356a23f8e14573ea03c3c5da0f84792c8acfd4b39a5913bb8c3bd6ca79f5573b0e61e829dab4d7cd04ad3305e4ad9b0bce1e3befdbdfcbe4d9b20a6b3bcee5b646f34ee58266698f000f6fffdce46e258f4b29ebe8f7dbfc5b6641eefd1fd3e3a72dcc6b26d535388863d488437c06bf9f0df3d61061c7e1b51f2897e30889391f5d7752be09ec7322a2e028be8a5d6379876a8ae22706c0846305258c1916b47537f0c8f0f47fb6158115f57143e82dc9db4d9796e15b47f0054826d5ab15db46d8506fe6d8ea536b0d0597d18fbb64129927dcf5f7db6d8747f2e25cd555b55d98eb738a1997ff020690216e32b1770cfc04205a17a294dbeb161ae82f206dd291749b831f076f71183c36273297c6bde46ec06badffd3dbc2bba880471c493d8a2889dee4911ee9d880c29206d13a08f51386c95ac6de64e62335be222120f91d9760dd9e5d4e6ce874e6431db6a9dd1915daf6a2cf65b2a143b9ec866e9d218bab0fe20eaff904f4187003f333836fc248a5e91bdc77de67c16d89fd92ed14989f4004f742d901f19da1cb74c857195e7e84cd75ffb96173e2da2c8d8ce90a9eec06be3024d7c01e1fcd26bdecae1587322dcf13a869f96a7f07bee2f3aa5568f484315a7bab0fac39e945210dd75448b702e030ac8e719172667b728c9d81ef435a3e915bcf643418feeb1591f61bbd78a19edd629887dece959b2dd097e4621c9abeceb82d7875b1851fecb0f377f52e3c89c18f838e5e9a2724dfefacc06128a167e349b44966ae2908ceff11c1ff261207912cdd57ff23d7c21587fdd38dc1b58ff5d4bdb52641884e5b30f42e2ca6d3b5a0ecb3f577716e616c76915a12cec4efc2410ab05602f3f3dda7f9d6f73c407a3165601bace03966859b760636d4e13baa9360543acb5fb8adba53aeb4d037d53e4bc6fba65c3b5dcb550b7ea98f9636920033bca92335c770b27360b771753cbec9f1ac601af11cc598add673ba5a9be731c2787500579dffb56d80698ece0d9bdc257d90c5cc9b46731beff01a494b10149fb1a468af66327c80969d54c578e7a850d8a5c816e470d572a97cc953c939572dcd56711b48a102c3d883678ce240eaef7a8a5ff379dfd3ba1fc98bfd0b35bced1faa3a3e03dbe5d43c2b68832ff0589ed8f3079c3e712ec8565b07e1dd674ab905c64b146cf7c278bb8053840b3eff30c8f98e374767e84a378df486d44d998c1fc8be89e73ee9f6fda117657f757c4b809ace017dd6cb71b7c98028804d2b26972ba8439a2fc8920ad6e8e0d68daadc8b967bed6a1eaf33ae7782313fd36ef3a63c4a9e3134642067ad5dedd3a261254312007922bed985025045d8cbda509ad6ba84a3940203a02f0ef249ee889f765c89c27065d92e2f3ee8ebf53880ace9ec775387983dd53309bbe496d7648d3fd51de89cafb46009f8e1fdad5a16cc2c1e8ae4c2ab3512310a311226d304cc1322e7259447b1b646e2896adf01bf2d8e3a379bfdcfd488111bc7d8d4d1b288105c6e48bd5450845ff9a5cacabe3351a36946b59aebf49374096deb9e61f1abdde97e8e4c39881338276752136625dc38fca59ceb357d337daef39a97f8124050e91ab4117c2a7ee9430633c774d4d9e833f25516d26dce7789c1a2a22429e1722a821c7d01cb0f7ddede86a6bdbf26fefe3394761b4e353abc2d6f54cf2965c65b10366881bfbf648b8ffd34988c74d88f70ba81e2d355a3543f72a588ac5aceebe74cd6a7166b4e6f2c72b0dcb9f974ecc8ba27e882e3efcbc641384892bdc48061dded3d5843e794821ba9dbf384a46178c7223f3f4676e6ef743bb47ffc62cd9eb549443a12015021fa1ceef7d6e542c227690bafa5da0d37dcfbfc981ef65ecbe9f64154c973baf39adf1ff609fa7628dcfd4eeaed7e2cfebb369ed27b4c6910c70827b6dbe80c5466f744c2e0762efb76f63a88d1577a682c6781d3ae33c0e511c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7524d0d4be0b0e18e5f75ceebead053f7687eecffd70d3f06e6134358528a41e125dbe69f068a7818710607ef6ce2b3e789b121129034411e6ff7e7aa83c1f54cce7059d718346d028c8d941ba431f0d8707b8bd0bea398bb212acdd1794d0d491d9f06b3051e7721b958adc3c5667445315c875275f1f755bdd79d7f344b1c67d3e4ba69f0483201c1e3ddff01e8450d2bf0b7361497c50c7bd3457b85a0c4a3a8c1ff2be7e71ea73b39c2336e20117e6ece90c75ec9c8326150f1e5c7febc9b3f54120fc53565e5597de9195c462431be820df641d3cb0dd189abf9f3ed7838e168617b1d18e2115370b501abdd852da78411ee6d654d2862b605362a4c51d3f5bd929f5b307cdae511d90f67c2a03cda367a1615ca3f14dafea385ec13a526aeeb790b2cbc9f47a497b4519efffb84a5ada8c94f86ad756060060d3df92c9c4d987fe535e7a78f6f18207b23455dba36d36a549f537462bd4796dbec928e8e3d89e32640ec5856fa7b95aba29724f411583dc6e54b7fb5886ccdc727af9594ff52e0e8d3a0bda8547f63d7146c636116583f31ef67fc7149b50ee035643aaa1f0950e345768f9caa608342d54e24396b1d148ae5e474c1c5e03613f1163f0abdd3a993e3c48d40c6aa50dbd10c617af3f3cde65f178a803b8d822896d949a47f1b6e64b7aa8f248f079cde5a7803c45af8aabb6566f7b08f0cf3ce16222983c4b94c180f66cafdf1998f5152ba32be1ee40be0336eebe68c28dd843ad65be080ac18bd12f87cec5d164d2c3750156dcad076341367b78b0b95521066bc775562a4d7c356abde7e34f43f042a0567ea7ddaf2fe6d13a38a708af4c90798acbaa356e9c73fad9474f8389aed65ae5a6bc8c3d2a707d48e069d009fa7ea5e0b56897ca63f2cd972461bc87d293bc3f25494d45859523a0df2f18afbb0fe66984fce0601b9a2a6a866da778cc101ec44fd5adfffb9f0a30cda91f28dada40b1e6cd583f7710157b2d26807205de0333346f03956e52157d433b31654c376bdf7fb73f9436850d1c1c6a39e4409c7ee36c07a6f90c7244c63b0ab7f6a9d7fc47f62d6945ae627e3174f50566c0c62b68666a7897876729def9375364c877c7ea8119f3595bf8664c07eb93feaaa2f4af01921ff647db557cbd49fbae803c9122f81b17fe40cff3f6225d3ae9e2522fdbdfedda90e49eb3026fc86e9c29903cbc7b71efb242114dcb33433f4bab3f7176bfcd29756ab1f960d8a5f5f9135635d131ae2381f28b991ff10969588e860f7c6541a0f850d90dc23a8150505b6adaf5e3f288ad6303da7f45e793d29093665b07639dd5e25f334d93ccba9cbf1eaacc979cabd8728e5ed105839ca79178e03e094f9217394cd9c360626b8315596b0146dd9be9bb3545b3dbc9f067fdf6bbdf0816f470cd6e10960c38886e260635f117e08034fd84cfea9ca27f523d669b84ad20881ca67f4f0d977ce06882986dabad9793e07f99289a2c1f60f30a01c97f0d534e6d3641be27daa578ca4410862c07046aaceb2b6f7942989204b20aa9204922857e8bdbf586570815fe6730a507d9faa765e11dd6a0d4c5902e4c411f485070da615dcfd5796973a7a930130183e4fa84efc708236db36bc972c695ad476f36efd648bb60252e8a9381686c329ccd694de648f04bce690d113358afb1e87a61249358827809eb573ee79c826af266307ee62833f17ef2a222e4c8cbe9798f35e13d49fe7609a61e181d8209161b17b2c83448f25315da0228cdfc24ecba328847d60c4292ee2dcc4f156163ba7e8851d9b4078351291bb12aa5e55834e1562cbb4802f0e2c9aa1819ec662b497d22a60d9ccd81625ae9897f105f5295143445210ac7b099856b3b094982050e15fef1c7a1efc9caffa746ccbf9f636716d09b910c264cd90ed81f4b74b566ba141a31ca58e94dc82b6a48045d2a9b0eb9504f8b5cad000a255ae84f5991579ca02370660b0adc74fe653d99ef59a782f1f602660d0d759bb67db740ddd7a385a884255ad651087b06932c0f9819f91cccbadfe286c1ffc89d5f1c089ba361f7f6b8201863dae5f9a37cd4dc57cbf9bbd76a1ac1b2e42baab867f5b0e05ceb26f1576ea25c8faea78df9f126ef9580a53a97adc498f30d6a1499be3b008ad034b8c6660bfa89ca96ca965f07716ee76e1abfa0a08f7c585ab6b6cda244c0ef1b3ec6dd918f61bd76d5f49217fea54da967dd1bd7ce33e13fd8f239d6ab861aebbfc3ec77df2650c277828e53ba778550a332cf3146f5c13e2490de1bad44c593384d23c03210621b61dcc6e732fa4ec88f1cdcbbe3283d6f51b833530457ecb88a34e7bf28221280ee9898f51a4cdeb739e4bdc59bf69656cb461d328196a4ad1f6c3d60e85356c2b22a460945f7015df43e908a25125717da8b5b770fb34b312eb5c65b6a6a76033a40ec81c0f0af1256e048394539a5d656008b5d703c8d50d1561b655349298419c5a31a130345c82d00a8714cf3fd238b273883debb4db68f31ef61880de7397ea324b0b3ea390157027e473eca279104c78aa86917a853e3f26de748386f8949796fb2ae541928c932a57a704f54ec51fdcdb991e4c50542e0a010f452e499017e3e90fa0fda672bca37975d5d7daae081024ea03cfbdc7ee0b85be406a1a3adcb74e54909b834b37984fe07da98eef05f061a9d2b3e45f7225cce58fce1c4e52b1f1c6781db92b07897a1d41377ba86371d03f7d760d6a2c1659a846d5f2960765567a43d3281f5a1558fee492a2a3752b62f373d6b5877a4954252f361c46bed8dc0067838290775a76a212b814f591386f81b4b112cb570301300961aadfcd0dbb0a946e678574a676e64a61b011526b085ef3ca38c46a27e4dfc68a94392d708b9e2f309f3ed0ae3788efdd2733935a30085cd78842f05051735e81b4add18a8e4481501234bce04ac008b153c866f1b0a48d32b2fc53b0d3c83e3f7f0fe1f647b9931866f4a8e460bdf32aab23546ea01c44a41f00d02ab91af827071d232c1231868b27e4492e20aa6838a82cb186cccc350da19006703a1c3f409cfab204a48f37df0e7ee1146f34731d0eefcd15043d892c6fff32fc7dd05a3a5bc4b0e78950032275072993bfeda764ad206c519a43802a0d36bb928b85e6675c83683c639d30c66961d7c263b5bc2b2225a68e961dec3a570aec8fd5c72433943a48b92c2800285750f228e51d9d0fa818376c660159f2d0993cd4ea86886ab3399f2b721d3184aa701bd8955860eeb6c0f226813596fead9a20f0f864c1a352f2df19dfdf62889a57f531f1c1b03f69caf4a841d09c49fe4ae8b4a2993455da0f6ca57173ac2c874f3ccd8886236e211fd289f377790d45ebda3588f55f03ce14912b504dec9e6a1957e4f6115b32b64a4a1fb33701006834c1295761aa676899a1d6dc3b416269c64adb9dc809afc1f407ffebbefdf65f5d8176c60eba22996e03ae588230addeb1a0080b6944545ed6a52510464439c99fc5199051784081ca841e5c3f4d4ca87d2456958090dcb788863e8f5a5ef81638a99db17626b27613c8064621033c439b51a93fdcf6c03a5b9c6a74a871a777d4267815d169e2915ce9d35234bedbc8d53e3e52c39819eaf6a9f7a2eccf8d78900067dea5245e69a0bc4496cd370ad9d3aa15730da32179f47f9916499a1ff494e97034ee28b0379aaf53965f8838e9b2df3c7596b65c71598793d884becfca0c9f530e3b08af8712ae8a176a5245a35f6afa9b4fbfe21d2e0f1b238b39cd9a292958d0f1e1109aaae57aec30d10df995edea0deaec92937256fb78ef0b909e7f8733e1d8b7abf50a7575604e348498353a96cf6812c91361a086ffff07eea4728e6a3cbb8d7f604b4e446ab290afa6f908bb91dfbafd163691b70fadd438306c43a4f381c6094741e59f0a2bb896dd5afaaaed0d99a45e3d6b56984b41ca089ea5835242af4720f8f025d6a83fe7f195a0c452948db4b5c757bfedf836e92472599f47c77a8ca30b0f8d789909fd342c73d9737c561031af7302ac8bae3606846d8a66e466aad249434860cc20c6927a07c7ce3b5d1ee5a9c64640b63efdc9a4cf393ad583e09c896c1243a6430c8932b96ee647b008abb9269d440ca33eca2e4676015b924343c60ee5b1071bf8a3d55d6f27bfe13f4664f23fc0a45c528e51138f3b25639172cb1992ef48e00a952765cbef8fd448fe7301a27bee483bee58aa126228905d71c1597fe2792d7d3b7652c784f6f693844aac83eef08a4f65c2f7ff061e2730c9966303c261ccf4c8ac4aac48059f24aca3e3ac17e88eb25e6fb0fde6934da796244173173d9113707b6df109bc563df30acf133a11ce96aba8c71e1310ca82a0b1819e55094aea690b5b2f22ec0f144c69c587c871fc62f91cfa02eab323f8324c7f39dadfebcb9ee59d7ecf5b18bf498508e680fa338af158f7fe55699d2117d1aee588d85c7a030a6ded18be20a1d546e8ab5f201d75f87c86ff42fdb3ac44695e53f3741a0dc505888d5a8b1a743bd8cc996fc0760bdafd55751911fd660e6927015a80f995fa2ff166f656e96813624b491eda3194b60aaa2a8d81b7cd6266ebf82c2cfcf87950dd89f493c308d753cd0af2dec409a84592ee6f6f560f1182a46a7a6a55e98a5c25b4cbbc39442587ff9909ee3ad65cf33b0bd196315ffb2064d0f2f03349da3675bd6f9650bbee3c615ea1a2f769426a90d7b6025d59d9372724199bb171284ab4ae23056f87af8d0abd570b3299469fbeb5be46661ee26e7e66d638ffd992fdc65e91a2fa41692d00d3ebbb0e6492ff52a2466e6dc8e6ead6da60ca03899f29827bf28c9cbc178355e3fe58347e2c014345bfd782a4e679831b043b7ad0fd64061d446439d1198103ef750938c44d2bfe71d0ebf0f8efd4575371f1943df120c510ac8262f2b44497e4ba888c0ba52988496fc01966d8241041108477a02992cc775c6ab7dc73750d2e785f15617b98548bee18a33cddbab626bc3fb716dfa21d1aeaab986d63b9682bb961eb93a0aae0cab81d72349e877d68c07623e0c707f2d4f023022670fefe260c60996ee31ab262b2d677379cfae7d7c7b238bb9f222a98e74f1c1bec26f8db7d89b04ff7d30ec81fb0bcf5b9cc4dd848336b3186580b7a6548c23b580dfed27e2c8b0c692240cf73181fbadd0161f4df10b729782cd2296252fba97acf60ad657a0a1ec311b481438a56142c87e74583b46f10ec892adf494e10d462ef0cca458397314de97d9d0eef237d2d9d4391799daa0ca062ceb97c24fdaed72e70d738a7962b49010963402f105a5486ad8a9b567cc3ad5b5cd226d4996303cfe1e844a915d427d0f18dd0153304aaeafc840fff4d8d601e4976d4003499ac1adc15295435a7061ed176a2b3c39b33636467d883b5553a51c459da31f0e90fa4cd4e783696d12e972e086889e0952b78857cabdd587b71142c523a7a79370e50541422a96a21f548cdbe6e440fff91a34d94a18be6f84b7a2773bb844bc9143bcab6da28b0c96c4fb595fb58ded15e475974c5d9d6bf115e4c0c3e014bdd4412f052cc34a35b0d292bcfcf5b19060bf060e3db5a4df6cbde1fc7a92c58a0efd2f0a292668e4bff7899e0ed49bd04247284b602ad2cec75c9ea41ae30d5a1edb6dc07e5271cee85cc40617de724bfb453d6cc40b46280e27966771cdc5d553af5c05a8d91ff5716fcda57714c14747eeb97b96ce1dd9901c3265c08e89416f40353be64fea3ac4cd001f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6fb7f2a92a4cbcc47508a27cb33553646d310b7232f9db8a621697d0878642ce80d8fd15cdfc59af4e096be9f34803b38175e71b85abdaf452ed7807c44c13d1db98ea8ad608a3f674d7924d2141cd56cec5db70aa16e36391b86449d42494ddafd04dc92a183afc46b72f68a08b7f57831c3d5c98d341eba1aec59d6ddcab0df4b1e58efd9a2f27c3f1af2a80fb3eba09ced085cccb6215e50b8aa2629fd41cae722826aca899ca92435417bfce6acdfc62db3e8e8fd0336a9f6d607a3ba49ba1f6f25893d2ddb6c8dfb3640391246195b6cb7fac5b92a3dc12ef862fac19e5cf73ef2672b8d9a87bc0d51844c5b677c3be35512d74c37d5036fdc732d21e9227386f921dc6fa805cf0539c4435b562c00fe64b67d01ff2d384394c57bdf108a5e8d0c0fcd170fbc84447a00c297e944947afbf463b2eacf49409a1ea3e5be64b83fd461bb0625baf2f085973f0858ff708357633551de314861d0aa53b2615f4f0d7823a671c5954e86b61ee9c7e353b05f8cb3aa2c48a3105cb1dff12d46d4f4625ae54cf60e97931e14a5783fab397ac39a4fcd7010373b797d6de83aa646f26fb4ddbdb8b488169327e8a14775a8845c090d7eaa120eeaa119dbbe2846ed788926957f4a5ac4f0372a251aeaf45d2f6023e22fb9d4db226c590e829fe7d63249a3fe745f79525d3a8ab571c69cbc0a1ce99a3ed34ee84ab7be55d1156b6fcb974bf15f0a4f18a87f3c174058c531ba3e586daf2213f299bc7610519d3ccca9fd3e32b1426a2491291f6178546c81d8a65aa5a61f2f5ae13241d37e659fc0e0605d95bc5ebb1160f7b3a95ec36276ba9b55abf6845d2e8c87bf689a103e1abfd117ec021cdb67da14a92dc7206e6810cf65226fee4c90948586d668af692b3c237a3fda33213ff2fe8c7a03dc543c7e95dacb1c5d969c2ba09d5b521b0dc8c743c390127b652e712233b1c90720816963fffe4ea7aabaa53b4be7e930681b0dcf9e327475075b987559f3e5480547a99efab2d21d577bc2f948e4e215aac01f527a440e0d44c07f037dd3f471815dd660ccc529fe0e932e6ac3e42c725a80895abd2357d1be60f94655c7db3b2011be87f73ee02af677d8a3e847e0b081909e4149a889314ebaa9253e5613f3b127422509d537862a0907e08de2599af1e40953aa607c2f61c4204a41b2a16358a183aca1029912c8c696fd3676ea7e3688186a7dd6154e043514ce38eba3663360dc7788d21f2c48f303c69dd6a5e3eb7303d014781a6a4de7310a9a004407ab38bb22e40256a3aa2b2af10a38884970c550b2b2558312745ba24b4ef60f8eef7d498da20c12e2b17028cf272edcf0c8fb22aa445f772fe37842717e5a2aca1ec94b1f690c7f53b49aef6ac219be996499aeb5ed56e3245439f546f5b42c38a756eff07b3a14f80a4623900ae6aaecb6f56fa6c2f6281ada02fd8fe5a1aff7c13c414e6071467fad060c5e661ed76521556fb7024ba0c989d7de2857d6762eff9830f1238b51f7583ac2d14790e5a755a30137d9c8c66e4de95f959d49a15ca5d25e1ae42b4c134cc2fc58e6164467004be87c6bab204bd4155ed4a373719be4022a73740d9d1517802fc1284c7f4c50abde1e74f5f0e20ad2a7c92b717a5b34d58d73b3022e39ee9d237d646a47607dab91726129fe9710d9debc7abee1769cdb9913214ef638a566963ee85ef30ef70f362eefc62ba2ed6dee76cb857372b56e78898c0e0663eebeead0d7ab10d26f15f357177ba6d8148ffb2b78828cdd21700a3a4dc15f8e83ed1d40004a9b1f427f6ce705853be12951729cb378495a2debd4e0cee8486c6c6f4d1551f615acf651834139fb1c72372b0e1e3c217486687d4d45d14e07c98256d738800b1ac106a587056dc160d219492eeb0012e0ccd02c9255c1f83a01ff6a3317240e1ac6d7f2137576faa0916e436fac5f1675e42fa2d695a36768ed233514f28dd001e237173a708f72d559309d90762b4daab1c95bf99bc277a2d8543156e207374fd258518cc4faefcead9259318c373d61a8765d3b3f0b55c38365f74e924f8425a60bb93048ec4877579e66a9b1467af999d4ef0e38408e02a52040a83870336ac95cd9ed8c00196646fc50b8717c7327a512881d290712ae56a5d60243d6cb3acacd69d8c98f745fb880f7a072bde120668389a05da3109f75dc7f6442247e3706c28a7013dd90483320cd0842daf74333e3e9b2d60ba381ef97126a100ecda0c96f4c16621e191007444463d83f191df3ee1b2aeb2be9ae64fded11ee19f35f9ac8011f7e28cd6f476a61d67bf41205960d5d56ece8bcf94cca879df7634f8c8d17d67a49ff5f6258facc69e56a4a24742efb9473ad86d0c5a7b26e330388b44d9ca3eddedadc42994865b2af9fa1ae290b57d17bb847006e7342d4e92b43eadde403d1c5e395fc2b109ca6bf1d3d02a69c7d222ed53e996ab2a7315063f786ea6d93a4afa528252fd629c56ee35118716bea4c18fff4efcd8d8754fb75e8444ad552d1101467e2e69e7f3046c7964c046827aa020aa09a026e6b455cd9c92a8684bbe9bb85352298d106c9a867d9031bd699f8cbfcfc91227c83c4ce3a3c767862ad4ec3b08294fc42bdc6bf8d90ea11a0f2263e237aeeaba190bfc8b24a5251954d8425dce9248c7a6ba0238e57995745e328446aa46c82738b6656755088b80d29214132ac7255d86e18344f4ad72c32797dd2a4c5837f6863b16214c9d633a5186b18ef180ee644cfc679e2443c6459aea636f1a499354537860c3d70cbc3a6894ea6e345b6274e9ef8aaa39d84ffab7e6c8086ea44a1817daa7e3414e53debd191a57f883f6ad24b1c412088a1dde3a3c1d0a5413a80a6e9b37971d077b2124c4632f453f41a5a09752534621c4c936a75cd438c5ef27c326dc24a80269c674b8768b74306b89657e34cbef00439e1bfc1c3f6231ca8900dfaad4497f90767583a761c114aa4b3fd625e2901805636dc5cd6df6e9cbeeb66f0473b7464bc43cda2e22a69b96c89600f84fed30e4e1b2aede7985cbf2a6c2be35ded47a491037a02348e3ccc83c33dd19ca1fbaae8f307a0a6175da3936494a4895c235c8bc99894a11846cd59e5a01a09f74fdc4f8e803f86fd709bd1b29e26267782a191744c03ee89eb9c302b589421c5dfa30bc32fba68393b39fdb56ad6a27a217a1712003df279ae33fe82b71b75bbbbb821198dd6b134cb4f0e3fb53218aa1dc93a5992dd73e8e6b586a38ee57c822bbd1b5428afe075030e4ca7157cf017d1fbf3e8220f5aec8cfefb0046312caf4179a33ae849102c27550145fdeacaa401e8ed7e57ae9729c311fe26b02512df26e308d6e4f83a3e639f1f5172e5bebe85ba2830d56d4c5d43c8b50c0266755e01986f7d61bdb32de7d01de7169880c60511a93190ad266a9f88c519d5558bd9a8c76b63150938bb4bdc5aca1e5017d2761c3c42e54597aec420a0b81320bdcf8eebf963cd8374802c86f045a76ab7fef41ca352e700312f64d93c869ab13ef142d7ab1eaa0472936e5275df00db938fc053ebc1add8fee4e5aac6344abdd011688ec1a5cbc457ba0ab89a74c3a2b6f448d1541814ecd33b1864de20bf3c740d691fd8588fef036bd295cdf061928ed6c854f20a3231f41387450606341b05fc696ff66800258768b54eb3544e1b9025071e352e5163c2b9b42c24b0faefa59843ce8a1d42e885b59fa44cfecc8a025d50b9bf2519366dc7d2dfdfb6b380dd109953fea1a716510c8d49355a5fca8eac644d9665e536ed02be9f320a394ae959328778792784176de5dc9a464fa33851b7cecb9c3188198fe21b0d2b7dfcba408d88e7e23cd0fc3ff6ad264ef1ae47bb616803fc2f3c40e0a6d50ac246c5036ddfe4dc50cfe1af2242084e414134d5d2d55ddb09333e9f39722953b5a8547f0564c7bf0a964c5c13dc810cf7dfc9e237645426939fae5a41297b60facfacdc3f700bf65300ab8653706ff964fdd2ee1a7c6e3ad1ecbed6e12f3ef81cd45c5f2256f7fe94e1c5141074f92d0bbf10226e8c474b9062323249468ee4a78ecfd4dcf4da1fd11ae11bfdfae1e7865c76dcc35f64d6bb02a95ba1a744563ac42fefd2b84607f0b2e98da00525a28d662972fee7e76d789eb750552aef98c5581aa223def16ef6a0749c5f166622bf4b8096d613d9c8443ac013dd16c400c8ec6b432a9b1a9d4654f4a88c4dc3fa129ff5df5caad5a428b67ae357305ef5f38fa5a4ff026ed6e131536a37127ce47c3f40f8fef853fc6935971fca10b404784d736ab9a87d7062cb3d2d824a76d478c61fa6d77bc5fbe76fabfa7ddd06b4d6722555eea443caca36cbb3bd13fe3e35a1301250cdff848118f9be08311b27450679148c9f708b99a25e64e3cb929e257c9320e00144563d6d8b39e3b02a3a345f4cd420717a7b53fc139734ce2f0ff12ef11297140e87a97073b8b1ab6a1ff3bebfdc93c6df986249fd42a26501ac1c81a93cb93c401ed842247b6727df9405f08582fa52df5ba880082bbbca37e2071b056957e4a1296b0f1cf80283295f6fc12d6f8bb94475624f85488b1f394bb20324bd1b575cef07230835bd2e773144c0c7943c4640b8e2696e1d2d0f15d5e027eedc56ce9a4b2a6f447138c91ce3388e4cdf6c6a7e208175a4b3b8135c2421397f73d8c37e3ca77cc66dcf6d7902fcfb3a21683146757b294fba96e28d78ab2d4423753f085f5e712f2e08fc0ad904cde7229e36a882ec138a49159efddc5984a2b00a9fda4609dcc0a147b842fe85ef2c24376501f3e0f5c1bd61c067bd8bac3e9710581436c54cccb80f88fc0b5374303bea0166ec571f0f99e726a9929e730f74743c0ac19692d4219d8b9c6c87d3a4bf4b9ef89dd213bb7c5ab35b30fae8916de7b505b032c4d38fa47214cf45b97c10ce2b6e1e84051ff72cf1f756710bd9846d52e0fc25759e03b9c3348851d32f164e5d0612b0e730b4ef93e02bbdd4f54112c9fca37916df344447642f466532aa916527abb67bd03a14694185c01205755ba6a9158dc0aa7751e67bca9b19da3069a9231003855e4c77cb51d9747b9eb8b309062ad548cf5199af32134cadd4e617e326ea1bd45d432562395b3f2477a9707b15a4e375c92e0b4bad4c086dcda58533e93b3f382f11d5e286b16e02835dec6c4e14580b14b706570e4f4fedf853f373da685ab2c0c2b5c8418ff85f5ba1b24eb407fd24712bdbfee3a0617c9fef6a538090c094f0e6dfc16827576ac8923f33884cad1b693b7e7ddca55c6630cb3b83b758b7fe53d09192a480c72e2950f131ca5af4861d4e2ee3d8cca859130061aac5f5dbb4dea698a922dbe03246a324438d84233c8f7bbfba4a13c50f6f075d6c93cba8955cdac36b5994bd55f6778d24d388ea1ac3c934708fb2c3bc4015cf2cce1ff1778dbbec3a20154d17264fb9cb904b47478d45e5464bbffaccf1c9add4165c6fb68aa666e773ae50ecd43d353d802e243d9e17e1ee25b24ec88db0d47a861d7c161afb883b7b533c265e1466c2e08a5285b6fe429291c0e28130452504cb0a012ab2443a6dee772e4fedc4e21433969135bf61c9475bf5cba70250037d9263c623403925f9276320c63aa68c790f808bf821aacef30db379953a43300b8ea1a8ec7e6418a9c9ee91067ff5a8fcf6fbd392a046643b488282f8487c98e12b2af700d6c235a46bf2a97680afa0de043c185da596cc39d6c3344e4552be8f2d530fc63ac08f80e0e0d02eed8d3f878f223b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he2f6a2a9da2aef455e3521a2e6098106c4dbf50f24931719e1f9d06088bd4e78a4d8cdb5631f3cfe2efe4beadbd954d0a05f2c24a65cb3223e6a1dd855ba483a16319a0f538c7728e2b528d5b6e264606ef8e4c1e7eebf28535c3283176b49792027f0a2f2d7906d4fc795218a74003a58d2e0dd398aa051f12fd1f47e3adc018c30f7221e0c36e013bdbb0eefb466609f6ed04ae83cd87972c726ffea7ef7effce16ea2eb8bf41ff71e563c4b3eb657ce0cb1ddc55cfb677a2a18216bd0dcd7d807483f72c26aaf11bac70fed7f5f53fe5ed4bf21a7a5cc3e2f7a25bffe0e6ee2e03a17cd211aa3ad417bd8349ee3d43ad7e0a7df4505c023cec92d157ece9a3bf0a5d87d8ba634bb814b70587d99cd23a4b0952f28b5c22805cc9b9f613c1d3d89186b7a86bfc070dbcb89668110cf23658111ce46fc3c4d847e08625469a103b0f0faaad74fbd69e2e6bbe076c69adfd669f46a27ee9550d758b59ea995ef4ffafbec06ef003864e595a441946abef49964749eff445ca6d2d08a095ec43e4c63789ead67bc195056fbfc57423a6040a0f37698277a46051e738fff73ddcf2e1d695b2182f64170cd778c3d550bdc0243e38651f3f51e2f959d03451738bf2519485b36bf567531c2203454bbec44c5b95b6b90220bd743d434efb454a227c9b7eaf86fc1dd392e3b302156c773ec5b6e02611ae59dd5416bafc0d3cd9f2210cb2b4729ef741dbd2a07c67cb740085171f084d49b8885009037006b14cf6e95d44c258444a39e3d7665e98992cbc0dcf7588304fbd1d6f43967256a6dcaf3a6d15ed1030c6ff2f5f5dd3cf1735ad70f81d0ee4d229a19bd4dd566dac8b4b58ba1bbfd2799bc9164367dcbf1cc252b524ea3985f302be40b11ed4ea015fb19a106fa283fb759424ba0225689d538e75199629ade7a174dcac2fbc5ae944981320f64995cc7cc439db2f8f2a69d33ab381fc43f4a378c47b8f85181de372561e47f65aba5ea127e60c796810150674b00320063fc26c671ad2a378f9012747da49329a577fd411ba43012616c48b351c2ddc24b70decd294f76712c148be684a06b07ae4b2ad28c496ec273060da422880a290c16de473e30cfda50f60eddfaffa012e2980be19ea39f086dd0c90fd3e504e1a1abc727b31c72d22c67244d50feef830168ad8732cce1addaf80ef77a6df1d1de9b34e0c75a49982f18d8baf55753388764c22ced041dd584a969df53cb51865ed37cec9798253337a690196fb2ab95e80ff571d3543dd6a01574c5b8b6cf2da488e613b8971282797f91bf498a40a0308d796b9a3a9e2b047beb3d05532f6d62e6597a169fcc79cfbfe972d7b68da21ddc0abfe70615a33bd9ccc3e64e21bcca8b6c5553e7867ed09c330dd2cd1c7e09db5e707597d41f985ee644760a177b8259671537274c2ab8c0935202477b505a074536e1b31ce16a43994944041966e87e0f7707324f1ded5398d626b5d3a642e0584995ef994cd0a8b6d6176d03d685bc1b97270ec701e8906d2e14d57f9147a6bb9afd811cf1abd4607133321da597f4123994b2cfce5b04560a748380b6b55a3ef59b3b2688d3505ee0e120e49c0d000a7c8afad6aa49f2e9a6a904850a2a4609efb1b5ff2daddd621b894df75320b26336d025e783e8fdb1dc22deb10b6bec72882ee0467dec097e3cc9cc1b7789866ba142aa81168c73ce63171ea580ca391e6b8d02316580a2f18cb4fb65a586dadb8dffb04b2d66bdd65c00b9a3ccb2faa0dea3853793b6e83bce0b555afcc287313fa5d8f0fdadbd17d1ce55b7dc387541d1a0312c31957d012d546d426f2c5c8436a79a3435ecb808557b09c8f2414adeb9a5ef0c4e7177ce074b3785b94e49ee659d22514227b68bbb9e9a7c8b2f6f9e252786e9bd13f5e1958d3389cadf0710d69a3515a3d758661df5b00730b848d7988357e3b9b2973a7f67f2b133dadaf80199b91ff6dec896bd69305d08ef7cbfcb7f5499142e27a0cf4cc419c4432f66846a1db8cdd7fc62be8d5869fca17d3656b55106c5ea95ec9763c624b3342d20113980852a9c30de820817c4704ee07ad8465dd5a1612e9ade971593d8543b055181ed6dc720be410ce4eea58435b0755834954dcaefb4d762f512f1e1c46336480cce5aba96e55e09ed5012c71b98f2e83b1c2eab2bde14447d26103f2df204adbdce55966d1ff351eb5623fab74402ffecf8137f069efdd602e29d95d46623a05cdc304d3ba492f3996714570e1de7e6a481c8cb2d6b051743fb0b0f6c524b1d6f2fb4bb4a79796caa7f69e69ed812799e602dbecf5d32d638867100560aba200583651bc1ca4ade8edc3a90483e98c3ef56b9e72e98d234007789d38560159e70d7cc03bc4153a52d66fcc4a8b66a52c563aeb82aa10a12bb9b64eeaa9f5ae3ed03d6d07b983bff0f3508bd1aea545af21d077e19b190945395f3b11e3e1d4a7df98074bda40c87c16576cf55c18f98f4f68ec38f1e3eb43bc461b8f852889bea23653b7345ded7ac6abc9a8c2dc474db1ae60057ca185ab18ce9c1739488969e9340da91926ba98c2f0b2e019961466a133176b180a4060454dca3e190c30a4cc2eece8f602abd9c474ef2407025e4dfdba83006dd7b9196dbbf1792b31250b508aed7d2fe3f22d0b85970910717b1ea343c994e7526988c9109352e32e8f85bfddf48dc0ed58d8a977782accb1640f492b08b7b1d68e0ae61a89344df27f245755ae165dfdf0f3150c34544e3e82c7acd5b7cce51330a51032bffcb87ca4c0bbd2ac002de9bc4cfcc3416ed67c4b246d1461888cd579069bfb2d4ef787782e945ecac3df3be0881ae202113e5d2cdb3a60fbcd7ad1997646310155c707b58ec9176ec20b3ca667d6890882d5466d7c50114858a9863179365b1aeb70a7b082cdc350b47a2bbd656b656f8b5df8392fb20c6bc96fb3ba7cce47388cb18255900fc558fa8ce69fe20a14021377178c04d2e911a5c6da9b4378e790e2cbef48171266401a500d5c1ce528551e0dbdab3550a24475f3036f415359a82cd336d96d616b72e0300740e0a859fad56469c3e7fbb195e409c60694f7e1f85f99b328435573c4519d8877b14a60f2591aa03976a9d11d3cd05fe374b7ba64fff5ae1b0c9f70666c463f32713c7f1adaf8587b8686398e2f4532b8afbedbee235955d592879fb3bc0b9125de4a9ae090f04bfe875c4bf4aeb754a94a3944f7089c695fde693cb3f0dd368f0f96dab22c9d7b78bd51062055fc6a7965be7f70b68c1b59403b013f295267a3676d49ec23f2f6c87b0df53a3526becb0455d09bc800077242fc7c57f53068444c9088f6a146e5723764e4a468b6f4970f725746aa71889be980316e73085514fb8cbe28f9245fbdd5400111cc0081a9223d9fd7a041108bf0056cc0dc1b9637a67d2a4f9db3e7ee2a79e110118674af5fa8bccd7b90e67bca49bc16ca008a0d25319fe9a434958706860dcc51af0958865c274fb02512e0b43d64b538271c4d8128230282fcf1bf5081dbe809c96e07c11482f3231b83fb5bba956493c177ff3279c740c3d9e6912a23aa70f8e24d5c29bdb8ff46779b46bb1d5752008373fa8f0ba93beb61031587ea2505cc7d4f4dc6c5bcefb5b5bd1460b7ff35bf2704449caea5bcaa964bccb40ba9b86ac00fe01b2d1f2bb80f94b80cd314a3216500b871a8905e5c98ba16d229d30cd2bc7188ae53249fd012615b40cb95a7b48e3cbc3b2054c3fa2e0a2260ea0a047b95bf4b44c8d89b421c04ba363e0e53fb4e92edf61d12501576932873cd782bbba3e0a65829f6ea03bb029bbffa00b6c141172527c496132e67df247fde9c926fec6c858b08afe4a0a50d161fd0f8106ce6da16503395777436f5b5ff430a2c5ae8e9fc451431a3dca5d21378ae506bd3163e733d429e648b6341123d9e301f255982fe253ed9860fae411685177356e2ff0888e9f5e93380a8638241b389d824048935b5e701ef38bdcb206a8d8c5ee5eb154877be73e197319e9d3130fa72b7d9f525275d9a3d185d5fbf77047b0b691158624c42f77f524fed82b7b2aaf411aae83b8ee8840617ae038322895dc482606c691f8e45026898769a37b1712a331f20d9f45f5087667a68238ff52bcce9b4f3a4b0d990c1d9e72dbf08217e3319a94128fd67cdf7869519882ac62a5454a30e053d2b7d8e61a8439d38ca19595edd0e3f1d40b65ad70b29631b004a26e086bc0fb41102fb14de984ac8db7179e7c117964d7890bf7618b6407e074c776a3b68ab0a0ad9219819c4c871875d342c7f1a3fe6a6289818ddcd2d340e7efee101b50716f70389a9e6145e7d2ea6dfffadaafac5f5ae63223369e6a0d97b0c51b4239eca5915e0f495df6fc7349216a796c4246e0d3f3599224cd203a4fa9b68154854703972ce7c79e3be68a127b104abd8d66a6f7eb4a22bd38797c012c6407e6904a780ce70da9df58b1c3b35334b1ac2d68122b30485cf28e01f587ba829b87b6b181f1cc83a623d1cfefab365e2fe868c42c096559b33309126fdf3080a5d8d3c4def2958f6b0ae190a62285f596489dacf4c5f085cc8312a6a7bd362f8006e1992a3465d3c981d9365e7b3ab00166a2f555b7a8ebc504d0085f4b4c2ba32e82574684e33674f6d8a6c7ee9106fb7f491e828d122063331cd6fbdbb22c6ebb362e56bb95a40075f5b3ccef1d9c0e9c39ec5cef9619e118a6607d5122fa96080d5ccd34bfcc55bdb4d3fb31cfa2354afe271d860e7ad42e152d3f0c48ced9225038ec535cb48b5d9864c17ceba1e081ddbbf4d92b3fdd143d811103f616cf918607e9836dce7efe3473b2e076ab19b6364de00c8dd08497f9822ad542c35374695e646647d2207ad5e8aa82b808763cc1f20a86639b14db19c27b6a021fad77fb876960f47da128311f95ed16138d9bbdf01e5f9bc459cbbaca5a8383ca8335a4521b57a1775517b6b4af46634b3b8584b7b0ade8a81bcdf3a193987807bd9aacc4ee0a56fe036c2865159e6a737eb118f99f738b66603639b452c897ce1b1a5428dd3f52cff5f58ebf53fb0246889dea04147bbe89f9d8b0b1f33b7783b7b167e825ba257b10f10032021fba75793d978913dfc1ebf2cd64bf989e45a33ac91ba455899b3aa555ef02a896c77c15ec7d67d42163fe8815a2d07c87d18435c106595931750b848f618523ae2affcf4025b363e2c910ccf55d4629b1318be6cd6659a4cd82db111a6c320828e801c0012015818832b58e7f0226fcfc427156c378c7dbd0504b540361c0a6cc93a7f3874c8e4713117874d2c656b1e622cf00974e4a4543a637f52deb9634b84829179081fca13062c730e8320f880d908f97f75c51cade36a0965f49f354a35c92ad2aed5cba9728a03210e319cd24ab98e4afa92efbcd2b66ffc84b213fdfffe6e82c8f7919e217eaf123fb2cfca8dee267b5742cde058ef4a9eef711bc23e0d854a4636eb283f2bdf47f439000f833a91a646c361c9c25ab8307984a39f001de794beccd33ca4ee8448a091eb49ef49e1a2a3d68966ce686df930bd6f0728e3c452132b57455dbd0e9cc8a0d1f463b8543811087f1e51f9c82eb05ee0fafcfede9d1a98bd2cfe1dd2dafdc9ad4a0c4e7514e967556c4d5708274672df69660387d26d7a8baf6545661468782c2686f77c5b3f18281f68082bb55f9c95752d6cfe53eb0731b7b4767c262aa36b4dc511b6014a248d6c31a89a14220a69c2f126e0c2125a9fb30c59d5e1b5865b6c3e5a376f40912d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h97425bea3205411434c8c42c4048b2801d41af208d43511073993613a1f598675bbff87f96c9d50e48702a193cab80d96c6fb87eac02ce6535b574d987353b23b088e49b36026e781e797b9b5016331d8cf82217f3c2c6fd1f73a9a527ecf08d97ff9d9aee904547e4143a63e6ccc6b864a8d1ee8cd7fc51be370be8cb838008e570a49936900390b625dbf54dee78fbc045c7ad3375f1f91167ca5441296584b5ca86405b28b60f1c6c4f824a1fba1a0259b7563318685e3f969733ae4012506cc185457a6993146129334b86176b206e402387197e31a27810ed1e312f8c2838660079a3de82d816ce0542e16273ed236d1e2b697d717fc3482121e5792dacac8feee81dfa7e6f57d2c71bb4a3dbda56906fd04c6ad5ff25ddf259dce5b541fd1be50988d85778c67bc4ea3ddaccfcc21934638b1addd29b4397f7fb24fba6aff857551668e5806177c8b2d910d187ef0e8e4158625dd7307990465351ed7aa1f135458aadf49b9a696ca0983bcb6aacc742ede6900fa47f0d8c5aa8df5a19a52af45699663c39752f882d499948362af6c45d77a743b651b3c4f81175b555a5d599d2acfb2dae37a653ae75b056dd10a148868041b5ef44d25ce2ba3b61674569c3b734e7ace10487a96fe2276eb81b156d882ec239a7eeb3e9dbf1cffeca65dc4b6f369028791bba567da85ff9b305a527258e5d559afe916415eb19f33fe45a6b5439b63deb86e75f541fd174df9d3c30b57c9463bae3f0d8504dfc99ffba24e4a4358b365b55d5c51211265a80f6b41eb0015ce2e6da6524047cb95f4fab777b7432b95e2a2f34536265a5696895264544030daaf22451ebe7268e80d42935d70d88f1a97a45e98c5ed8012609734fdbc61cfc4cd365df225b820d5659fc4fa5ab9a1e0e186cfb45b5bf2d699d56607904d04e889f05bc9a0636fde9c5c4d23f1f406350f2d8a85c60971ecf9d10908af41ecc71e661b488e4b9ca21d4f66bd9dce02ad014946bcf2e95b3a4e58b081bb2adbc8d9883160adcefe177c2179248b663f96d0b84acaa6bd682b0cb93a3a6f0be462e48612de099867d632dcc468fbaeaf54bf4ec6b32bf69f9510035b52aeebc9e765b679ba6c1db6967db99ba43659a9383d96c417d5f37699463a2d9d3d849c35cb4eb8c15036b33aa01b5f6821c81af6ce2b00393b5f541ac9dde850ba42b66c12cfc86d8ebc3bc208ae148e92ef8f39df8b1f863bfc99c5d6bb14ae37b39d4ada734fba59ae5577ac9328a6322d7c8fccb4b67391e4c53082d5f2a52c59eb0e5059eda7d3562ab13d9a5c0868c7dc9326a7aff33353c14cde85e0a65188c1e3774ab0ce375981b3e91d6fe4d6ffff6a97e5a760b356622358636f519fb5ba76eb8415da3b037c85b305d2929c0916c2a8b809a9164cbc5605ab1c582c3791370fc975953e867942d10d8247c036d2f0ddf66cc64bb132e33c49a2ada02d2d62f31c36318a6c48ecf58ee83c4ada780800aa41776e5dfbff26c19b8d701bf88b632dd1a358c6c56949b9c324aee3cf92bc93a69c22934c01f9765f8f52521022e3da12636ec1fe17171ed1e5ee52f8aff9c513b7ddb27f671346589907a8a4bafd97443a32ccca80ffee33f6e71a98a7d1cfbb7350964c029dd3ea8611c4c2f5c33b2fd5059948ca5273c9fe29aee6849413e81a43f68a79bcc8dd4c7c256ec80f5e164132af79513637d654dee96cd0378e1391433d1f93512befce29b75c3c78a8ab561d97d54ce2864c2ba6c35ceba98a6318e102abc334b06c2a4e172ef51717f630438d21744434cef7973822f9f5cca3addac90f5b6b06b57086f6c3aa9d87b561f620a5d711e3623060cbd82ab0af285009387bba36982e4d512b837c6f365615522ce9f90fcb9766248a0ccccd8e5d73d85c5f987c4c13062d3fa4c0fc8d107990f371036067a98281085435b1a7ab97e563892de6797ba608967c1fc9243c68d958314a9fcebb789407b6673c84cbd33c1a5909b94ad38b4b59083bda95477d425d223554e986024ac19a7535740888dc8e72d28926e258b42836ed54df0572503ac4b9c129689875b355203f36fe572ddf4f07403902317b2f0989b550b953a3ee4f9a0739cef138bbdbc6b0cc6d287cd4284baff07c59d0feebf8252d8371a22d1f5420cf1e19e2ecccef2e6a21e657d959298ecc4e3b56510cc4fcb1bc6cc4646e545f64042f19c6a7f6bb030af468c1abd7101360c8f11ed13ad3b23a22aa1f6d2b439f86d74bf836b3c8fd3bc1a3ff9a71e34d72af3ae392db656c2ccb710b644c2458d40573b51dbfee4c465982d971c02dfdcb6bbbb82a6188e22e49d5a097c10bb782775243e942bc937b95c664512d009a8f2c28f1c3bf3091557b0cc02a042b05a4eef816105959edb2160e5335627a2254b02bdf985aec3ada1be64203f0eabce3c6e446da496bd78f6b2f6db249ebe3c1db11d9a38d5941da1863b693592caac3ffea64824235638c878af557023cd1c4413d299e97447608a4de7f7f6fc642ded07534e2944f6c26b390579504264a5622132000af0b1478c8d8245cbdaa839641f1c43dd1398ff2d059dc80064c245715154716cae64fc17c7313cbcd55c9963b75634b2373e3230727508df6e1ad5a248ae8ecd7cf3459d1c77d2a81694e6339c4fc06df7ec8606d855d6ca6bbd799bd5beaf11b6cfe59fdde0f7f20a1756318a14b81b4cf3d4212c64f20df6b8b6495389459e68a78a4964685d7385dbeeb04010d4bb9b86797d7ccb6a345a4f310f416fdf1f00164274a18eb544c5666379ba131862ce48ed9a0a02f527535509056934dcf6a74835a67d341aa0ddd90839704897d3cafaebd2e3ba122f5ce98187c3519f405513d144f6b8af96387096c0a8143fb2ac41ec53c268e8e466d67ad6a532e5e55062becca113ba47e4f683ae4c44cb9512bcaca6b9b892632049f7d64fcfaaac6ead47f699691e410713354dd4bdd1eae2056d1bbec259c6f497217dfb70bc002f253b99917b4dc7e78402c9800935c384e600c8626f34b40be8338f625d21a78ed4ec6a133580cbbbf2fe366b4a00d81949299e153482b56c7ad6ca01ee5b598479a642f236d8655cbd1bec62b20bff68dac77014e4f88f7942b10ce71b7cdabf8c5b6ff4f9d9b1eee0d295e255fac44b2cc7ee40d85dc8d24cc91420d97b2ffd29adb531309f429684321d170f7cfd2fcf7ea1bb55715b9d02f2b246c603b87f55796e2fddbe7df6afc6692d5fb6d075b3d542e955b34db0cc6af7d92b0b804569861f2b65c9ea6e1e991235d7cee0d7e4c177d0b3af3b1613f93220e485c8592eea13c42c420915982a182240928c43e4b20d9ee039e459826def29cdca76043a453004599014f8a3ad68c9be004c34b9a983bed6a064220027ed13c98bd111626c8b9e1f2be76765084d1a4740eb399d35ff96408707dd6f71c3fb0178d788555047cff01d7a58c8a8e02ed42d67e00c012510d906e98cda4c6d4d6811ecac8b47232de554633f8c1ae7ee1ff985799d439571c71680a3b50ea863c136686b40c2f6f88e8afe834513324193a30d613c629a552c31cb899645ca780bf2c6324d929068a90644986d5d84429c251f327d1a5d5469c54d969655419fdfb174279dceac93c357ac6964c37b417c78d37c9b020cc07b5c7a3d6fbb4a0d9cbc7758ec333c109d8d34dfca09495f2a2ecf28c2730461bca7e31a65f560908b6b9fd5bbc9e52f36fd5ed3b4f44e74c613156f57ce5ed7ab469748abd3ad3f0c77dca727d0b52dcbfea2971f9e75d6a50fe90290d7669d58851826fb39a912c78f204d8109fc4080af88ef3142bb86525111b5b1110c8542f60d2ad8cb19b06877abfa62266d462504f9c972d76239172f8a005f8e0a44b93449897340961e9514eb6751ef6a0b9558d16873b432146cadf7b21a3381a4938aea95fde4fe226ac745f68836aeae1d4ab4aa23f2025cfce3a8bdc0a34a31af87f9f0925cb3d50a898c4684f561d0ae916234e2ef7e3c9c9dbfbb9c34d560bc68ee328e65418ad3577e07c2f4346887407a9e3c003ccb3afdf9a30d755cc9189eefb4691465963d08df325962ab385f52bc506ea07616f9a68b7dd0897866c83489a349a2861266026688f05f4418e342960b8abf5d0a59800783aa9b08482fe6c493afa8c761e1b14dc5a8d85db395f7b4814883dd389043130a26ba2673884297bfce21d12334767db34d060c233fe0b74b49c342f2b8aabd84e66a188eb381b19786180251d7287e90288fe267ad2553cf3d76d8db41842578f8e2df8f1a6a80c8892011a3876c3419f84c488019cf0c906e4eed88d4c5611661193e4dfbd268e58801413c52deffea1ef9352942ed18cf7ac087c442d2f3471d114a5e1e77f27ca630e206dee79fb515f5a1083bfc6922e87f3ae7d88eb8fac944b40afcbb5f6f621afbdfadf152c94a02ea67130d2ef141c124af2b3ec346da0a0c6237044cd62870a614cb84e7e000f1ce0c1e58a4660ceb6a1c2e0c400ec300b426f8a66a4740bfe512c18945a847d833f691a095d5a2246d18dd7740fb8cbed08625e8b3e3d4e3f21d95439e7009f47142fa4b3968905e01de749f701d0ae20cc5dfe280e8174e9f39faf310a134828806fa75779ab6b070802b9d61a3033354243efee70eacd3709943048616dbb77b7440d6454a2fc097c603520bc5cf82ce9b0e9e57cc10334d0b7879c1a2db1067527b607eddd6bf7ea1438f6ae0a340902c3747cbdf00e4499ce623cd2f432fba1c69cf33873eac7019282ddbcd9eb0e77a8930b0239539a54130c1b50827e7bcfa24c4eff9475d54ddf408446fe99fba0bdd6536428cc7c4a118e1aa1cb056cbd07da56d1a33964932186a2a775ac34068ecd775423e227f213ab244d430485c3da9b4818e395c10f6073249fe926e3a3cc5ffa3d4db6435db4de54e5bc5e43518ad1f24d5b89762ff478cfce22e25d9f88feabf0ea254578ef7e610853b65da283ab3627bd4e93931431017067448f26b9deb33736f4e4efc28e5585571f054c8531c34faf182ee3dbfb53856436f154722c78a75b62a1b7a625be2bd3c4e266c1429b1d27e62507c08024307ae79a229ba0f545c5d133f0d83226622bb22af2b7a5066d13a8e4183e39fadfa064c56c51da49c52963f1738f8ed1ab9384a234530d7958fbc3dfc6f3c831485e41b62e5bb204ff07b225631d57125eed0bca8583d92f7951fb792053f975a25e740155ce7d1d616561273120d3dff783a47095782a4b2188c7b437d7a4b3b921e3222649f33410360e4d9e13f555f687a7241b1a9b51e7b7901551c431d89966b0ff03aaa5b5afc6b5237a23225204ced87debd143f8cf7a8ba5a82f26d00c9c23f18ef0dfeeba5e7ca89272c85f831312908b52002f3b96b82a05cd49cc7fb94d1886d3e3f0b83d59ee7420c06bf80d345b99410edb1b6a84eb2336dac23b59d0d4981d80309eb6cfe048cdc0f1c099398b4b4d4dec2da5585c57ffe688c37ed779a1cd1e2ccc79e9dca4ad4b80a044ba05261d6114e9300033805e26350022a922ee9fbc48d4b81620e91b190b56a1df9bdb4bae84ab184c279ba2e7f57c0c0d68aa7772117ce7db066b4b65236fd6f9d7e4728cc190447c3813ed03add6e69341fd3d2c9c0d1a747497b80df07d743e7c8cafcbfd46a843fc981a9637a5678c64214422fbdf77970ebf180a7c7eb268c5af129e2d96afcc2eb551108c2768d1209f316c61a001875f7dadc19fafc95e0c6a17cfc7fd7fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc6af7c2854614262ef0388a9233a876527eb9557587bba2f1bd42274b701a20b1af398ed24fd51fe35d834deb178749779e4daef375f1015fbe20d9341b7c7445347abc1c04a5e02fefb8a73917eaaf0ace0dbe7d1021a91ae361033bce2a7d8ac675cfbec58c4002549346e2316a4057c5da4c48f1d6d7b7f765f79fac1c4d0746cbcf9fb818d0825ddd4059c67517c37c532e6bcf03d6fc32b57d2cac70d9f660f5411b6e97514bb6607ae8b67996de297bc699a268dc760b8d3c77deb86219b57c1e5e99b677e465f4032c9d922187faab819ff2185c01469778f1d9160d816baa13eab82e89d5f718a017612965f05927ffdc53d0934d1cab4f7b9e9d2c34eb04843b7fdd16c5c50628c7583fe0186280486e13447786d37b9117d8eba9aab57ef5efc6497e1a19767647fe4ba6844076b526781b3e4a1faed8473e2662f9e610b5dd8e47ae85706fbd6f1abae1816baf9935781ec9cf169eb3d821bebb61f429912656b88d6865b85a4d61f83f1d70a36fb1604d6f7e8634d93e239ff0676dae4f2149d12f3b667a7b57417bd1b1b94caf91bb1421ff08ee047d30eb218058bf3147c3a98483a7036020fb1312061089db18b1ce3c04a81a54e7d4f91bca8c49f4b6d7e2da415f4f9fcd8371ea37aaedd46f25fa9e427b2b98d41610e08d1553a16a81db0f88240ef4e9774575a0bc16bb5408534d64d63cc64d1244c440b86f9b546c499c32ac2fb77bc720864a862c39a1b698c846afc78255d7e686d68f1b5fc45dcf18e4fb57de3b69d446e14cbad781f2ffce0625badb68539f4c0cc42903a03b585dbbd97e259399a9e423ea584f6647c6d5a5b58315f9ec11a9551ba80936fddd3fedc53abbdc2146b6e42947df5a32bc586fe4603b012168a41ca4957754f553410fc10ff637c622d8a4c343d83c21c84cf3557080ede9733b75317be226b716c72ddc39f52d7f26f0db86cc6cbd2bb3383a7ca75686064a24dae114e4055404000455dccc24506ec6495fe9f430235fe7a7f06a0d046b97bf4cdd1249599e6cd96dbaa1685905fbcfde4a9db65cad5911c7d45b9ad675f5889d1c3eba605ffb06f17994043f1c4c4b6a591405bc736f52d7135b1a4c49a0bd359e93bd9b9d30a8d110006acad73d9cc7001334598ec9583a4af5f66fcabd371466e94f4e1cbc9f122ff9319a5ede1e3e1cef2462fd26a501860ec1dc2b958ab7355a4a6558b0e95da15c4bbd7d576de451edcea5345e75424fc452c3f8216e74ec5dcba45e48e5b288a066aa24e7425ee4f990cdf2a3e479d4e4bac6d7db052abfb0ec567c4197a6b5fc95afd75a38f4d1f74241eb2bcb0d3bdf2d9d30a14982e30b1af4b5693322ab62b837f1df7db06dab399c94f6b1203c400348b952ec87a0d502b46da86f5780bd694851ef8f33526d7d11fda7715e95dda4c0a53303d965bd59503e40785445c2d2031932b8f3f3803bedfc037458d5aede5a366ae11029b75df3ae14484972f20595e6f4f44ad05cb5a1b2c842b6b85e4f52ac50626ef4748ca23c48f0fc6ae1c8ef72607c388a00e9d0f0f6b7221a70cd13033662174efc203b4fd9af706e7d9b3d0c353bd20bf6f8a94051a8258f5f86b237342a04bda1ffd36fbe9b9683f49c0973f6e94373b5d9b4b0d43ca7919df229591157ad2285823feccca9c1f86533ae9a9624bd654066d3ef7a7a11123e23ebc5039b7774eb8ffb897423892c7343e76cbc06bcc2c75bb8ed2ecd158ec95d994632fa76a4e158839656d514346b275b380105c46b095649c98b69b98d9eddb1f37caf1f78ea1120c234ea25c280aeb76483d5e1f78aad5864905269c452e175091455ab268e2098a32aa1056b5fcd18606f95e1a52c5c0e961c1dca6c4dd6d191829c1d5e14c7fd611ba4b16f12c752c8dec39d80abe4bda9b87e0d06f842b25b28fa0d4f1d99a4d67b8cd8f963f2ee9bb9a9819556c4bffa7899538c2bf1cf0386c04e2206a00119694bf8cc26468046b0b121d9bea334f061fe1c1ef3bdfb38fc62de655c225f472e98fcc3c0a22983a22e914f0b8308c6feb1b743aed0012c7ffc226e214536283d66339a5048c4ac4d7cec65dc24fe4c9166c7210a3c4362d4cfcca50e40bf8c58d55c3136f5e13407dbb2aaf8f180396a6ab523d922cdc102fbd1f956cf662003dc3f24c42e005b0e86742f70fa09ad20501a5bab19da9e8b74e66ae774ad94f5c12e859e5b46b04619a4a0d46910fe91e79feecbbbff54210734a0f67c73e67df04d465449062b7b7f1b29d0bae0225cb9601037d1043404954672e26b227222ecebcbb72ec3a8cb47263af356ac9a77f672297f1ce36e7c6448278faa08f5bae529facbac5e15d311d443555aa111992d60827c9f1d12e1c6060342d5ef0b65b68b4b74aa61b10ab135d64ca78de2f79a4154dcbac943e5302f7a46b6c9872f675424375fbaf935a5d09d864c143ebd098f710ef341651994620bcd09684863d37c065222e577c46011d06c42afdd5f1e909accba3892a797134c2567499d206ae34397987aa33956ff4e1d7c2a2dba14ee577cb63e01c0af9bb521b1387e575b2ca5a05b19abfc04ff6ed06302f1a9bc397ccca280f8f58eb283bb35aac1b41d48f18af160ed74ef114af5292409c570572e1be7099676d6d88b0dc49a8e8770cf4a0b2931084367e16d1eeed8adab5a38be7892fa52b7528463aac4b5ce2b55a6665ac539d55c5b9064e1b10326245b0bf43c3d5d053c397f9f5f95b0f01bcc3c459d340937afd8612a4f5b6aa047ec4916ef5cc8b917355ef87ee28dad226aa77c5b24737e1e4073798e206c883c4e4b71b3bcbb1e32a36e08a04c92a3954d14603a78a8482ea2492759d2cf0112c23be941b6e70a296719742eb22d2c4bce6efff3b798f87993bcae92d2d4a71c0ce1b92f0d4974fb5cff6278524271c26ed737efa454f55fb50c131c5ef35eee46632e4165199da5e1ade6f4dd26abc1d9521706234f414e422395a3ebc322c17b528458d2a1c7f99d6709a39902a6bd48138ccb53132b0a8a6ee33f7544d5cfe677cb07bfdfa15a89de872bc1889f4f0712b677fde91b8871bacbd92dd7ae372440f5ab2045efb1c76b3a4f559a157c69013e13fd5eab31f7329347c0710b7d011daeda5d5d4346ae211046eb064bbbc4a1434f5ad1deac4dc0553d63ba8a002693979821b998a4087d47ff88c26113fa2b7e94ce9185e5058b17fb2903af8876948fcc64387a8deeb0b2c56ac49f0a0fba27fde48bae61edd04eaf0d20d9065bd3104c1e0ee14d4aea9a3fac1dc067db2ee37d18f735a855769618c9aa6fa7dff91ecf61d40784c0458592fc48f421dfdedb250208d222b50d56588a2a607991d973a2cc8be3e7bb565b3363d318db7d911e28cae095d3912d6fc8cf43c66f27f01c0b0dc776302237e4cbead8ac6633fbe1ac90a67c7cf4af059e60da9694f0cf1003b55dffa1a10edd431e75600822ad14527274ffce28010567a655c97e449b7774c209202b7ea6a0ef3dbbdc4d9aa787eeba4c348ff92ea5f2002511a5652231d9158488e14252e55b5431e85b2c97de63a94b3524ede952b0b881de289f22ce564b6621bdd0c52ab17d4251158dd28d81f70368d064791b21d1f7b613ea3216799a67c9511895796d4f97b4bbdfe98fb871a45a41a0f833766b3936c736b93bd7bc0c427b41b7ebc9b8cec1aa09b7aeede0415b92dd056bcf1fb5ff06d35cf4b9d3880ffa0b6252949a1ed377f63a3d003b4573bde783fe40dc1656e127568e108c4460ef2e4fbcaf4292c90690c271d91f9f3de1e58935fbda4a7f17a46cfcbfe1fef6f24e1d9f4c6de319712d9f2919dadfe263743a81d53f48ce30b2fa83c65714cb9e1d46a1ce2188b4e7a705323b2501f643ffd12d3d89ff78703145533d5895c00e547e2966d37f4296ab1d95cd218312d463920215d4b92ce77efcb26bef8ebcea35967f78fad36ca3d56258ebac2f762314e258e653f6fe398a7e18a7b4ad0bb0a53feb255a58f8b20ef8491a2807bef03f1e475c6009c20f2cb83181e86ddce6ff1ad3505f30a35c7bdf6d97707260d51c67ef36b7c29705b2da7d0d53ba6e6556a4dc689d4867dbdabd7ffa95e76413978a63c3a1d6737ab1dd24b58de9365838b1168a8acb4af9637e558f179f05b74c6ddfc95d5eccd1eca336012ee73de138e527194df231b3a1058f3baeba10c915c33f01b83f91b2099e33897e58a10fbae52487d5d703f84c112f5e697b88660b90fb1692361129ec469a96e472f929d38908cee4824382c0195dd55785a636a78b418431436f5fae980e375ee49b80f45f0ea3b679768e08c1b3038853ffad0bd11379b78f0f37ce6325af2e840c3591cedae1a9ea7df5c2a954bd7c20b47e3911ce7d08703de503353a0a51478ebefe2c538987f86e7341dddf6e12d1c60b97fdd4ec893551ad1f3379d0a8723dc701d2e63957236f147fec2a9fc40bd9bd701c5843cb379cd85fce78ff75971e6725a9a161bb6dfaa90fe4fcbe29969f6061e0a790b03612cd8762c9b9f84456818a8f6c9dbef6f194396ef879a71e7bed80aaba8cac4e4b7744f4c04b873bf8279cb98d49d48df91208e8b68ff256e89ea995f10a430c65b0c4f5a50d66886f351d538a4468a3488d7252371f81179858763bc395c74dc6838c0db36773fa59d12cbc3d44d0f32df182c34b651fd7bb8d0206cd6939d6ccc07069e3d8279ed48a69ac257192c1051bc4332d619e14dc8cfccc6584207f243cf11531c455ab7902434bdd57fd675e7a619e9bc8c6cc777f09efdca0d67ca9190dff4152fd06f07c5773f32794dc5d63ee484ce4e2170ca8f65440e5d12b58ef73975b8ade8bd3922808df9d5c2f69b9aadd35f12ed6562137d846c2c40ef9ef38030299926e3a4b207be2ccd3e5bc3c9e505c087b46ee68fdf3cc7b7fc2e1515643fbbe2a9239246bb9c690476b9965fdaf008224c42d2f74148fd8e98fd310f3f0a04513c4cc089e08029f5cd4ad4e21bb1b8156c9057ed419a9e2174ea328f0af2a1db6b414dc59ba961837725cbdfb0e2dce338f428137d41f7815b0eeed5f411507c09dd3544a7836fa6bb87c67bb8c0ecd436e3531b2cdbc8460357613bc9f816517017a858da8ca2271b40410aab49f183aa8e920925be255c409cc6d23fb27c628495b305b5ba51c41e8100fa5eb316e057d71c32ef394618e8d213be1c2ffab968fbb92eeb991ceca96e063d62c64e6657dd8c1d03d173b27b76d6dfc644f34b46530dd3e144899e825ac77a0bca0b084b86fdb70c5b0c00303bca5cb1bd5fe421b6efb121ff458fe036cd151be1cc63dd01a10e6f5a488f085334fb58eb423df71c8b99ba1d9c4b5990877d333cb1ca5d2f17093285fc918679556636636866872fa75fabf2234edb15fe8e6fcab15c01ef8e2da80d8bc85ac1fb2e528efad492a2a3347a036dd2ffd6850718bca44c3d6186ca4c8be97d4d435d5f9221771ce77717538f852db23c2ab32bbd6517bf174b006cbdd4838532dba74455d12cfd52470907b3db5100657de4ad202fcec4e2a0949b9b575f24f219d05a21a065b3e66e0643e651e0ca8969b9971d73c21e90b806e057437a9b41c370c3a9e6b8e87e4cd67192905bf8da3b20d0a22064bb0583955cf4d30729b3d288706a32462269ac3a9bcc9b6ce3f9658a8e2844acb40426f81f582d19999a89fce5cdf90d60c727afac566141e2218a51d29aee03cfdfb757dba4dfc2e6559f09faee626531a923bf7ce7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h221044ec6d82911cb4cf8c17b8912351a908ea291ac43420137917ac454bf72f90e3ba46bbd792a66659eb514c4eb45044cc9749adf6c9793cc70ff3d27f7c23f26bcd4152a506e5e9e5fa1a276dcede8d233b1332a39f648f887229b54de8c13b20878adfb0d8eccf52b3f9b6abeb836fd302d96163a3e0bb3614c109762bd515ada53e3368e74d7624185636c34abdd4175fdcacfc2d359a0ebc03af95031a4ec3a498571d9397de1703aa07a3d37128b967a5da1009a40eea0869d695cf85f97b9ac45d9c31943ca803581c81a60ecee75c02c370ccd02298ff7b9df8ac6504335ed5d9136b860f3881ec06f8fdadb3433b1bc63dc5973014a69149b0b7d48c96a14b32afe96efdc3d07f478a1ddb46ef0d6231dcdb719f31cba4281ddcfe0d73a54e5150499a9eb861cf2516facb9d34ad3e58fa098d678dbfea8df345dc7fd76060e87c98621aac53fddb66bc807294588efc79d4404232e242bc6089c538012b8ef7f971d643a39bc895ffb1bf7aabdc098d7d08457d2f7678dd7b14964b2e9f368523628eb60bfd1583d3206a086229c976aa04a7acdc64d442ef3e7ac7746007aa7851a82c1db9d76a80372ad67d3f3a17a1f72ae9dd3c89dc9e22b69649ece2582d441993feaae4ec2301c1dc24fe5f7f08254d23cfa296cf4e84fb4ed58e76d32fddfab0ccdd96a7f8495585791dd817cd0a38d288f77ff75420804ee138323fd6bd8b01bb616574384ba66a646afa6c2a169f34b82e4cf35115a53e5d35c4a9d92ee6b54fe4c406906e2ae987d12f71bc93fd2bb265700720f3a1d3a28fa20a8df06af14e98a11773301d14ae0b05cadf968d672f3bb4681fdf74c31a72d02a9f0a13b8003b91554c83f9147d56ae252883ed8f487749bee570b6bd310ed80abd4b6cde5f89b317f132210ea3b5f1e869d33ce4c5699adaf764aa646a22dfff3962e5af8287c845df2090fe008d55b3f8eb8eff40dbca915819cbca6a0e71b1f827a7b10fb4ee1ba188e0de4fc62d8b4b631b91ac3e46fbc500ab55d221079c1901d777af9460cd56fe7b35fc2334743424106a22a34fae1b2549185ab36de33c27744248b970d265e0a7d96283f8c0c90f9c3425ed8b93ca2f1423f30d7ab2ec4e6b7dc025139cd78bfaf808b3d922885d9deced8649ff78ff5e27554c3153e340572de68a90ec359b8113b55d4672d188db24ce3c827397d64df8e511c71170e7cc0335992228f7952ad60118c8a51ef95a3718a8c79278c0dd8e92f29690492c3ee917cf567f7e2c7a5e48401c6cb41c60349c43b60afa700fadb3f3a65fb0b59207ebc7db139f7acef91dfb8d8a6438fb3085b00cda4150f9d341e8f6f609e48a66a5039619e670ff8bc2095f2e987080218069694f3f10abcd1f053d9e0ebbd9cb4749e4e677ca1b7744a96beb8009f8e60005b20f5e0e7309849c3188b419dfdb89a7c0cc44335375f25e0f1c71ebacea2ad18487c83f38b415464a376e60dd9bf274649ede1bce2e35b2c398d6bc957c03bf914f0332ac193dd1d034d53346b084b4005b8edf79b012db856cd59279a9652f2a0895856b5df1556f65bd5c5c182279a25a28d43556e9c54614e0d2447f14f4c3f3f4b8fc06ba1bc4c4882b83058ba1722a5c9b7ac9a437d86011c6c5b343dbb87cfd9daa2ac921e137f19d8190d92e375472d9cc62f1aabe633b8990aed8ff91114e27a90cfc31a0d3bc30b3a205c43148ad55ae35cd46f2271818e22c6f23d44c6db08485ec26d5c9de75cf6a013723709450d3cd8771ef2001ebb65e997a21ceb04e43efe05b553dc4cfae6a76315ef8ba8adf0ba996f2f961dfc848813fc4d6d4f74ce259fab801093bbb4c103429e114b47696f5d5b4cb03a15933ae2cd08c632a727526389d9fdfe836768f44bce4e8b5b904d41b2434a3c2b7d5a7680cb20e25aa30473062f9bc4b88c3bb0c554e9ac65102066f4e93293f91b9d933894183aedfb060a1d80e93b7d1b10e80a3de04b81e9a24b786acd854cf9f071c36a5a7df5b80c51337d4d3158f59ea88614b9404b76c87144087a05dd6c6b57e0d7968672f1af04ffdfb1c00e4734eac1506bb472b47a0501dbeeca2d2502b69000a5e42cbd1b4f3d58dc613a2c2f354360e49330c8448cca0637a7561a2aa049b42d3bbd9e131e1557f4d52e7987f0b872017edbad5db80c50852009650a9823bd0fe8b0039c3f184f2286f9407b7417a4e984d9c6811ea12e2532f0151cef6d4ac8bc37a03bbc5112bdef1cd19c55fa052704d430f4207514e1f40faac5a7f598c9450692fe49f963ca2701304cb56065add6f03dc2d22be88f20e5f34539e4681d62cd7fd68b0423804c26214dc149de6e7376d87a54a8e298249836a181698b8f6f479fec10ceef98234890b6e5b458035a2c033920c54e854ed3c0e7db3e9dddc66aeb3f53d1b2274f6271e8942dfa6334a7e59dc007ea03fadd334a417268d48f22a781c70d7785522fd14b30ca4921a311abb25487a5b53c03199ec30a9b1a10faf202b230e113d8ed44abdf7236f329f78249706a0fb8d5ae029ebf57ee0ceecc6df00d085f24399e31acf7459e5cd13149f16fb7eee802cbefe7a78475d1cf30bd221b74823cab0d696d0ed61ceceebd9ebd310af32954705838066187bb92a66667787a1007f7cfb7c27fdeffaa1e42fd8dd91567e76f7a4aa4c3a0ceef28e491f5105d25e091648a403d5dd18c158e4cfd5a8ddc77438ba5b7b653e0c0746f9ad35ecb5a93b9163b8e05cda934f7510bcb53d7786b592aa17173f4da71e5e1be217ec187fb65ca71be9bafe39f9bd97fcc921f6ed9c2085c24d6e551d6c9380c76ebcac8402ca8137e3c0bc4c63713420eb7fc839f903c5cf6a2eeb17ffd5befb0532016205505cd678dbee35fddb2cbfc1920a7516347df4632a52ebf526ad642072d1fe7b2b21457134a4cfd364688d305ed2231852ee3043b0cd0d54eec2d6a229877ce96c5a00f1a36dd8596afa335129bcf146c046215b8b8d1d18dea612438eaa5566b8e6d188bd27a9985edf94cff6e203946f70c075bc8e71f430ada303e26f2df610f6a9906be1572dc33136867df407a598f7b7ff474dcb5c5783e93a953b96801ac649233eba9872a2ad31938ab4d4e17e36dd0138fef52cc43c0569f19c099a8b212b6f6159f023ed718ab01ee874c3a09057366df15045b83430b5465ace60d89dbc004b285c2466d4c3fc7515898c36792a79bb0cc12e78db16de4e45515c553116dccb30eb1129f906317288607009874e3483d19237b415db3a42c7c1c8a99c003f4dbe198d968dfd469fb1a73839ca683039b3d856ea887114ae619df9eef898bf35c8cac0a70027aa276f226dc1f828dc437d45089e88c95fb0bdc4a057fa3f07fdd2a3b101e2ac7bfb1efe19c503ad7574d5eb441a1841200d406f71745ce97cca9af4a3f62028480e5e4d1aaf05bb5127d3e0085049ddb9c3e9ad88d112797beeda381e20794996ace5e421b51c4001bbeca2749e0718934f417b5fbb05ff4a581a148bba178eb64f0822ff62262d8b70c9e3ec48c711df8d56f92cad1245884d3fd1b96748e5ff04286e9362b15091d1b01264b0b1887c32585fecc3628814058ff541d33d92e8be4481d9aa54cb540f0963ce2d7ba0f6254913a2b0107d4e13765625568896f6866d2cbd91c0dd668f9f5931c5626945ab1816153cda5d75ccda5bef0e4fde262c0301e76d75907c3350e34c9ce36f8d1c4d298e3f6ecf6cdf4ae015a15924f5e3c2835aeb1725924c66ecdee1b64ee8a0cc0ea13355a7c6db5882f2e3456ba9fd5550359b5093f69f8c0a9639fbbabf0e52a4fad903afebf742f596b3632b39a42a3799dc0dd33e979f5ca1503d55d0c60e4a9abb3a3ed44b0442da073de72873f2276460728b66003a7cd76ba2006b17032b9d1f9931246a1b16495f800834705523c39d5a7f1a7874f8945e84d41f1eff5c898e542e86bf1f34601163b20f05e22a187179aa8d465fbab1e74f374dd10d0881229eef6f0ad4ffe86a71651fdebbc60ce9c98463d91ddfe32e72ec5f4eabe591bb799369673d1741ff01d735200ac537a0ebf615a5cf7059cec49972e831a227c00818c82c509b0509cd7149a07e21db2189989f5628cf33a8b8d787457501aa03629f8723aa958b5e9cd161a232cae10fbcb9392ae92b29c93042fe845025a526952b26a0e0c9deec9703c58f664b1e5597bc057d6bccc8898a894495b3ae3787fb3c736d3056a4ab18cb785cf84b1a4c74675d1d822e76d29f206c6ef972375e5e0cc30a7fff51a023530fca65be75d47167f5d43194d9952905775f2518fa4e080189b9e79211a9f2f4b478a88eceae6af3926505636d16595dc9cf7e83dafa2bfc63512e55213cf0da6c2b66f87345d0d621a0345f305708a60ec2f174caa56d6c9d90bf1c4f14cc5802e92500ad55d3c837f49fd44e85edc20eb0ea2c5f45ec3163ea5910cab82862ef7537b9df53a5b4f5ce3732f795c6f9cb1b5098d6028633757bd26d428f26b549241e5f6acff6d7328d101688dd2cbe5829df1964c61bebe59d93480f5dc2cc5dde1d7068575226adb572efd567ab9a5a172e33923af5e9abaa2a0bab5eb0b814c7e5f30660048d04ff308857e7028cdc87f78253b081138c0410f858e7010dd5b0d4fe9913a4406b6261855d1c68702c3bc6f06685738f2636dc3d694d7d05c2ac1df6baf61cc20996c2657b6c08b07d8559338698f54d4022c9e23d4d03d3d75bc72c30ce3895a30e643ae144a76d835e213d825e530e58d8c7303492e8c345f84047dd2433c61389a02ee6a47199a89a6128fe7052804dc0e0888780bfca3ec059cba1d068dcacb1c19e56670d62e04e0db949f5fe0b057b2e36d7f36937a5dddd527646c685b4037a6d72d8b559ffb81a53c859f9517c287e56a2dcb7d17b2ff0056a822b89b05a0cef3c59d44ebd889a427be114fabb1878558770e5e00345025eb014ea588f85601ac8fbaa2aceac8a3e71d7a2321670e67ef6738ab0ad6a428132df68bd7a1e1c6409c0fd379a7f8893e3607e82cf560b5d828b559dac941db8a901ce7f45e257606d80769efb602f30167927fd38694104475af9a66045f3b02a532e0bf8271c2fb0498d1cdef1136ad04376125e49ca7bd52f2493bc354d1374f3601746c199ffce8dec5135ac8bb4e947fa13ce6de9c4de9f9cac10a3f5ee95b6aa87466894cb0b7e37441d00fdb6042fcf7c40aebf0c7bc65d7c5e50b9d3174ea4f3a4b3dc871a5469ebebfba9f5288ba728e40861766bf835425fb8b6d101b34b71dd6d318f2d9c6545fbfa6a40bc4f0764aa053e1c20ce022522f582ceb7f73b77b22968fc9ca919bd2a9f8a7d446417fd4052d8631b13a8753a00f054a25cc308834c6295b3e5b71598807f8194b189fa17ec7a10e03bc2ccd2b376a0ab246bfc5f07873e3b5d4024db833f1f8e7720a28562784dfa86c014728dcfe08298933b65b5ba217b4c25d3814b027bf0fc19b5b651eb121377b98373a42f70d4a2147c24081c581adac59fa5fc5f983fa1b071e01e239abf79d6ec33bd383b7843002b2b2efd9e028cf06e89fbfd17a6d7a35454410a629b3f59c9e02e7efe1ad036901d8b998cda2fc847c9835426b8dda3654ed5febd742db85d16c5aab281f95026f575fe5b03c070af06c13134b216895e1215e79e580775f27351969d117d95f3809817dff51e683e174e38664ce086cf150ae8f382397909844f003c11137c4070fc2f5b1e2953;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7f0b00240aecb0b9c607ffb2fcc42d4d2e44361a4a38738b3ea416b2a129ca14afa97ebc393395045d2192f53cd40191f0d03c45e560a0ec36e13828e75bd7807b6d9481deb4a1f2de9104aa801267afed1ef3fb4d05c3ad5dd68d8004614ef3ef9921f995da84a7108d5a11c5277dce43f21a7c8abce3c5e925601be5d1e9b0b548a694655076ecee383aa10010347692ed84f3ef198431076c68e3c73a27df82464a87ad4dde7c78e3f2a4c8dc7f373765fbc0218d93e0fbb079a1cdc316ad78fe7065e966a2c7483a185ea3481f05b01592f289ca9e314f5529fd0382ef9bd58fc2465a4ce39eca9bbac06f3eae9599a76c7802854f225d01a12445776802b51e099ae7db5928c4bc1d55c8f4912ac14a951bc3d93507069ca1cb74c0c9e5b5067e4e335bb1338cdcf840e5e27a49e2974e8051705fc02505131f9c85437e1acce18f4e95d629f705857ae6083c26e01cd06c7b5a762c079c5f2d5a382ee91895d91d7d31b4f1a901c0f6485dcc8153e499bdc81a8f0148011aad00f4ff4d114035ae178e4859f9068bf266ef8dfe47f421dc04e007a874db6cc5d7d324d3fe917f7fa7c909d4bfba92008348a013d0ffe68221fb0bbf6f2a849eb8d35c7d85bb129013a66bc4da9cd51b0d92c20681e1cf6f55d0dceeced32f1dfde5c9d48d45da3094e610ed30a8ec9e5f4cfcbf50697bdef34406e4c7df7a9206ec08bb3fea4588d2add3a4405a2bfd6944900cfb6d3a1abd3ffed920725b32fb265c733069dd68a361663c15ff94853b3e2a403fb166e53e9946f51e07b16e1b0c1b992349302a55ae182385b20899c55e41c7a4e73f5d108333589b369a877bae0cbe10d05fb864aa06832781ff066937d008fff53456a997de4ada40dca8fb33537fb9c6a59e61240c6baf4d48a39b4ef3dc72516db08f4cdaaf7c9e7d93762ec9a953dde632e180e685f87e3368386fc642dcda74bcac39b8676f4271ba27172e30af85ae2380aa56ccac794468a4631e98cd172189400424628fa79e4d1535af8b2ef0483516a681cdaa6c2040e91677d1d2ca2b48d31f17b6c2347d7cfda704528ee0f66ef912601043338d4051c551f8987ee14cb6dfacfa5ddff5c3579e06591c91d271cd89fcb6c49899abee752f0755dbd273c2dff6f810af72aa2233d44bf72dc6a1d8b72723b63bc406485655e20c0b7fb5133996de75e1940e3102c50b24d47dcdfaa1bc443fcf0de6d3c725019f6459daf9abe66d588740b3100fb47e7cfa0beaef897656dfccdaaeacbdb49425bb7b005e8fb9fc7c015e5c39adee05f321cd00668e9f038f9971091ce0f0b594ecdc4204ecc31120df8b0c5881503619cf34e0727bcd86061e5703622d3d007319f1bf104bb2e1c579128256b4acb0949ba64ff6ebd407246aba7550917ffb9d8d49544fb9babd57c5c0688a6dde854f5797178686be0bce1d65d3bf37c4952f90f2ce28194c99e197b343fe56592b3db6d5e073aef7fc406f5198aa5a1570cdd959230e429fdf50c87e2ae38e76e5f4c2f247c91655fe569de5ce8270cef737cce169ef7602b1cf04cfd45d0dad049894ba4bf10a7e80415c8e5193b085a4055e316937da2affdc1cd507c37d65de4ca6adfabedb2c00c8590bb51318953c6fa532ebcbeb521b2fbb01ca94b2806a4255493d6cd95cd600314e6f640afb4d2423a69d61664ed34418bafdc20f48369217d6bdddbce34096e28064f0f6ddbb83b1c322b50ada3cfeecfd6f7e8f95c653d9a6ca241f44d6e5bd0feb83e044027426aa2aa6211b8cd382a249933113cc1dab002e76b6cc528153d34536bf48bcc2a65483a69600d876e512842a8b18c37d801bd33f8274479c0d3cbba9e739103888643be182aa58fa583af70638c5b5c43ae9032e460d6e98c6a0fa1c60b936ed2e4d16804eb9ca36622093ab4e7e098a55161f5ea16b0c96ab3dd532ff3e783a3c120bddfce05cab585168d71195f159e86d53ab64b946659e7f498a87bf62dd96d094f2a75293542dc44e872638ed9b29e3d659db797e7bc6a89073e7906218c7c031589fab939ddd6d7eed096acfe91f3426f458d5a3e31b3926e59ff287519d928d7aec2591a2719a7391cce1c2867d5bc6fc5814b37266a42e4a4e282936bb834f7c6b06f44259ceb26f91e5d091711f79fa816efec1f2c1437675055cf58de01837f8a14eabae53010be458132925296b3fcfc7e269a21d2e7917961b5d382994cffff8a9bf6ee2e85d4392dba3abdbb663a9f6d862aa4fcfa37ba1bf55294453cce33da4fa070dbf1114f9ba0cede5c363fe832f5b51ac002bea7024bd89870758930833a50243c20acf9b5c647ef4fd5732a2ecc0eec125a5d813acdc52404ef9cb451495951cbbd6a6d5735ca043f8dcdbd65a6735ea7eb600ebc662e69fbcd5c2652862ae3cb1f166dd3d9c9872abbff4432ec1d62ea4b74d05c4e81dd7e126b31ccdd281a8c8bce301f566e6e8e8ba2dbd45b43a178fee6dae86fa7025111cb7391c0fa9ccdd15ef3fc83d41dc90c51d3de50e3e12f0c013519753eaa9b4a3938a70c1c9c3d13db7a91509fc77c2f59490a665f1c7e0496f9b6ddf3f0be71ba32feb6556793b9de77c185e51ddb3cac7620a9c86244fd15e35f885437a6f41125a90aa9951ddc15c894dc847922189bd65de000b71305fc0e489bb0502e00fa2181dc718d689f1b7b15d7f6077a0b56251894ea0372e418d8d4580c28058a0e552338285e802870dd519d4d351eb227c04e9694001c297d6157498f31c73b97b061914d02e2e9af1f6c832b937a0b59711b90c59f556d4a2bb021a797a03e46734276dc3ed90bfb8ed24fafa5d73405021e808278ac019ea848dd94c620d190f555e42599367cacadeb461e2abf89d994f480224045bf668f14a14ff6fb85af7cac265cd28742a28bf9492c418f9a4307b331d55a7ede61fecfcab71b867edf3878eb1db9627fe3c73b1a7fb5eb1a7211a8704715c01f9ed67ac90f35170adad477e356a4449d60eaa10b9ef55539b3bf223da10554f120779da3be7873e08cc3ca3f50356368c94809b03e49eaa29015c0d91cf11d0c9928adb6fe4133700efb90f3c39fb0b5d63e35526e14e161ded1c20416ee98d26c48f6c3d487c09b820118d9e45e0ed4b45f440f1e98e78e9cc3770f5534305b250da9b068e31759d87cb842a3c063135f090dfe7538a661049b3faf9f43d880a6874cd2f9c5e97bd39a3812d532f1d4ec61f5714b675bed04d549b995b25d8f95a53eb1d35d618fac8e24627e4b11867eee8139c657e38aabb8ac086043f3655bbc05d04c5ded6af7e2b0483d9e8d65b60d5f39d4c46db61604ceb6067c9578961565b452faa125cdac81a98371c4bd2934e2edeb83ce2539368ae54fee61fd016beb450fa6dd4f9bea7095e4679052353adc023f57040d8399c90856be267bc7c10aea25f5cd6c0bfbc5079fd8478305e60b572b3b39234b6f249a56fb411cacbde7bdaffc5268c6fc34d38926dbf4ba1cbd3d3a3dc301b3cae17be3dca5d1ab0bff441af7870878f25144d9143876e3d05b8b6a93bdb154c997d3e2a6ca7ba2441c6131a929be1aa1a69304ecc25363503ae6b9fadb83fda1e1f6a3021624713b095850be4da4b16bcd437c4176b26702a1c78a96367c29d3f651a7c4db0e7154ef9609e3bf696f835dc33cd91d35a772eb2e660e5af67f1458f522b3aa311217ba4a9c3f9970afccef2d2fc091aac3c706e72d43b527757cc60141053345569fee5d53d0f35206ebbf762e90353939d95040fc7886b78e440c0b36c1a4c3a74b7fd64e79370a427514f51000f3bd9f67326fde3069f96cef3ffdd5ec3e323f0265d8f6791793634d73a56006c789b4c8c8eda171e2ebe93ce00042de0ece06eb38473d07d46b9140a4ebd16cb3a36692f1a36f059ddd7ed5780a63c5108afd3c5c7fd188f1db61023751a1d86811599d101359960f1059adfec972ab8b8bfef82f42d457cddb5c89044df9c49a06ec9ae36e2249b3461a4789ffdc7779d12db303e7fd1a872cf6dd37f688ae361da56b64fce20f0a8e06bcb0716094bf3fdde3b76b3128b82b9f26ad41e720923db19403072fb5052fb06b3ec90d2ee675b7fdac0be383384b9e0553d36fa05287cb3d48c4be7330aebf34c2519ee543b64a327b2a4d8a005eaff10b6170c69f5188050fedbc43451ed4e47fcb7dcbdc1a082a550d344ae6807394a3aeb8ecebff75fa334fe38c4f3582eec286d79d6fc4fb52ab53991cee267d320ab32ec9d1e95d4f726975dd41fbdea3d678b471ecedb10c7cc805a9c72cee4d58c0093e0c29176b97ecc92e57349950f4980263ce4d160a1e1c7780a9c5b57528a7ef3a8f9b80edeee17980ce41b0ab3c12018c1451723f5f6728788b55d56628a829b913f27790582ec8f7091fa9802354d8248b9b104b15c728df29e29037e0a2bfeafa5427afea83adf75c9246047c8acff28f84ae71f3af5332f351acf5682560a6423b8cd77662bec3e0508bd48697925ce26dee15a5f014dbee45b962a8ca19a1ac3f561ff6435fad4fd98f6c7a5374e517e57df88ddea55b43210fda01c3d033a0a7aaeaba065fe41e21cdb2063d7161eea37af28eac137827744b3ad8fa25c029e2f17dd71755eddf51ce2c400c821b09a0639cfdee06abe0cea533f23c33ec5f05a0d497995da57341f4ef49387c6eedc508eca56244e0e91ed63d53b71b852e99464e4c056c4a5e1d8c46e79890bdc4d54f54fcf0446551e0d2487a8bea60c3f098348fd000e78e4f1c189707837bd2e85f8f841f0f569781191c6db4b29fe3d2f1563ab0e4ffe0254080ada6e1c3452b16b70eb76f684268c31040c05f1901eaa4e746a21b3bf22b4ab2618492c5fab981c6d400d9e6d60d5c777b84f464b9c0596f1c4f5324de698588e3148e0f80b1b30205023ca4236e48440a250c73d8049f4c1347709c355707d7d31523d4b6a182eedeb795379c78e341e3ebe04fd58704aa39849008be332ef7c20a7fb9b94dab1e3ee38b4e23dbfaa42e34d7a42c100bb38879e8c336e92b46e1069f82068b09c20879b98b2251661f7cbdb6ad947b03408bea623ff227e2d1ebda27e54edaf31ab3d9ca907b901553e8818c7950580892437160f05734bd262deea0702fa9ab46586a331db8d41d83bc1f563afb7ef0371e75edb66814135e4ee9dec8d47bad1c2e2887d438611238520e294dbf57a1b2258f6daffe2f7b4846c233e2bf6dad6178e938d6e4f342698fa2941738d6a3b67c13ce79594f5a23dc1a88ebd3bc30b636aa12da3e59c4746d9a22e0e4c9e6e40ff64351a6f69b82fa5a02f5827c909b18d8218aea16d06510c7529f9241b200b86c988db9a27a2f89295767f648e83b2312ae870ce8ccd30e45a0e6b4463e246fc839f86270cfcfd63322e9a3970933159ac23f7cdd062014c5e09714ea7a6f5d22bfdea44ad61b238eaa5fea678513f42d0f1cb5ce4383d62bf7b532999709bf5861b0d80cd839cd450e07c7c2c28be380e2ef63c8ac26b67ab6555ec6e4df3dead344201501bc37267b6ab9b4b23d08d3408eee82397ec8297e804eed3dea2333fb240348a7c3414202349c5369ef674d7da373aede6e4a118c07a1257ab1c3a889a4db81f50157691adc5a58fd7668d78ce0f956f0d2b252b1cf9d537f9f7c5f406eebe3bbeb46fdef493a3180b3c31687ff4105d3b90d31e4328516c57efc33cfb93bc4eefcd9ba0ebbe3184978fe777c6d0edeb5e9a80aab7500cdf26a340;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc336c0bd35912d902fb8a0ce83741afc71dfa207891a9cce57cfb8d0bd14ec2f668b946f2987c5392ef1023bf87d00052bb8d688ade328482bb0742527507a5fc7bc9ecc83e9151c4f10af761d4a39050cb13ecff4c8151667ffae6f9bb110b1effaaff15253d54022e785070d9f4b0bb0ad546ac9503160d8c5fa5607300723655c74964ce35ac9f62a76a081bbfb55229fa5d415b4e27c76e4d562b325a9cab5e2924d583308f1834a5858a01f0524360fdd1a52d0c81dd836a3985d6734fe3e583e223ace32bbbff17cb4098f50d880644f3f47c0a70d6aa1d51e45b29ea7764398f1036681e9e302aa87011956071664b50c305edde3192fa160a69440d3f5406606f50ae451cf3781c78e2841174f95bce4029feac1c5f5c362db6a576c6bc64a3b50269afb1bcc78f5fdf53b0c83686b9fcb0d487496c6e560af61d74651366f50ad4be5590fc159f769c2cef65f0f0c8968d4e65b0086d7a43fb67067a6e23602b6cdad2f4039cb0204f9558927fc870471230bd143686c6c6648434feceee6e7944d9c857980341788b6409a9f381373f6bacb12aac3994da2587bfc0f05150476242d89cc4855b8a313fe08087a3654285e74d5a487fa03538c354083afe9b267df3c52ed02324ce042fcbb33a3d8037afcde31632a6fb7ec76a003e615c19d2d77994ac33e47144bf511beccab81f33cf12faa5983a7e1a42b5532ae78fdde19367268a434d0615c8eab3d16041b0905dfc9b06540b6b8f4432a59de52592c5a086cd4eff2329884172b24fc60c92bf1fd8415cee67eca19b92d55069241ef24828e87291a813e8921809524b707726f5a724a7e4dc562aaa4b442a4f48871c9ae2f667eed065390e8e6ce4e829e2d359abb4b4cf37a8883ecaa624556af25560473c1f7dd0e1bc3d4e8518ea6e6292063faf42452df624b938cbf6ea83da395550ea0b6c17b6cfa7ceb520556d32f86d00db809d83e6ca401587376c30a122d50921b503ab17e2a40e19b74e934bbbad52141ae9a488f7cb9f576e6b3adcf0e06fa88b54dd224ded7d7107df74ebc7f04ea160e4f5e3747a6efbfa4db02c427260097738cd2f0033a73b1cddf9690f73bfff37b5df11c70b11e2ed93008019aa9c4204db14871a452bb2cbd29c537ba75df74274fcccec975a17e2300a01ec6c3740a4ca80a30f9a4bb96d70cb4ec063d1d4b71f736870b6569183f2f6547607cbc3cf6b3667764c23d258c878392affdafa2004394508cedb7a28640ef87ebb05b2186c45d4caf8fa1c95f1172be2f01761e1462315ff86901cfb3157dec315a5c5d5efaf940f96a6ba53527cf63a1bcc1472c1d1addb50744d8b8d176036aec605b4cd2e74894902ad69f74fab304a4941781c6eb8fc10964623a3e6bdc7462fa1ec4b692270af8ac66b0f42764e320cc22810198713edb9b4289f56c5ba6b34c7c8a488e7d6c4c31a67083e42beb217bae6996b9487306b4de323c3cbf7ae5e271476c5d55cf1e53480570469a0bf80d3ceb39ff4b71db9a7209231d8c25f9f250ac789f84a077edf0b245a9ab068a3a3fa7b43b02a632e44e0a4bebaa2ade4a5881f88deff927c79602eac134f9e233007bcbf1947f6ed664e83ae14061c9f3976d5dfa1563f1b7cade7e8c0c5002a8618bdcfaee756cac9f7e448ad0a80433db20b6c579448a5c8e24241e6874e5e51c194298bafff637a7cc03a7e2323ebf3ab66e7c75114713d0f80c0e3d7bf4940cd712d560d71658ac16aa88dc78e046af2a0d2bd5ad83556878a3bf59d0e1ce3d8a52d28197ece613d6cf70aa2ee22ac29f5131a725312a4dee42cc8988e124fce3b34d1e6f072e073d106bfc1a146f84c6c349f9943582e6cdda67ec449fe6818205a9977a3a504748724bedb2aeade4a2057e6118a6ad46192870ec998e85ae6f38adfc3cfa0e76ea95380a16571c250202ffa046849c2c11c60fe78d573084bd8c4c7956b8713686feabdde59136574dc0b64a121d1609323abd6ea37d59bd1e78bd1e9c82b2266713580dede5c761a699a71adf19a2929b814252c19f1204a1c7dd7ca2191bd52eddc60782c28bf52fca1ad208f7fdf290a97fdde872675e894b7acfd6297f5dd25beb7ca1e94c3008999facf635f1223a0827250a59366ee5ff9c5f5b171db3f15b676ef88c3d558bcfd33b01fde22a8f818bce0ee7a4212ede230a8b96067f3e1c36e94e1f8a6db7551d01f71bd1f13aa3889e6188d9eebf2bbe6188b9ebf15c14b9f241e352a4127db334ce83d69fa5e3319462fdf22b5c0a69be008d5af7967a6cc04b5d1a21079aa0bd7a2436b2c49b91ba891e49c925130229f076effb9607426bb3ebc437ce60b96f391a36fa678008ef836956b4afd6714f3bb084dbc7e7bac84272211fc5bf6d45b027d108f6b163bb9dc88bfb5040ef6741967e508512baa4262db4700ebebfeb62e01ac3c6fc37b561dc993e5009bf0713d5dc681a8a001492b84459dbb1e3bee6b304d431a7217f4fd92df70f741c7b704f6f616cc1938dfa73859294597d01a9fb023df435b9a1695449fa6852df4f86bb976250e8a86f78b1492a5c6c5324977deeed78dff6d7b12035d0096c85638d171a0b87bc95abc8aa354955599f96d65da4bcde20616bc4641989c993d66689e8c468f839060112a6da9a3675bc784a2d2ec97b0ae815cd7234c322a3f2095560be39d5999ad19c7b7e49ecd3c2007c722e38ff4bf2b8c15ec8f39a6c63a9635de9ad2f966e940d9139bfd316132d2ce2496058a7fccd880e43afba890a5e725775d7c0d863e6807bf8ac94835c57925fa36ce5f2af0e4e184727b5284bd9ff3f209b3c530a1665b0f06ed34302bcee2bb023ecf401385ab9bb9fa21c8984235fc4fce4f78455695e00d7cbb5d9f58c2638bf2f4b4962c9c375a793063f3808dfb6621a548173b69e96b78920b66ef214f42394b8bfc2a4e661af7a4de8c301adfba6955c700b11977627b79a03730baa7df256219145fd91da748215ce175bbafa81c4658ba9057da4eb29102a01b98687b8c5b0fde60d1cc2054e3a441aa4f82b43350081c1e7f13931b40f12b48f19ee9e42894578384bd64ae416a4ac7d8640cfd7e0f84cdcbb724e617cd73ef84d8dc182d0b5dfa4a2bbb29a7933e5eaf9230da1f1df56ef37e5c1b295f29f65e66616a3404adb4f96038fdb8cd6d3da858a866a5d1776cddf83ab659d920814b999ac4a5dd1b5365a9d96275fb0bbfa3985c162e4a7bf2e54813d7ea2ddf004234c1fa39f2091b9615f0ceb5ab86d829e4c0332e60492bd7214af39121af30ce97f8b9505bf8af060151e2fab3f2632892e66fc04ca42ebde7f674fc78ef780b23c8be84ea7ad7d93974e10a6240e0ea0c0e166e4b596d028f6383c5e421f3cc6341b1d0a175ccf5e6a47921b4142a29557bf36df0f7fd8f5c8fe42a1661952d07b46b2bf934f9ef78dea3ca3acbf03d2a8079341cbdfe358b04d9a26412eb1a9d3f23545eeb62dc7678dd5fd676f450cbf761cbd652051ce201d0d9d1e39bfad0d207d5c8206dea4866b27e8c2532936eb3abc0647e59075ce436ca4842801d5100a57a62066e487fbe1768361cf004e7323daf00c3ef544e6c8a70688019ed2b7325e8d1d5efb8f6edc6299e108d55170e94664ee11b859ef2c4f3649e5beeea44303fbeb48fd0f5fac1c36309f9a93bb5f29bf931a1dbd3865e88fbb1c0add037c1fd50836425388a1c5e8c8730604676766ef735f01fbc5fd5d8807bc3397db4df49c31ee7383990497a7b21241404270a5820a177df1fcc57576cdf52a7accc404359c9469d0bed5811d5d614705312fcc4608ece21bbdf82817dbcacd6aeb0ef9d6918030c65f2c9093044c341785449a9863275ef0e06afb3ea8d4e08127b905405c9f5453839e168fbe67ed9e632afd207c7d1472c9c873f132cab655533946b91c855977f386bb8c6791cf8a725bd1cc1a8bb6697ef74671384aea63164c406789bbd3db38d27cd9191cdeb046493a87476863fbb0fffdc6b7a7af414164313f4addadeb3bf1b4281e56a2578cae5c8481be64c31045019eefed8417bb6125a24ef29a0408eb053397982ff820b1ba311e2a8ce309a1bbd12853f395a971a759b7227d3931873bb423ea3e879a5f899b64f26b5e6d462448f5a1266581dfcbb4743de952aecef392ce9858718f254e144215360fac84851e38f547b37cef97d8e38cadf4870a4d95a3613c662f17d09dfead826a5914c211c4ab7443800cc4704a92c6fd05cd997564b7d51c490ddea18973bc9f993a5f2ea2011f008e92cf6a02ef3f6ff13698efaa9fed58a7ccddb4bc5f993cd3289ef5933d233409ddea9247da24042ce52b5d8e068393fb319a9186e3e14c7273adbd57550d4616b4e4c011880adc15b265415d607e7565c433f699b3ea3162642a5e1037a1e893dc540a639495254162d03762133769a327f6bc463a9f9759c406a8eb66a20e3e48181778726c10248820f15d0de0caa71bb9026d948c8a5c6b755305bb9e6810b1bda36bae6b309672108411a628e0499b241dc8bf436f4029b5025142fb36fa1123db958ca7f1aa2e87cf8aa2832b2fc4797b9cef3880e4487b780cd5afaaa4cb4153e95fc957c6c5d004a0d0dd949aee6c3e18267bc761d92f2d71c77cd03c363d62524afd514f0a6330a5020796163d65994d9421dc88c21370a3285da0160ca1cb0d040f421e4b904f4ab4452c4e224637b266134976f4ce29147e6151fe576e3ce2ced9fd4171589466ab5ca4e8137abf35ec58b1791ae62e56e8c8b044d2ff5db74098e142a99a8358e617e8c95e8bb538ba6424f6d6f5dfdb78e4e6cce2d8ef8771feb62b5e0cb67f0d7de2f65322c9b0a7c3c202bafd6718b9371403bcb0cfc7513eef0eb3e2aad1b2b7a60ecb84e73009357d55f4a36e792967556124b81922afb960ed87ea8342b273cf83e45c689ffc69e679efc1518fc8e57cda3cedd8e0d912eaa6c4ed10343803808c30de3b50c51b551d828f0f3bb705ddbfed8b568870a1f5c20015b06b186fd0f3182d7e89668fd83b93a426766707ab5f3641bf1542bc12d2cd3ccd526f6830ce2e718d60a45d25d59beb2a5372625941cf8f0b53e2730d158ecba337b5a4255078f1e5bf526dc947d9dd45154e4314cdc8afa93cf79acf0a331f09cd150736d903de3b03634310ba5304a38ed0269c1bec8c6ce3faf2342eceb7722bc36b3d373b55f1609fc3c5a30ddbb034d9170e0f728c75e10d297df3edd6a3e4625b05170d029ed20fcfb48057a85ee1ae1b7c2b551a51088f229c5204336d2fe4f97def5c03e249b809af353df3808aa38e9c22da31f4890fad95bbd3a005fe4f96e1e1ed8244d1d7407196ba420e8631ab397a0e06c08829cb89e5c50d7a322a1eb5b303afedad73939b40e1c12d1ee68e8bb7a0429f64ff2b638e1778aaca772426ff40e7071ee5667384cf52b57ffde01300b6f93657f0c29351c0321181046a2f65e0c22f9c1259eeb7b405b8f396db0dcccafc9a04358f60b1ac43b1228ee9dc3806f291c1904d99e6128b49f9635906e8adc063be5827df714cb9aec0d2281d3ba8c2454574324a57144dfb44aec8eada55c336588584ee5c765ac3219c900f2d02e0b2800521859ad48114fa018eb2b757c7686d3b6761ae8ca82df117b56c8e4e62e690073f59c07a9dfe66fb312a5471b28eae8d3e3f6dc3c34b6cbbd39a281982485d090b3c921eb6cc916f970b95d77c2e389f709875bf96cd8d30e03b18f7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h8099953a6fc04de8fb54cb151f370a47fbcec2e9c5429e27b0082e734ad5aa11f16fc1f225f4277f35046ef809097c5b27da8a3817c7f6d3e81210d9c57d3c3360fc01dc522de2be8ac7f1d2a31ca13621148e6cfd8cfbc4b4ed9d80eff884647f1db5768069fb5b6d770d84cdf54c1aa76c05b9ee559f7c1dc10b57902d073e185617fb63416ba78cae9c17f8b34caf66b65e18f01cb87860b91944c573b15bd6df5a1c47e725e59f15f9c085366eeb1f43df93b43b17a7cf55af09073d6db63804bcd33e70703978057b70ad666d1ce69cd9eca5212c2b012ace187424bb4bf5a65d694d107da9f3fe64c6717c5e3aa29772ab4bbef359cb31c3ceaa4b7a4d005962331ea21416173718684f562da5af5e6612ecd22ebeab2832f843f2b07a70c9ed770f4a7dfbfd668cc2a84423a56ea71c1edd6c9d83b01e438191f4b7ac00c6ab6cd8606763a52ac2d6c2829319aec3cbcb005c95c46af80030cfcab1aaa26452461c6b1408e1b0f3cce928a86b2e0f1f86048ebb3101e271f2f118a0cf8a5fbb1553ebeae8b90a5d273b43a097aa03bdb66fa876c92b301226dd5055504ca5795ac79ddf4c4903b65b3caf4512dc28cdb5fe1c035b6ea64aef795335f5195293607e7b14cc09c09f2ba3706e5aee1e945efce97b76c055aef17acc77c79f2c91c9839aa4f9643db044a30fc01759729c0511474b522f961b3ef2b7a1ee83b818713cf088687214215b680a1f9a84f4711aff7ddfe5dd3abe91a7a5c1d4ac70289d178cceee3bf82377db14bbee65e7ea2656d5593f70b6f7488812bf44b6f7e4a01b1f481c88b8f6bd202e1326ce3c82dcf221babaa79837690766469efa070eef74010e003637d02977f2f697775d3733072cddab06762e2d3f0b7262ca37d25cedfd4729a40710fe115b6de7d583d9f532e71d78211751d68befcd827061d7521eb1023624af88a61af10ec7f899179a004a9a5679c379a01662a6bac711281e34c18407aac250cf963ba36471942cac7251804c3d86b5d04ca564407b7f0caa0893973fb3a8701cf429574c95668b4428f927302f7d017afb56dd091d0ae11acd699530d2ac3eb5c4b2336f43fe70364f44b5c39eb0f1df4137bb1faf8f05b99077fe6ab315f3c27ffa292823d63e902242b00db538684b897568ff46e3b5612e21b917a93a1ebe512b9318a41afc36c01313fd790449494564bfd4d40e6d73fb1fb39e956cffc5dc7ebf5e563d1f0a4e47e4f8f6eccf56614b5f809e8c00c95ad43eaa8f9747266232abb6b9a618e535f03f3272401a1ac2181a52bf00eeac1fa8aeb5805a3aba93ab271f285fb4b9c312cd112f02524002bdcaa8c2ed34d73eddf423ff8eb1bc57407bcb640a8ce6b5cad918854013bc3503cde693f3e8e90ea694e9428d2f96564ee7cd4375e9562fb8707f6fea0ab16f8fe4f16f9189d5e11b8f2e5ca978ce9ae6ba78fba9dd38930310409e0a678e97a67fb1f0cd155163e183aaeb06be6b8aeebe4f95596e55d23a303b9d135de1df29379b089a18bce80174ea82daff63d8811f8c723b3e5f2fa2d4f32cbb361f6a9db3f1b5905ae606f7210309c9bbe33ed80d9b71df0be3c74dfc954cf842df195fbda5c1f4ea673c37751f41716794efaf86465c75210a5170145c058d224acd99eda51252f1676b07df57ff7f22c88e083884ddb11f4dc2d34836ff1e36b8f364b124173059ac7e409ac63b8613ee945f2974a45e7a247525ba745efe15a63a3976d818916e2e487d3bbe7c189b13ccc34dac26814be8f629db42b0882b63cfc24bd5a6e552c27966f6fa4f49ffc6c27b1dfad46b4ace817ead898e4baf5590e3af7fcb23c9290d98eaf04937e3aa026d3103e341ff1aee186aa7798ff3e5372ee55f6c72481432d02c4c1e97cb1101faffe306d7f57b98a5259bcca39bd6f1d484b5ba2ad19eb24f4bef125b8551d601a4765c317c53de3c665dba86ffc60593b46906df70d07a131a1ca8413c252ce1d0230b6582a9c5d6e4a03159e4d8931f3e3ae9375781afecb3dedbe20020d2834a083eecff884637e5e811a4728bd0c407f6181fa202204fd35cd48382d2ff48cde00fe978bd7e09cc57612aa9b815893bbf72ea32f5dc9da4aef879ba6896393f6dc86dd2e2217ffebf6cd758059c2e989059db3572d90a6e89020bb2b39339e9a39b9cfbc8ef81869416f2db644dd8a9d613108a2b606c40cff91a2e3f98fe9e6c3d86281243eef757234661654e28966c162dcb42c0566466252e05ac7fcce9f6036150dc180c06d4206b1e70456aba357dd34457e7b08c20bb48aab087ef79c280ac2ffc110c6b325465c587b669379bc186629cfb94626db6ffe748ea6515c2bce89b7f0ee37c1ed531e16858908269a526ba06a692df5346caaa780803d50f06f81a959cc7e1802f41db8eb0af6d3a24990066fe04e7fac5135f252d81508c5b565488dc404ce6309017f9a414ab1b2f556938a43b21fffc9b9a6a7b7ba6fb6b92f5f3286b25eda05bf40397c8fb7b89e018f75b57cea398444675fa08b979506a76952e33e18f28ad08ddb65644c76475b6668c355a98ba1087af2ac3b0a71e2b9314a7bca033791bf000b410501fc1388ea7f3767a210e4152714bdf8462e183cd985f164208d2d4f7bf05b0ee7bdd429e1241e1218c954a66b328c1412455b9ba1c3c64d532da0f2c5e6b7c24b62b910cb4e4a80bd243e95a5e3b27a29611bcad625e1c910843bdecea3577fceaadd2f309d0e0aab2fe1c75a79411c0c26dee465ca0630eacd7cacb5a95fda198e25d60767d2730270833c3b8babd5879f34ee4a075362e202ac8a9279e2718ac035b93fb0890fb7e744ed5792d52ac541e4ef6a87b9b32072abc18947e9b68f5cc265c3cc4d167b53ea82a547fefaa0ce89af01043c2828590ee176331b5a246587d4bdddbad9be8c4bfc5ea4ea379f2d0b5b0c2a423915a34130fc46f7d0d4c6fb9af69d334aa77fc0abb469acd63e980e4bd9a5ddbb5634bb7356dae17ff19a65053666bf544847c6f072c927826f2dd850b309abb009d3c63bc0abf761018930948c656d8e89a31af4ca5b816f14b4e0df0f4192e1341f8a737636390d03e04b1b976bccee718389c16270935003ec188c8c9ba4c62fcc1d71585e2ca4f9e6a8a47ef2f864d727f9417cadc36c2263e3ac7f0da94ebf5b4dcc8dbd5d700aabb28e0661c3710db70014aa700fea529a864cb43c55cacfe320c67b2e6e3d1f6cec2b5010fdfe7086be4b82901a21dab0d0e8d7cf86e834274a7b228390a21eecffd82023ebb372d62259667a5a8d7668db2ca57d6f734427640a1481122cb0f4bde2b6c03360c5d0870f12073fada84781e40396baedb26c8965ef0fd81e3172e235e16f4f25e90b0ab48bb3c0cf765adac18dbce82177f14c354cce39def0fa7109379a45d5705cdece26ecce9c97ac60984540e2c34f4d8a2b510c0d976a5e639a3e7812d018a21b8892db9d7bc057976f804e5bc48ef16c8209f9c06f2664043c9227b8819f06da6857b436f7d5ed7f2c0f147599ebf396bbb6605fddcea6bf39bb2e4769cf5c49c2e03e57453f1e8129c9b8ede492999cb5011a190b78226865e01576f2ae638c8d92556da619ddf6eef9d0c3c3ce2d239ace1710f459d70bc19ae4fe0f0522e63cef0639f3725c335b445668d9e1132c8c517e54dc31fc073f154aa883cfc138658c7edfad99b31963f628cd7275cd17ca4374e5f1407df7b99f94b896ead5209be856d91f354c36f48aa01849c1ef96ef101161cf254a5b523883964528400ef7ff650039628a784e434a952d79df45b5aa9f79891bd6d8ba8b9ce3b504c11ff1a5e650f5388847afe44e3083ee7c24c179740515e22c609daccf31096b2eeb199162ebc148a6b5edb0c71b58f3dddec257036bee00cbd843a4c6d5ea459f702cd7534bce89b7466b95e657b54e424173d880e6944d2420cad2bd88576475d183408cd98a327f2282617122d82c4d6a43139f27acd387c9aa5978e1e994d246043d490f3d46693f68e224f1738a6232ff9e0c6e97066298681fd1c4f026e06a07d8cc6900060ac9506a43e4fe45d545ae3e22a3e9d44afd4d129415b822f5add18ec846ead4f062bbf13be7405d22cf1ec3faa8da6c672e842a9dc125bfbdbb52b3ff79ec3c5ceb6a432b9b0c55e72fdc4f261c05eb9952b0afcd0f36c3182c112e9f0879a9da66d046dce0c531e7accb85ea6005fbf2e0fe5c5698c0a6d6fa411c50b227e4292700f7da532cb902210ac6c1b8ad4bbaea325d28835b1c82dd9c5df048e5006306aec20ede2c2109eb4fbea5a22f1fcd322c7f2792510cc06bbf53b81a17f647ef7f7407041861bf015c27b05c12d5920711ff820ee6f843a494e3037bd2639d4b512cdf4d02bcb1df0f9682cbb68509ddbecb254899c271c7081c03e991bd320815e753fc1f45d7d951847e344bfcc2dfed7903090d15bcedb010cdf13464c8f4a0ad35dbd2119a82184b58c3e24b03e52bcc95e07b3ff1051dc3f6461777ce2ed8f45d279e35865ecc65fe61f5c3cc5b28cf721cbaf7c8529f5d3ca560abf716b228971c6e9106f38e98ec8d5a8237024d8418b028085bc5352e7fa6d2eb0d88ec499f8b20e145f4397c6e21ada298757f37553035fb597f128f381e807b1757ba6e6181804f8f43c4dac80d2df687f2bfe43dffce1ed98caee089739239cb8f60531b09be3c3e43666912ed2aa20075cc55b8e2ea15d7201ec319f9f76ccd9a18da722f28d976db2a40faaf68aaa2afc8f92eeb6971360babbac0121afe59558561380af061a4df92493d2a3b24bccfab19ed4a523c93b82a583e5734623554a5a14b5cd2b8e3327aa3ddac86b4c73a591155ff6f8c8d62c77bb48d697d5ed4c5830634c06e0cae605082b54b5e23f5847acfea954b7327ea4b54b82c40526a80b030a2ab5e2a661f2f968078eda995503bced71f8af013681cf3b9cca25950704bc391cbb575b5bce232760c1a90c4446d2fbc2e2c3f241a83dd1a7c3b22cccab8053abbf6c23e21210274359449664219d147b2c7c178590bd9ded55bd74d4755bb2437d7dd8fa356131016d45aa84789089cdb08dc0c1401d963a9d226388dd3aa8453df9159040465bd8612e9e3d67c8a98fd9134725f43347e35984359036edc92cc61a7145c850df4b2084f84e0cf982fca222ad8821cb387c0b65d7ae54cdf6a06317a37bcbbe33d986824b9ca2307dcc406cc2087679ac447d7d9b55ec6b19795e9684ba78cdefcfb61e4b6e380fd217a9e2edbd994985621a5e0e881624c6bedc4e0003e8e597ca1d99235347644488fb155aa887caf1c06342632d42f6b89e3ec144baf7a1f3de2ee87f3ebc94fc097536ee248a6635f544a6af0b9b19c9600d5394e82562f1ed50387b5e47c13ce1c4e8db180b0fed4f61690f1c49e663414e8f2480b5ebe5e14d740333ac85b4534cf1c5a0bdce6aaf8c8926da4f67b0781730c0268fadc423316b43e0dc977275aa5bbf8197cd07283f5ce772598cd6f1a48c324e8580c3cc2e53dbb68cd9333db3b89c98a2f825b9478c4236b3798e46a770b8c21fda65d75ca8f7f93e3f6d03be0fe2245477778992b6a557a5d5b9cc63ff657f5ce981ddd51f0a48baea4b57fb8ebbf7a0cc01dac771efaa4272ed4cd836e40bec12955d26e9d9328d52f27a072c6d301fffc15cc605a938b46edfcce8e94e2e84447678058922feb5b24ed659797d3c6491e17c35522a9e6f97e3710d8952c9626d66b0a60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'he22eb7fd328698578c4357ae45a82d0465757efc6be28a0b19269946e5d2602ed26beda75cff8e9629f11c741419c051c8a8e30ed2a5a2f4d32c12c75d530eccf6c9ebc4e0c480a87ce71dc966f148b3d5182986042109ace2f80c238b214054ea7d7be7a3cd43f8d1a1329e9360970eed6af2d8ab0f28c629ef92807fc32b3c745af918974a6135c89d3204f942a7adefa401a13f9a8fb099bd285b4dc25bfbb174da1471eed83f1cf00de5b906f91f427d24702ca26edf11275a4ba96ecd6ec927528babd86971b5071757d8f3ceff9defcaa5ab5d30aa6d2b636de0d10f314f71f0f0d8c583f818aa4ec27bb731bb8cdf5dd74ce08c8d1d06e62239f7a847ef2ca6ed3e7b0e6347f09c209d422ecaf615a1c9cdaafb25d3588e0559e4ad9a56714f48a259fc25415e497008d0acdb1ba7ef36367af4751d8a0d9a65f2ac4f347ec9da9e41bd43205b6f38c802b79f7767163d7515756a36d22b2e89c205e56b47d4e07cbccb25bd1d730c5253039348e46d3b6f401959c9b778a3f7f1fcde4a230cd2e38819ac7d8732d8ebbc4482fc65bf8a51d7fb5a207ac8bc93058760fa797c2803f72a55104022932c9cf771bb82373724426655af4764333bf111c03bf7cd2ebfa03c2a8c45202b3a78c714c400f6af81352a553a782c2b6266f59150041e7ab82523d0e814689f67b96cdac8bf9171ada2065d5db9e282b5b8ca2e521e811127d91e9581f7be5914ff58e245fbb0c1bbc77bcb722eb70b9f46de620c9a440b0b0adb7531e48c82df49daf5b1672175b3ad31c8ce091dd3cf15c168da7565bc63d4711d07805240e3f96b09764dd943412b54c2e8f9055332ef127b7bfdd5148a886f226761f7c52984eef985663098b2fe983b7d3357724c1b04278827a52c74981c52dd7120dd9db93e1109a253ac730bea82f67bbe9f2bf7b0b4a8afd755b718ed57f6342b66db6e7977cda9a05fe3a78bdd580f3f74f59a1e53cfb003b50af9878445b2772e60a1ee0ab8bb57384b9805f9f8fe2d20db63ffa7837b3209339e825cb0a283d6f4f3e06190441f27377594521f0cbc0573b4e197cc892123e0953234d814b056d709a60f03e973af7e140161d5db0e748a04c7ed92119bdbc754eaae0a2aa21584a8c7dda8143e973767a943a0de56a34fb9af92e0cce6badae476dda1340b74da54c572d83c99db07210fe563c25f6f6a33304c6130d15f5525ce366b688a4aa8ec300d0eec25e00f6e353fd3308aeba260e1e61e7a039f26b94df8f4f4c2d85b18a42f866532fd297390d9a18bb3e9a4e8102f82c5e9b8c117743d26fc02aa5413cf6514bf1aa58e9f61538600f0694ba01a9be76804f86ddad7c12e2e51cc7f28b725a95f952d1c4cca61266d9d9fc3a4c522acac7f1c8f63a66512980e869e9bbeca2dac823ad887f6bdd6ab6c0bd664e5f031a0322e715a81216556ca7f384482a1b7452debebc7a7c8b33e27a35ca1bbb40496df66cbe6859d96377144e38959c01417cabc11d013bbb34b2596a2c72ef8b98189830fea6d8a812fefe91b10e91fdfe95d484fe9ca390c97e6903dcdd078dfb8d2b4d30f8a76e6b5773ab72898a797ac5cdb84838e50e9e538f699851cd701b3facf8f8959faa1d556fd5c1b4bf3b17c1a1cb280a2acb191094d88044e731acb4667dd8ce33acf17bd43a778f5f7d73e6cddaee58cbf642def49938b97844ef9eded5edd96e3206f6e35095b08ad18e22570ee42dcb457d129276af95748b8d5f0f6ba7db0c904bf1576eb75777753c4ea0d93873a6194285a551b4f06f1a286eac17d00ce6a236636023e52da7fce3e7fc5c6b8847ed53885b3d8539574ab6680a2112fde4a09164df3de3ae2b815882739a4341853fc3ba18a714cd6ce055f63704f76bfdd3a3cd23ec3413ba5ae45fcb647bd44d315a625e82ab65e42dba56466613eaca18cf691e61c6f274ad7814ce5186d0374e903fdd6e95be2dbff115ce9abcf4e27163e774eca29b289418029b8dadd0afa2456d9a1f28fa003c77a734f8d2d5a7839eb79ff12d8952ff3d863f43aee9bb00b35ab32e941f8e4a5c2e8042d10d44769c94b5677dda6c90b48590c5778701464fd3926d25fcd858985c748d052e2754f66b153006d2b37121d0537e4a0e03cb11eac6fbf39c4bb134a5e154a09577e8e86ec4644e325b4c6a5b9f0823fa378cc524fcd39c15c6e32f6e0625231b100ebe8756eb6fa1171dd04a54610d824f7b33e0d8692d31466b15067f529659c80fd79804252f1ecfaec982980b05b9e2d1a74fbc3ff81afc2952189266608445501ff0463a802b07fdd7750ac24bbd3258ad32a314247e7213c27f2f61bc16c6dceabb6b015a3e6e1c509ca561f8e78a9cefccc6119cf16371d73e76ace73ed6deffa3b0a554e10b9f5676b8d642f7240cdd548a8127a311b9987570437118f19082d0053dcbe9d8abb4e829abee7525b7f8a580b50e0f347ff8a12c77ff74bf6e03738d4cee81e24a535bc517a19e9c6a379967b20d024a3d9ae1c65a9549ea546141b22308cf7d7ac6ca89adb13d774e8d567eff6c00d1937203fac121f7dc6f2a56a03b89f9691caa70e9d0e5478b95b7a0c9b784301f75b0ec95a57b1708897dac4f315eb766d0c6cd215f85f4b2407700f809bf8007e832a25079b1f68554a6626c3cd3fe93ce0c8984d470c73ed7767909d7b8db957243ffc7918bd2ddc5402d4ff06012b9d71c0e7b4d0a907c2f2b2fa6cb790dafb01c2e7d888a08b7fee2a9589a213b762526497673ef723ff77729ef6c7d6950e760a8cd04feecfbffdd8a20a8e3c1de01fc767b809d1dca1764a271e179816fa043a33796081a605e13e9156c823a074d5bd89c39da7c759bc51aa102f05295a9571421253d16e2f16c041f13ca5af601162dc10cce9a7b2848dc07536e6f4e00f58084c8b29f9363881de97bbd7a264b291435c7440495ffc7e08526d3fae2d0710c2f2e0e41e13dc387c6c54b01a71566e92d013e04d99218019cd07faa41bf5d761142db532eb8d97bbc18bed16d78da92972fcaa30d843523f2c2be6ec0d342a842d9fcaa71c860adeed446bb59828438c424c5a151083f907584d3d91c977aaa46bef18d30f0cbf4a0f8777e9d05fd2048783212d29bc0ff2e216bfed5afce140537c46dfbc62bdc2b9ce98fe5646e79d484855165bcb6d88fdb2eda6da27e314d3273c0b24219fb0de40b244ef4f3b751edfc7638e340e334db30f821a063f4bd101ff6cb216b150e415a7bb251e612adad6ea3d0ae6831b07c18d23fb2872e3a9660897af926b0d64c94cd8d8cf7e9caddda65edffbb5bc561c8c0121deed54f5600a109a1457c70452e77a9ddda572ffaac445797a9b35b9d79ccdadc3464254ebfe85e53d72caaca2594346cea4ab4fb2c548f41f68ab1ff4ebe737b12e2d4b1fe9c270161e4a8bc87fa53102d6efe841c55a56a779e5cdcea49d5cb7ff2f6d968041163026da131d57205beb3277a506abb5a5d8c0bd7e6386785eabd1b7518d2c27af6b14571c5ad9784c08004bf4e6f17cd3d12538c4841b1cad7be0d2ad12d455ccd48fc5cdfb643c640125adb75ce49add4834ce32262aedb839b0622ba5f6576ac4b3303ae4c7602761dcb25162a039fbfc4e566b719dbc4f160af8a4bfe0aa3f45c2558dc59269336d1fc3537e329c94f9aa7034f14257ad4f71a0f451bf345baa8e7d133bb890552e6b45223bc72c51251b10d15961d38e4c3e7df52d46237da4918f913016cb4923079ce9a35f59207e205da66fa79cdb8f82c08a716d8af1bb9e660bf0e4081231da322b995f39735daa76cf83812ef03b5bee24f39c0845225c0a25a90593fe9ad0fe987f91d2124f071024c8ede29d4a34c7700047b4a27f407537e64de3ef687af2b87635298a7c02944b437c0736c3ec69aa82641ec8c266a84280c4acc298b9f2cc6554c51ed4e70a82f801987c994e2d76146d0f8e283c530596ddd88069e99f234033a915cf21ffc2a94c55761365c026debaf938813dcb6d9072fadd1fb68c2c1ac8b2691ad780c66533bf2ef1ff85e58da3fa3b3ffa614c6fce2f94dc818e1a708f6976d0d17f9b3164c04aae7c49f87cc70a19c77c26fa8024af8ee22c40ceaae66cefac47a50b1298547886b8aaf604e6afb43c535683c9da37640815c3b9ebf0aed848a6fe8f145f1850217039655b36c8a664a0bd7fd26a903c2889ed01daf12ccc537e5d4f05ea3b5068187c70f60ef3c3066c915a97b5a7c045a015bfc622c47c6f5d35bbee764567f16100b3cc10e8e4e6570bb7d215333476ae15167ce6cc0fe14576c21e482fbf6e1a4dea9a6d43dd51361910bf12964097ad472856dcac3de7790b4a54c3973f987e8e7f563af21ddb404f31858f640b2838769b0122d94dfdde2fe8ad65658aa540f198813c19316bf073b0882f9c2db1740263e02c7c113dc7bd4a939cf5178b2a15e658b250f9f614814f9757019a96a8a69317bfd0b34e1f82d5744d16ac9f8b90dab8ec1c5bdc113a6e20a289536a64fe6875532b565e180dd29bff9f2e51ad8c7e1921ffb124597a27e041239d3c90b7c477a207ccc14ea012eade32b4b5994e6cf36e347bfb4c75f5faac6908bcb9008a3c00d4740d8550d0b71f69adc21a634a35ec29c022b118791389b6dfee5beb68fc670e8b3fea3020488cd27b8d1a318ea17cce6876977fb9b2c1f5f57a6a508ae59ded5c5ce4da0bdfbe946785b65e2ac9214efb33dd5650b624f0907a6daeddff4a79fdec35e53e47aefc931b2dda65a4bda717877d4c384c117e8d3b573e1728b0662aac97acc9654ac12c811c985e89fc7b0d1f24c492b593a72c74fbce65309b6cbdbf70ec232a754465f9a43c9a03962e0ddbe02b0c9711ecb13753a72b8d0067feb3b2dd5c6484263b9f97cdf32846d00d67b0193d01015f9922edea7c29e9df4cdb39e4f197d8d6408ac2dcd605cd0276b54baaa1fcf813e6470d9673327490f8ef7f4673e02df9d3628988044ec98ab702cbcc2383e0b4fdcf2d27f1ec5f9196cd08d7ba3ec0d73ae1929d16e6c98b4fa9943059446b2b55f8303a778a2c05ab03d0fe513df7a022c7e8ac49d3d34a3b471e9894ef6bc41eac5ce2f9e648993aae9bc65b83951ca31ee713987209c88282cb7875a82faebe9a40dcafeb8596ca7808451aca8a89396d3c2e1e679486649e6d91d2d1279ca9fc79a4ec108fccf3a207d8892efde3a351bc83518d43d55c6de47fd53e0e48ca44dba63d90bb9c16732c87fd6328c586d8f354a0ea534550d67ca33bc4ff6a3cf36a5387a3d6850563c44c78a31b641131ceda02e484119b8aab0f30634f4d4b2e07a130e0b7db5629f99efef8e7eb473f5e8c20d25b00aa46f85391ecc6677ef0c972ca73956a25977c0fc99f292be59ad21656da1dfcf845fba0d80ca19836012e03656e1a35d31a92ef9a9b76624560e2e5576d47761984afe5063ff21b57f270137f9817ab32fb11644e87a97a28021e012ad15831b433928abf03dd776430e03c5a3634a93efc546c3b15e42c5ef5943375b2fbc0cb66981d636eb8a92f9b1468dd12cda57d76ac3de1cf3f3d6f5abb3205f7d5cbbf6c0d9ac0f52e89f1dde6d2e7ea76e488048bf974ff615b2abecdd22f5bcdd06d9974239c5d7199a799bae5d4b14f660495e7948b15549494b8b8397f5d83dce05acbfc8cd98db0a9a141cb1b602ac3d4b6cb25baf8749bacdd40e40846de9e924ec17db285ce1f91e1372204548c77790924735f354fff77;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb51953fb44d1e3cc131c86d464defacdd6376809c17429bf60aec7f50b1ebde32707683e5fb805e6d702a46397dbbe7d605f5cd8b9b66aa2261fdd8d304bada28436d9f5ae0edb5cf69974350ca7e3170a2c8c33563d5242e619c7c4cfb6a1c390e13780f871b0312da43aecd80ea70af846ad48ce7b402357a7f38f7c0a52b039374b04ab0f65a2dce8e802f934d14f67d8db3e81137a1cabf54913fbb8af1e8988926239f703774d2613de4a4cdcd51467dabbc7ea4378376379ecf51e84858f6dd47bdd9910fa2f1d29f11425f597b97128789db8fc7a3389f386f32ea43c5f203337674c5c1e431412f403521c7be5fd94f43467dadfe7eb1086557f2d3386ac27113c6f64639c5ff62fba1f6307f3244edbdee45cd661377dfef99f6776c5b9899b22d07e6f1275570f11e6f5a20d2a8236f2b7f400e77afec8f7657a54a43d73dcc95b442c2af84f8f9477ced5dfa7d78503b01cd5725d7883b91480fe7b0795238af5ef3ca052f7b0ece754fbe4fdddb5d03ef614a09acf8dd0ca38c09b8aaf4f4282e953f275788d4e593be46bf72a0fb1db75592bc2e597374b425df18f78b02c53de74fe26b029ac73d2091d6f277f5ee8fb8de8964c086951396ac8690cc372a6e8fe5ffb3bc37b69830529c633626432355937cad088ec819445266f7ec03733ce2e1327233fc3f79c25d4b78e2ee1493ad3015285b586aca435d2ef480d6ee8572ee8908c1e307ba225933cca36b6895628c9b0978b132f15a179124916f4b5acb1a6668f31fd8ee7ae26e3fac554865ff7c846fc74ff57296369388d7b9a76c204d5303e94d22b520467175fba485177a036e9e1316d889247facbca76411956172e05b9f79bc249112aad51c720999dd2be209baae882b3f625bc9c0551bf8547c19994ef9bfa5f216f2f8763ae8328e7d0cfbc7f851979a6c5de4a462e3d4cb22a7a4d2bb0b9ccfb9a8f019bcf286dccec8d7a9369c2f78480095d06bbbd8fa946a201cc173c4c7b1dbbbd7076e69437cdfc98cfc4e04bbbbe43659b8700236401bb772f1048724c54366b05f5a4688b397be0a1d6d83230db0a4abb0bdd55ffc8cf3cffa883a2eb0f9ab9701736c12feef6f862974126cb32d7432effe7707be6ef3781b5141334e53ac0e3cd1c80d2cab07374b60aca0d12df1a90c5752a80ab34823cfc06a294b5b5e64a2629ffc2abde5218cbbede84a90df493b91c38009164db09ce10cddc46491e9e46833b5c4df21e2c8684be0e72dcdd2f47d4aa38a984c5e9cee252b493a2e6fb210bf6b0762d396e342954607c21531f2edbbe5dde6d560e6229141d63cb3e7fca2673942f0a8a7f406b163109f7cb8f2f30138cc377e552c92066a4acaf22103edba298a99e9ec5ee4333e8a70b94020c9c495e467dfd319633335dd2a7e5b9b1a1d9784ba54ccc31266aef94c81b8835d95aa077de063722dcf2db9e072ba383475b08d04d8400e9abe876a03ae0e321c925e57e3599d7b1f7651cf92596447107cbb6723bea90fd71bad8315af5b884a979adf5a14d4513025ac3d5b6f9e6c5bfea2ccb0129e409145d5d9ee8078727bf927f9230d25f259b43f2ce0d3101f975333471d04ac5cec9a71b90f33bf6276175caa7c34dbe12968c4e094b7b9e8de433c63d9c76901d4f7ccc11715dfba279a00565bdddc6439c1a11c715cefcfe1dda169c7049dbd95af904fdbf66681eb473dd1ceb58e159bf104be08792f103ca01afaab4d6db7c036df94b8165319d478e6462c689d27a06614dc8150fe973184dba6e107066ae1e702a97803621e81106eb9cfd175996804ae5c8ab61187e6ed96a9619ab2c22278974e245708d7c7bc5608f669de0cd047b4f68022f82495a4ef91e1d12960ce82cd9eae94366e880483511a1a5822aaa26d86a585ce6e1da6a6d9ace3fdd8bad279208592a1d767867c1d633998aece6f730cdbb78c50fb5ee9129584f8e881142e46297223d0fdf2ebd6ff9c1e2087fccaa769419258df99a5ac37a65abfc3c1d38c8c61137b97ac6c2243413fd5573abc625901430671b32f77815025eae49c41f37097914e88c1d834c208b58a20894082069686c0dd340edfc35c105a2446fa9c2355fb6952838662dce4608b769bc89096ac06f5733f2c88bc93bfa9e710075afb822f2336330b5a061617b16a3898039dbe06023556fc01c76e655bc99194f7661ba9935f20e9bea3c30bb19756fb1f97f5386a12fa2c80071a68f70bab9ab603e992d7710970634dac4bc4fc55eb359b83361f5f5e49afa4a0b37a212af18ed10704a138bbc2789e7c769bed09bcc8d895695768d4cc808ffb0452eda1128480ccd040ce620b5442fe10e17394350320431b9d7aa98c4a6d6ececf72c26c10b023b6a676522c31d879ee7ca9dec4fceeee4d16e277264edf4a1a449582b6cb8cf0f268ddb9cfb9bb3e55196d34e9b94c64bea94ca9e914b5804fa14aa783151cfbefe1b813fae984764812ed7369274c41fc978c365b0b2821a264f6c728791afb749c54f705ad7e459b993526dd671a805ec0d4cc97f32d27fb0f8cbb62aacf38d392904689bacffe5ae8a3c84b40cf1b1789324c5d005f7d34af470c77bb6b6ea8f909e8363296049c0641a9281c17e52ed9bbe01bda3d1cd1c79ac0ea78be7be1f2958e5206cd831ca19b957129a717c680a273c792448febf686babd2e5f234ab791b17cf2177f6e683a25e70ddf5b9eda24e4555834acc58c984e4e535fce77d84f0db4b8bd5caed09dbe249111edc61a4b4b47eb1c737b218ee4747e96f47a233b1e05385ca9ca476036e596f8b379ee0b37e8dd69e0979b7d9dd7281da57bba653f0d267cac64aef3f867ae187f07eb00636bedccd659c61e6b3b0eb95419b3984fdd1b771a2770dc14a9e8b2f7d28aecb403f7722284a4993f732234115458f7e9f7a9e1e07be1b5f3cb76272279f3fce1b52ac32ab9eaddc8f224e0916a1038979c8a4bcd1c861dc66322f58b5473424442412232d7ec4767af72085f4808d076fd9682e179f187c0d00f7f7d87728b522e953c1e97612ab5176e6c938c61e728a87550b145d798855e2ad3a046b600a32abe71837cb88f3927103b4cb5806bed945541210bc38de9b8e1ddb13e6c3eb77839ef6d6fe82c21acf5d0c7f96641e460137d04e39990b0ed19832276ce6c01e9568123ec3090c44fcb27ab1245418d07020569a062ad25c40e12f6a61af5071587443fc049099ba8d031b732bb77281ced782783c444666e2eb2f751e299cc4d136ac242f42ca606efaeb6acac60809ff726a3c1f67cf6ba08afd7d9c9464ec4c0e339540eeb2dc1d682b8ec3907261f8f4a39239fb05b332bea65c6ee9827b165b68258db688fa80848f0d1f239c86d0d4ebd1eca5179715ce47e79c5f4991e459a0fadeb916f67b4f4888a9ccc3be5f64fdb7eb1902af5fa6f156552c698f0dac12d0cfd1a8d10129125630db335982df0476bb2a6575aa5544913eeb81d67f90d6e89040621e7a9c082dd4df9aaf24c53d24f00bd182ba6d3ec1a5d5bd3397b7c4c201807492cd6bf511e4cd57282967b01f80067864d78dbce387bae29f3f33253c25b0ee0781fa732dd59a9ab54e312a3df3af9be6e73866101009a1d19f6e550507c5cbb1328793458d1568fe63220fbedb0bccf11ed3474ecc383abe7d8aaefc4f40d4aced03c24576921c6f5625d1454565f6e8d5f183288bd4f0504f7f109a110b4f1190c2e49aa44117de04c3821850e189cdbce99a27ad42d519412306938d309a1ff2d8bd7380ab424aa8fdc031177171f5b67a5d4144cc080aea4a58eede997b721ab2ef0a36737d39fd4aedff94c5ad02bd637580c51ae9a5f4fec9c664cc069d3136affbd0aba5aae7f507c5bcf14a26486a16b715060290426e1d98f7f20eb896897eb009a967c5de0192454f250ddc0c65e8f33de4585ec9e65e5b3b6682d34e0804724670db9ffd058c949e718928c9751e22971a465e4141ccb7429a9e8769758a77abe8ddff06284d4140e161e597d0234dbc8447d718e3fdb245d2da7275bb4459c13be76a3b50f9810fc05fd90950ae85ccd68ac690248e3bddd67916374266504e11772943ce4e8809012f3f5750d954e00c9350471be1d350df5839014ea8b7f7c274ee506cdb2354f84b4f54d27b05b06bc1f53b16f6e07b03d64742bb2a944b767b020bf4988c358acff67557f79fdcbf42361402fc3d3aec83dca7b00fcf38ec883f9f529acb29b94b7dceaf65715304f903db08688f2ebf085741c1e482faa18449c1c1d648cb6700d0a1fc7a439f65758b5606b9fee319de6a0950e576e7fcf10d2c2d2fb8c6c0d3922835e17075dd31f78305d7d348b04597ad93142f1ec53ae92b1159e316fb4cc6d969eca8b8d4be8da21ab0d5d55edb0421e3b2fc9089725ef6962c64b68ddd37749a144f1a6ae526ef094a777baa3d35264043c64abcfd8753e0319593fbf70287eccec6683f69ebbfb14a1eae825d610809d3c3674c3d83880aef088a09c398e659bd13eecbd9860f88c90e95dd265b3dc5b40c4aebb13f2a3eccc469b049142dfdc14b3b03ad698c1359e85126737cc0fc25b8fbf85ef8c0d64b5f2417f6bd572041ba802c60d8008d510fefa347f9b6bf0ff6133891f19951b9f53e53a0e5d590a781a8799450dcd3444eb5169784271b40ee5d62490fa46c7135ef7f174bbdd5afae73c589f0b281fe651b24e0de448a8d53ceb41bf427142b4e379199cb54ff90f5cad8f2770fbb98c1aaa2e4c09e2bb0e6e883f4cbb5406c3c0b38eb723fa6d588485c9820d984d016d16757e58d6f395c027368f6d1974e5b01716d4f0e9aab9155796749b87a67c5ec144a70790d4967a50888dd8bc693532d146326e53614a69479dc79df4ea1b532b3ba2e0498e16d310b1c9f68659ba31fbb1354e616e2d4a49b83422ad76f9ce1a5968b21634be85eb046c21d948d89fcf1b24833750e06e680ddb7ec5e3b00149d47c7e6f65be7f44a69ce9b738578378c6700fb355830599f2350994f4431f46831bde3cf49c237f20cd91aad84b7db3e939fa962b1cbb053409186b11aee941a00d6021d49c8de4455a1cd03d5e89019399f59766662b7544dde114e32270928c7e5eb5cdb42c7b79671e21176f49c7cabbc9f7d102f91c693e981d20742de1b49e14f5b2fe17aa7fb816fd5fa2224c0398dc587ac319c2edd2eff6f7845b412b008284b59e6140588de8e760e9027eb6aa13c9ff724059f09ac9fd955421d576745d7d00df56e02a233747d9151711f0ce7a39859ed15ea7d8e6d26380eea22771a0c7808f317e387256c49abfbe9c31f0db8dd170e5f1e0aeb838bafebe080f3ba768eec37f522dcd9a579aec663f9ff3b9635617cbf30940b0bd91ac41ab4bd27a2137370a4eeee1eb7290749b9e12672562bc5b43227b5a95c475a369071ec9a04cde9f102a0bd4fbad015942c2851a0952bd926d4db3b2f5a921e46ff2bdf183260e9a5965237f4ca9ce43bc9dcd4870cc8b6db96ac8cf933f909eab4a5c25ada5902212d5896f3fdb9e22cd48042d7c94a59956648409aef5dd80e4ee2a96be0758256ae5e0787cdf4597b2d9ea71901185cf85dedec60052131a5111d8b4eb4dfb8673e84837e3be891c3fdb97691cac6eb51d65524bd949fc58c8b0687c2a769837e7b1e15ed6d6723f69c3f9d838fe5c9cd22067a7c00b96b30ee091b80a38725a6d9a526ac0c50ef97a976d4e1c39fdff65dea95f495d5616fadd2825e78;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h865f290e73d038d0c6d628bf3a5ef72b2d70a7d0c52c01b5f29ff580e6b49da666d1a27658115d402ef7355e2b8a8a3277fa90d661d1e2357a2ad4e1de52c2d2e9095ab390933be8927b4c1e5ee311780c1bb4c0e6223746255a38e064945d5afe7d2e5e8c55fecddccefa449da2d8b0e58ec1fc1be230131f4bbe1dd249395a0bce495be2805404570b4866a203d4dd2edf6e07907e5554d3a1b693dbf777b1f0321e4d68dd71d27d6b8b20fefee30611b6526c923a45bfcca3043ba991272a35c84c5f37599842942d4184a5901774c9c9d4182ad549e284559639018d32c32512917deac7e989ad591da06b5a987ca8a54b4e3a50cf9909ed3461c05e05767106bb5a9de8537a245dc4f3f425202790e555fa8af25a0e3a9028378a77c88d7d528fd08abd41e0153fe9f5bbdbeac8fcca2576fd75156d6c9291a60b0be697e1b9eb308d32bff473a40c6867447d563849b409e024ede803f2a34b96f4d5d28faf22f3d95e82c5df70aa581f6fd4458f4aab1583a4970f2f36e3ed2f3fe470dfca42b481c552a914a7393d65272a3937989d38cfc1d77c5676d7466662655fae5d322189722ba68b9e1872245151cc4addbc351335f4b520c1ac6629dd98a3f7b75fab6e9b1c3a3c45a6fabc79fca5b298e11a801f81561b044cda0bc3ae717ced32303b18328b4adebfbfa43a28a9ee088a56a6e0de8f04df9ff85564979c40b3575d9b52e46420c17ad92d940c89f044414339bf193050e85bb4ab25138cf18b65de460f947491a23cdcb5db2f59246bfc44e505d75de94ffe044d996a52cad4cbd742583c14066b65c6688d64d3cf21990fd84739dcb591ff45058e71bf1c90848f57ed9a15b5d2756c2aff3a6f35efbaa0c267a449bd1a1911b4c2c3dfbf399b1e45c863f95e911f888ba5138a05bd0049638ff509b6778487fece35ef11368c1ec9a33e955c88c8043bf4f84e460da6cdae4f74e0b6eec7724916146f9fe653beacb7067df437d81c1b2198c1b49b8becfc795a3518b50a0a72c50d17aab3d2c95dcb095b93def8a7059656a137cda924fca0e784e6e6c2ff3310598926d233834fbbcf0ca92df0068eeae30f473704fdd13f941675ca8aadf22f97e74701db82500fabbaaa5f7c17aae1fdc1b228a766b6836849fce02bc95d4a41725a8ae945dc892a139514836b4a1be34ab6acef73e10074ba79921e15dc757f03c8517c56facf91e09ced322b009e0c6a845993f5e485c9eba7a3860a5071fc2c61888ffdd9c4a39ed7fd348330d563c91bba5a7619639edf9028f8625a040949a1fba24fcb8a931f50673ec38f48da08d0bc780a1fa88c8d5c3c738696ed87857fd3ad2a1463d3eacaedf70734c168033649c1fe5691853896b9391b1a7ce37294166115bc11e55e910bd2a93bc140506ced70ad2e60e7e82c82bb188d457d80f3e300ddb05caff2d6d4a6afd58fa9ec1c2412b7c7b831ca6fb8b6c25605a1f53caf902805991a92fe2c1a464e7b044c168d63f648f1669b63cd2c63f67803a1e2877e4ba3e5a2e79d27c026c78eaafdde30ee6af018d5433d0d7854d57a2ecaa0e39ad1ddf7e15fefc9045facb1cf89ce25d116c6e560781764f2a3bb518415f79986b6126c435c2578d68604c741c60ac0a9f3b073daa80016a650600d23dce03700fa77a02e3380c843c5eda01b4af69b2310a874901aacfc05d6956698c4682989df972695e2e521245219c71edba04fe29840024bd2a43b5bc1d07883b4aff9c1253d1a4b1892f2485f37d12e89e5dfff9860330501c4db40a4e5e708c6fe1d056d4674666e69c265e08eb407f235e2c0001ae00dccd7cae829b602692a7ac62ac618d6190799555b940bd479ed4ff7ed24ec77bd85f8042f567c42c4551f8593b914b486e8130caaae5c8387c8eea89cf0fcf5d656a58c3bdbc61429f81751c56596985bce28651845f21a273d4f31604d74f7979af5abf14c269b0060b2fce609e8e43da32ff775a2ab10ca5a341b84cae735351eecd01c8e00aff9dfbd22546f3445329359b6103d45994126ea097746bf0d1f64b93497f9768d5107b1ebd2865900ac644a2c1b67842f1915331bbab3acec286f998c96fed5d9b3619567d431701d3025240d2f966e2de33637134e221b75f9361876fe1d11207dcc01d73ff89dfe1300f934066efbdf80afe7c55f834d550ae82f0a93d92f118ec631d8b0c680d06a170983b80bfb2a6403cd72a117e164e59ef487b624f6c3217d5ae9a8ac82ff7a6d962849e83f57868a0c132fb4f28abd8f766339523f82bfeb7dc049b24c695aff34d3a32a95d4b7042dc7c2e4be2dc6dd270fe487d04ec2df9b18a006d18fc707262656ac2fcd93f5b9be27fe6a42a201d019fd47259ce7128d1c1f33fd26a04205abd970cda1e7d34bae46a6f0f94a15904241ef2cf1798835df844ca78f94b849732defafe85f1b0a2e59b0e69b708ea5ca83bf1b5313e321792a55b28fd9254476d9950eb4b06b8cd642cb177efa0aaea8cb35c2125b58a8592a2bcda92564246b3144936e94c7945abb2720e640702a4f4bb5cfc39680de6412bc955eef8db4e4fb2f97f16fe0b6faf277bc6a36184d77c06a937333c8ac090d164f7ed7632f72f04a26f3f35c0e3cd20557fe32de2bc0a38292e4583a2e8ee38974b7a43ca03f033dd1879408c0b39a0cae7bae8f8b41195ad7160a98d029ed2a583306a41121ad69e3fbfb938f24c8db693734884c31f2a9ba9340e02c2c00ab2dd7f42ba4f59b782e1d26d88f4dcb7a2365c5302533b6dbc1ea35bba2accb56ad851e272200028da48bbfcc6b7a6551c33896a3809b16d69c72cc0fd3ba2449d40a3bc4957fcfd082bb643604de61bbc144ff5e02362e440dad8c7e23c8256f11214dcd048c11e9a1cc96eaa1279bbffe0690a4aea581653761b4b012b137a68dbff71ed01418c2c4db1e3a710c032e47cbab3cf48425078b4e0725796f7a6fedd669023971a0576ea9419059b3c91a63db15048fbb5ebdb2e8fedaae95caf07a2c6c6df6754dd386ce6084a7bfcbd19d31aadee2f27ad32bc00cd2ad83297a1a041f821a6ee99c9de6e1ae8d01d5939d7993d36e786cce1ee9fad3e4738827d26a96734687958009ea254297b77cc70f913ca621757893b64206c02a82136a7526d49654fa1b6ab6567eee76abf01b0e4886c25deaf67e45681e0fff44dde2c6fce59706841d15e39cbf61e10461a2fbb65b1441c93f960f90adbbcc5b46840d67d338c72e5205a0a26efa72c9aabb57a04b4af57d5895382c0b846d10ab71cac5b8fb63e47ab049a1f0b05b5dfd9d6d73b9ddacb4dcd8776c1a18b295f111ae25bb8302d3c36083138a64509b337ae67f1f1a2457789bfff9574a73b6573bd3439ab8fcdb46fd3ba9bfd76589e5613b88ab8e074f5e13dba91d621b96439e376df0ac45aefa1f1f804ce3e753bcbe710f1548d2662cc17527fdc994e26a6318d1b9bdfeb97f1e567b30e84c4917af5f9b643f7c3e99f0a5b0062704e8484210f70e27123ffcb5d26e71815911285b3a0405b44a335eaf7a7e82af762991da3fdbe4fe89d53346e258743b99daac48c3ad73ca7f0084b57286d52595024113374e86794464d47258e77a7c27364671e7bb26b7be1fda2ed91b0a9770ec59358219829ba4b335ff51fd12e31e1cd81b6ee7267f593df9ebe655345ac6d1ba1254d54d2648e6415a09f561f5fe6cc89993ff1ce142e5bba8c46449be98e48d59492ee9e27ddb662446e2fbc4cdd027430c9293ac238d7d20bda84b1ffc23b67e2ac6b836f90f4c5e47ea739443f42a9218ddadb93e009c1bcc99318c582656c69a6938e78cbf7b9cce0c655dce997d8e0e19da2fe0f1d4cfa8fb0de6f92020dd90cb6100368980d56d7bf4f4324a4d1880cf21319f5a348a5a30b6d3e853dbf5cb0ea638244aecaf77e10bcbbafe5f66ed73041d2b0c504e38ed6952accb5747a6790faa934123d27df6351f2d272c2ef7def8367815af9cbc5c8add2819746ef55b35c5b955624d66807043568c6429e7a436dd5b759d02d4700e2e9b6bf91b890d4f11c786a4a49b31fe247481c7d621d9daa4588b75bcabcb263c735a3202b29cbeae18c3fd3d5b2fdd56b954c694e44c653542bd33ce89576d094045939deb9758775729144d759df7e5625b5845e69ea24177e539c26adac7572dfd3f75fc0f38cf86e7bbbba5a2285f98cc5cb025e7ead30b1d61f3f7fd19a05b399b253425a86e075d7068a9d181b9a0428861f676d504326580a0a69fa14c9b8f05853faccccd01c60f54fc04d5675d7bb58db22823edf21605353e1c96ed54f230c15226d2180f6c1512f994b7442652b64cf0582082b0de49a5ddafb0544112e347fba9020c02e4220aa1556feb419d9f5c6f63549b4ff576e4c3d0ad65f1c26c82b1af7d5a608451c279fa55253ab0f618a84436703829dde589671decf542d12ffdef382b40673a66c88805378f5a638e327a94bbbc10b3157c1bfd3627ff892ca202d8f847c0446527a665ea329e027544ae582ede15f074dd19907d3e1118fc4bd07af81813f3859f6f7b7ff3cf8b38c2900261a2873762d59fc084989d7f4063a205505a41966b38f739366738eb87fbd8ff5e587a827301d84405d0631371b84527548535c641008faa936fbf50ca56468f570e27a0bcc53046d2a314aed1e5de86680222378a6f75df0307b1ce9ca08db0cdd015a7a8dc582f0d411cc78f3ad79abe370b066652fe7e53acecda47203993d6f93bf492e0cd1726d232f930a9116a3d524e93a65d9f0cb75c69ce5edf5dcb21928f6d1fa4d900ed4e73bc66af91f7472f355404dc1e3065a102e234e482abd8a86231c9354ea7ae994133b3bbdbf2cc5b874fe27502748d02ab20d502ce88e87aeabb96cacb0340709dc5410f9e1e13fa9d9d61c56cd3cdedb6014c02a4b29a4cbd0ccf1efed2bdf9529cba41da535a02b1b3eb370000343d3898c7306bb9ed2d74b6be17ae5a40c1a26c4035b3fda5b071bd17ebbe6d466a460d36dfc2e6dd3b6137afb8aeedb1047c982e922ca40e6ef6c9f39ec3504930671d5c69feb85c7e5205301eb279dcc29e94e8ab9e0ab056a48a62e23a699ad16294e09cd642d8af45d4c783d501741d735ebfaa10b2ff91cc2816a96bc69e0e3851e1aa958dfe739d49c4dee500dd6cd993c851cb1f8120387887e87d6f8cfe565361dd8937cca69bff18083899c3d6c2320a77a8d4bb2af7db5cb7807736e72a2cd7d955fc1421b8043419a4da231a884971dec067410024d02d11a3ccf24ce6be96bca98c9aaa0b2ff21a1f477cb90c6f910e4c6fba94e16bb40f019170832efc463666c17c45c59b6713218ac49f9ab3d6880aa485b1f78ac26c04da001f0a08756efe41bc29e5315b9bc66825ed0a97aaf2d3b0dd7b09760992c89cbf08892f81aee53699234f2b52a74c143cca9276b2b642e3da9dfbf752df5956eb295a262f220ef30d6246c40004a97963a8a95a8d77a54681bb8f744bf2b9e7a9cc9acb782fa8c31959fc7b97d5897d1d24de0bb4e68842925f480aabd2bf4033747037a8e2fbb2d142a97ecb555f86fc2ed82a55374eba8026076933a5a6b679fb114ed32c1a476d8e7d0427b3fb1e47fd0e5d1298203b68926d93615eadcee574009b331eb0fe42775dc8b6c22330878aabd18009ed2b38d0f01b2f44248d7f67285606adc0f654ca470bf5bb55df59df2830f6e9331b2837c8e48de55620c7de2446e4036f9964460fabec02d49dbe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hdc5e762e36de08af841c4dbcfcbb7541c4bef89d120768ae7c9d5bea2c48f1ee01c8731f5b0d16f6b12f44754f2301b8214178801a3302c434d5414ad8cb2f6dede648178340a8d44db865681ee7b8cfbce1a30cd8e669bba1c774cb80f96bc79e03c718564f129802678fb91a0626eddb1ec35cb9dd62c407793b57b0a17070bb271dadab94adb51e9d27ce716f0147f06574350064642270a72fcc9f55b2f8621b86e7c7a12e55db2f03186db440fd50c6c99f8c598cd43feb7c562f6f608c1a49ab3f3f06034d046a540cdd5af9871538246fa4a5835025687d435674e97e9a7032ebc649d8c3a0bdfd935cbf7e0ad2250c08146a6cd1498ecb595507c02be1140fdaa778e139b029cf91de3647d384b4c843f061d097bd232ae01d85e96704aff86385d666b4b8f5f8d5a5ac2c7a5d9f8fcd33c237a5209f80e78c840ccb64511c2b211c1b0de2b86dac7e10704f52057dd1a84fa6fa2709818c90e9c919ecf536a7ec8ce6980f1f5361a869845ed7e3cfa2764e76e129ada4e75572bb173b4212a5fb0fb30b86c4f9d72eec5078390154b95dab36b682bf40dd29c42f10e02040ec66ffa56eff08197d37a22b44f906bf4ce1eaa57f6adad3a437e18586e408ca54f8450b948411dc865201698e1c4977569671e600b6362466036baf35416fb615a869825952c7765e7c1f78c3797cbe729548dcdfcb0ac56bffb1632da7a7a9dc37f5561922cc3688a1dd6f24917f9625e4efd1587e7f39ef7b81f59c1a0b472ba1a8a5dbd13ef30b0d85e1368b54e1e732244bc4f424f151fe5d16a4f1ef36d59c2e9dab0230e137b1160c647806f02df9cea79af9d31ec2238478bec71a1045806e686775930649c0d39cbbfbf1080ee79f7f48f452549f21b4d022d762c95b406adf783327666a2df4b023727804be1e64aaa0635b1c153a572c92296c5b2104d5a85333db3e41d3571193cdc65f01c5a3c50ad66ed8ba5cc75ea3562a561703d0680b4cbbf200fac6f76f10d1fbce4f4002e35ca9848065219d76e32f09d9a5b0ea46f2cbd141bdc78467f7d1f511223dd10821b5f8ad673eb647634ebb08bd998aa6b837682d50a42e78d9ee3677a2fb17411d57dd4c35c3e9ebd57ec183dd877bd6d4ae97ab102e725136f51dc67dbfecde8390a4897968f1e88b8ca37f85c42dfc28b26f83c040ae1b60abba5a05d5ab61d210f96c67568710a21dc44bddb037fca60181c05dfd373d0b8edcdd75fde0a79bdb3735713910f93cc1deee4331016501ab7390d954e012f47b42b3622dfb3907d7b59fc72dae80abcf5c9974bb533c63bbe74d06eefdaba99c5b96a538dd5bf3e3efe325e377d5cf8ebe6a54745ecbd18732cd15b6d6f0d8083a87e4975fe60d2d0ea5e5c546ff41ca01071e1503a2379250813716937f9afa46a860a335915fe37fbeaaa1fb91862146bdd9c2da5fdd5ed4bc35934502e91f18af8a1f9a1f90678ca122f27c9eea17df307f2a704f6fefa9e20eeca93941b60818267e353f1dd8adb95c98f9441528011b2c66dd6811212cb8e5af1207affaf441ff72f74fb87a5c266efdc082d1448938c72e2e394d430e412ebeb6c73c43d92690dbf6e34c1359465f1fc966444e65749f097c229530ddf32e4312fa13ba9a793e803a6dfe087a86630642705fc388980b65af1b7e04457a000bd9d2a46f159c61c0a2886bcdb60a46fa9357825c15d5d0267a57dec0c54cb1a09a37622bf32b0a7c9ff90177684db7346d4cb15d8ce3e1440997012dad095010bfafebdeab7009c9e36767ca6ce52c3b62dac942d34fc37524fdef78a76efc0b55f8d8602c0aaa4f82284667cf1135852639409a9a23dcd91f4bb535fa6d43b84c0f5a2d263a65f4d17820b7cc49eaf3c1c990cf288d417d0e08cc1984cd5ebce62c454716b0213691a601b8ea279cbe8c186b6005b17062e993a84a2c7a0f3baabb4946a92fbad6cda4333139ee1222ba94a439bba7406f9515706d00068bc5c470f744ae789372031550c3c8f7f378f194174d1964fb25ff906e3d11453bad9ad748dd25436ff02938d41225cfbbe03c506893341c9ffbbb8bfb8eb93ba93656564a03d657d5731b2c482cfee689861dadeab86cad98540501fad7f31e823ada8398516459421bdce29f76e8e854994dfb17afe1ccd8ee53b865ccff4354a96f2b8ad6554411538caf0a8ad20c05e6eeba0c214c8e5c75e27d8dc4b4f04b4f2725116c5119d75f31d1c576271a91aaffba5028d03fdc3ab739c3692f91ddf5ef2a7b3004b939ede9135bcc84e64e72bdc0c47078d4c6a7c18e23459ee016eefdd4ac6d6aa5e0a53e06e691459aaf56204991619e71468fafc4fc5c4a1c59ac3370751dfc02880e8fdcd172dfd472179bee77fdcd8703501dc6636caaa088859463f4e571d3da7324ce9f1f580e612a26b7ddd2539e5761ae08b16dc30bfb6457daea533a25444a0359b59612053b6867d91fbafb107f5c094a73b77501eaf81b12681a6be6ded21a78797732eef7f7d55ed911b75b1442be0e3e2ecb3b2cc69cb21c3d0e37b18b05a87b3c4e4aabf4a4741ca4f50d5633af2152a56b5acccbab224b72871172a13d3c37eb3194f842c6b0f3e5cc04a15d4d53376ba51fbbf2a956e14d9a897a2750e5a166c6c2c2e2cb7d471915a605bb347bcb2afb575b7d264a8eaf9ece3d0569a3edfaef5ced10a8ab478560ee77b1f7f21d8137f32bb0a4a667b9354a9621880fcbadfd93754e63137ca0979fe461d9e0a541b1aae4961b4c267dad1abb8c9004a063b1449707007dd52c2f8afc0eccd62555771c8b46075984362eb63b4625adbebb77b6e5c7dbfc4e481ab4ad45f9b5c9748cde98722b5a4a9c90f34b69a77ec89c829bbe220e019c3fe72e008be5f2843e49c111fe5415d2caa095b5ad7ede9d39ca681aa3c173f98cd851345e97a126a3d51cd329afed37f8fb2e3def69eb70343a7b293831eb4025e2d355f27680d916fca1c879f85b0bf37cc8d6e79defc1839196047b81d7c7c249160b1334562876ed007451023638c111ffd152da523f5c9a57d829fb197f3a04f67091d03d9c1b0bb36db7acb24d4af37bf0ec3bbee2e4c2ac583a6d289394fa1d9f7b6b086f9e64f5d0badd91cf9e389fad4ecacdf2894c7e4bc3393d96a852eeecadd2a128bdd6819a0c564d413f681d32ac1d24ae2d6dd16ea9e287257dd7d2b4385bf5c6ae340a13123c6c9624dca0e21d0fff93300787195e70eae413cfbb0cbd70c7139a3e4e3e2b54a213edf507c1ae84dcba712d2492b27d8a7cc48b606626650f96e91c83f0160436d580bcf3d3c96a554bcd23af14351a692e3e2bbf0b8ee69e23cb2a6c98c250930c11e57cd742c163c7d51e64f49f98caf1a0508710e7dc144cdc8a523bec6fe15c15780c60cbb3d208261ec737c3b14fa897007ee467d0a81136fd7029b961686cb8e602ce315f93fcc5df87676500152d026008fe60b5d21cfcec6609b28abf9dd1037a53f5d74f3f39c14cb35f782b3eaacbc00b0cf6c2a46d54119ceef348a540dc5b933509607f7cce61e6d5de4f3ce54fa25aa5857e92a82eeee77bbf37204c3903688a3cf1230e44a473e44d0c3ce264a8cd793046ff4ea1f0e77764a9198ee80cc37898e4378eb8db424cced75e92401f6bc2255083c49a248fffab291e3db190c7c65daec1597c302c1aff02ce2fc07a1fd5471712d2acef9d04555d9cf9aea38e1efb476150663c6f0811044376d7cc34d78f411d805dcd6637d50636114923a2445938dba9f136790952c0d42b20ed62424108745e6e576cf7f705d071692fed85e4a452ea46ccaac4809c01b29da20e44e44366eabc74b051c0d5f8b7ce66eb11e570a19a22cc971a09adf12783ba2f15f5e8fde16c5e7c2c40a6c451d6c9e7a303bd5e4c647ae564e0e85540a1dc99e98dc8d1af8f3accefa7ae004dec2e0b3915739568ee659ac320f11e36fec953d9e4bff8546a22ed755a6d5c6bf5325de7ec69c758501496d8bb46201bcbec30a83f5fc37236e884ef8c27b495d0ff017abe15e50d44279e8fa22fb8c5db85e20de32a93dde5e00da8c1a9952848ebdd422c4e42e456a987738bc5dd162c17fc8358d5e1b0566ebc21c06a5ec50fc7003c0c96e954743ff94f096be0d35fef2df62a2ed5a5d866d37d71b86db7d387363af65d58b146a3ff85f9051fd2980f189a9cc9434e579e26cfe7c24d82e528aa9f8ffa7b0324ea9a4738eacc18098f92c98645909ae09c5dcdba0097211c60601d7f55640b68efd56eece3e3fc6fe783f94b7fc6434c2994671c2d566955e2027209478d5d1581a0e19741d6bc3a412aeabdbeb67d7c8693416710e7502f92a51c8c824d24fbb2f7e863f5f119fa3797d9426479c30017913a5391804ded82f9302edd5f4a902c6f66f7ce0e2c023f4a22edaaa66b6de8522cfb5e28d29759c9bff229b5e6a7660f99216c16e0be6275ec419855a2f26ac64a9d405953c6681579ae6181c4d4c347068f46aa492695cfaa7de75d9aebf0cfa35136a3bee298b0f0e2265346bb4e0c0f687874ab888346067d2a0202e5425424096981c64dac43f2ae332117be439781e8e137cc85f9643ad6629786bc40bf92a1b8294cb54ef822580df0ad12f8d94f4a7c38afb403e36ee8edb0074fb56d7fa74036f69b18b60a6b79d458d6534cd8ba9ade2617f1ab94252d0403a8d6d95553b3e8631e5e28494df8782b59d9b238b5dcfbc3cf031a18e60c6d37103d6b1a6e7d423eaa8092384ba656bd06a14dc646cba42f6a3af410b964ad87e464222fca420f10b269aab91733c36d492a6f63bdade91dd6f97ff31013e6a2a047616ddb786a4598d35a2082a5b7fe8abd239ddcb2cd5fe9ce1b5057d55ed66f38afb185ed48bef4e800356969a1ceb4c7fa4e9d539e571790ad8c5f6dd5c43841f79ec087bdfd4700f2b9609faf7f428b35bd6410f4ced4b73d51989fd92722f46daa0a3a91c0efaf60fbab2ce04f3922fcfc0b9499bfb0ee4cccf0cf2387d64e10ca362184108cc67245d7b68f45a88792303e3ea71833c019d289ed0aeff7c186eb0acdeaa588c3671380fdad385a326d74b391c673a85100a560c2aab78297be29fbf46fd8ce1e5ee0b98f6e5eff5ac198f17c9da698f4e94566c476cdbd2b8789b8691197d89bc55c5fa14ccf9eb872e9bc374128b4ef53dbe433b849735e164f4a45c39882a215eb1a70dff34df5cc4a2d0f2123610e60e7647e5129718ae22be549dffe1fecef6967cdf40a89a8d97fdb73fab2eb3f8f4986498f32f41b16ea2c92384b534812d97c2ba233205d16090b11492010c8cf1ed73f23a621248a23b372a10007478d275d742e7ce98a616e652f6999befe489cc55b0d9ae21c3b90401c9cbafbbf7fe9cdb481c157d522b2804cead7142d5a0f1a0b726c493a2ff53ee40090ece81e578cf17357d3f9da103806afda90b22b9e78c7befe6251ada7f3ef43909139124243044175a9b492a5b62a7c22046da5f9d22aa52639a9c273ae03a151d7e5aaccc8229b953d828d7589469fa31f6f27d72bbd40b53aedbda06fc95fdcc29e42f82840283458e0546cbf2df1cf227a86814fe4ad7f655872e187dfe168a664cab29b2c201d6c557cb78b8d4dbd7146f9c239e6b98fa0e580032f6538041a6c3d56c25dcec8f36116e9baf8f3d445391fd2db38e1ac5d97169e605cf011c8e33dd45a3cd12ea7fe60042439b6a086e64cf4085b726af9618c789ae374b7f5749dd7a1f90df59448a6692805;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7ab14355957cd14174e35b43c48c598ffa0ac32620fa246c46c4c426157dad3a20ccd5c1561552d26d1c1fbcbb8df3bf85ac168c2cfec4709008fe3079f2409920ab99326930d2619922da48d4331ac0e64f127f2958e7bb9764dee697fbb0b27922ad107000f81cb8849627d45f8533f1b7635b2d1ef4a3f70090f0a86bd1de0b419185dae03d5077bdce184fbdf6edb1d77558be154835af19052d7c71fe0c4aebc8e86122bbd31ae268f7dd524ec9831a56ae468af87777112db201878dbc010fffe5ad30497a0479e6e40c764db8e3b5c3958e963146f0ddf9bbf67f7dc8a9013ab79ab3c022f75a550939b0992f8b314097cbf176ff881d2f8e556ef5d1d2fcc0e1d2824681317edf23f282d23b16bebebde4370e0376a5d631e05da40945c67d41a8e73edcaa5277845a6e4fe5ca1bf12116198866164081b2f1973f41861ad17b53bddf429a2a2b151afa6ef7c7e36d9170a6fdd4d3c2741b8e333ffefc9114b50007ed556a1194839f1530487e6cbd55ea8061fa30b69c711cac91974ba6d2ccaffc96c4811c6d3d514c54521ef8a940d94a1c16d9125ba33be98637d2bad502f478fa1e0635f13998ab4f907ed2eb0ed247197326a3c36bcdc21cfa1909d1736f942d5db7aaff5251c03d6c861233355396394fcd136ceaed2e93ce22b016071ad5c02c9866a2cd84fdd390a416703f0aaacd5ad76a6e81f83903b517f13ed1e70e00d75fc0567acb31c81ae40c669e1f0e1d7919d5d2c9294e367f289d00245faf204d7e6355f72db631e52daf914613b56bbe3644fa31d4c85a659c7c7ac358f810fdf15c7f15874afe12ecff2efae145f370966c61d0af8b8391dc439849921428019e0a992fde7d5d40a5c0ca3d2b10aaaadc927b867b7ace6deb403de0d92674a810c8d6017dce08943f92c1276bb039b1eb5332ca1db5e9d229943b641210c052b4fd34d05381f483d156198f167e2d02e22e2a214d9ab0265c5e9e26134d37820469f60ad80d5c8a401353c6b9e039a92726c35d98d10e760d53fb0ad2e0cf1a9171d09efe4359db3cf47d17e845e6c9dc0ef2e855abe00c94fd0b94baa1267e44fec8545b7c679a6264cbaf25b05352187fb81093e8b7322271b521d79c3636dac01542031f70b3ae70489b1efd03203e95bda5f2b179bd487cde1b3625108e614d63f085fd528474d98d009e5dcff59d28e602e191fe0dee0f37cc65585f60105a5f017bab0d7fc483e582fbf6c4cb1efe1de01f15d8dc482aea0a8cbd91b84f0af91a07256b673bf6664f554afcb02290056f0e58e4de6a308f64bd90a8ea1831992dff11d0468f229121f801944fb47ca55fab52693ce58287b8ba3597724775f9dec75516bffbf75062d3091a9ae130ec1f76fecb0569044cb2015b8577f399fa3d572c91e5eb87345350cde08c86c2446382e703d825392b2452d11a40e75c74ef32e8b67cddfdd0d36044a36b9241fd6eda7e5c4e2d963d362ef43ff821e51a57ec9eb43e8ce18c7efa376a01381f40529cb631bd9af5cfa0bec7a789babbbc1f7366c9b16d93d8a861d4b9b7fe5e44a1b7d47878480a59ed47539f5a756a6ccab52cb5a156e161cfb36e86d6cd94ec5be9cd1f8b6f2b961b166ef09cfc76f967d9311fe01b2f7b797e1d022420cc2b43aabcb4aca77bae702fa0da2e6b9fa2d0dc1cf8ed437b0cbbc9bd59b3191a599a79a6a4a4b470c821f1832babc09c23950340af8a7eff63bb19ee23a1508169eb8b9fc291375d764b10ce7e77bf28883c68c195b1aec1099d53b77516050d6b6db825dc9777c7880d3b1914c2138f85f489e87ba62240744224dff90f956af27276beae0c40ad5b2d5e8b2cf0d27df57a25bf1c63bd72bc77f8ae0d929f5d0234dd60720db7986e3f917f49d41cea9c4cf8201e84ef15ebfe703901019109e8ac4580a03a565b8afadf1ad53ee3045eee9e919462f5d287183c3ae438dd9fc7b175625b67693cf4c4b40162c2a6101ecd8305943aff820159940bb8a36a13ccac6b8dfaf764942d86360ef784ac519e9edb0dd3531ff981f4b7e782cc22f723155fdb32d3bc96f23891e94031ed3f84c9d7ca232cc88a094ab9543106e9c99bc151655dcbf6dfe8253a4641af506d4c9dac346a28663d065e4b572571c74acf6f837a5147dab9089feec67d8a4b93e1fe5f2c61914da10e134acf2b2e508c95ea9ffbe278d78c9698ea5b5d3fdb3c29a3f0aa7756e15acc54862c932b83bbc641fecbcb8e59c846a0ee0c2285420852e71fb0ae270cf56e38ff78c8933475b1aaa701bb14d59cd29b779447c114baafacb74ad0a103e98d9553f233373f13c4fe5cbbba0aa7ba940c2d3e8e933cdbfbb51e9e1b0044b99cc902fd13490dfa3b2d3bfcdf4af26ff6c5899b3d501678d24b8af5e473fb44a3d94badf03c9af3e60adf547fe9dbc9d786f23039242fb550e05d6ed80cff0a66ebac35f65f956a9d5ddd5ed6ee3c94c3c1c57a48859469665eae997c186816a0ed8e9764dbeb8dd8bc31b1ba1fa50b54255ff092e54736806cf50f8e78d9105d80dda6c2df7825ee7df3200f401b47e30947c191e021b5c4464837b723ce3ee3167f1b491636abcb48039d77949b511176e817d462916006f27182916eab1eec4c6551839b1c27313c171a026eefe9399194fcb8a12a7ad6221aa29c28ca183071c72f96a29b4337225c15d26ecfa41cf91ba740de43608eaf3f649f0ed1b7312fa503434f4da8b007681897074633a4cc8d19f8c26d32855f3a2a29cffa2698b987b507bed2d62b797f0796f1261312191fbddb8d74a07eacb246a7ee4f4925d7063e01652cab2866cd51623b565ba98d97ae2110f2fa84042b2f37a9bb63263f080769087b99ff6bf1b2ccde7fba1bb156717e7b0501ac4330a1bb16acd9c43d42d979af5d0e7dbb14f6fe2b797cbf27469bfa2619146ee84b437bb24e193427ab32abeb2d32c733f600e57be34c25027b29fc53cee81b88868c65aed76205def99563c4d0dff913a1d88ed451309ab8bac09059131ab63faf1191efee192b05ff76d4564475921f7619f86225c197358b94ffa44a093ede0fa3f1c84ca38a06a0a80ad802212874218704a533d1d7ee60ee3ecce233660f8a48c1c2dbe23fb0e802049fee915f03261ca740e8f65e2a8ebca3224bbd8c938cd64f5154c9a3f092f7c1968eb357055f51e1cf4bd16be0e30db4021846251aee20a307b9f9dfd8d6e3c2af6e071042c27d48cf5baf328b3d8f01f73e04120333211b47b4a26ff0790d0f420927ffedc395db9c67db1420c0a0a864990cd618cd5905ce38c1c735a1001f3d072f03202bf5ec657ea188baaf87732e9b209b5612da4cb596956a847e0f31cef0cf64e1392f1c88226948118a897daaf9723accfdc205452b2dbd2785f519925a14b5e97348b319dfd3fdb603a43e10b72a377a2896643abb79934005f90a031afdcf2408be6e10b592257664fc1a7c35c9c5d8293c39c4953ef05a9c83c8f8a64de4108639ff3323aafa20c40c14a30b8e2bacbca8f2f2c85c9870a8d374948e0b6e98aaca3e526ca229c663e89681061dd0ac8806419e2fad98d6d131d94401398f82f88b20c663e9e79eadacb449f45eb23ab5a2e656b3d740489eb3a28353b1c3d1c39d4f995f616805fd0a9fb133add4053106276e6aa24826a274cc87c1e0c6937fb05f4b2fb8f0758af999366377fa368c3ebc76bdd4ef325b63ea162ef0b4d39870470b74e93e93dbef636e3fe2a8e9d1836e83dd159d478a8318bde4706f45a01bd408c99ee80144a5c64af75126e185906e9d3774b7c5c40ea58690d804b8fbc7b74aa08e17434fdc27c12a84635b4ad9dd6226f7481968d9612a38a3d0dbe78d7086bbdc22d1b0ea89972747f986b2e0f79a580eb4d100046e3cd79bb726d08ba99637389c4f9851e09fc3fe9f3a75b3e62ac189db4a76bc30ef1a04b52c35c5f22cea8a1fe3e7cfcbebcef09a39e1a4b8447877cbdf3de651a63db09bf68a72192ebde22b991b7521a4a37193891dd2f7557ad9217b9c136bb4249c0df03e1145f7b7b5c7be5db12f695c22f3498044c32abdfcaffb3e41f0e97b64a48999c80ca0498e1135be5c431fc564706afe9b377821046f37e1665ddafadecc5cf30c89aa83428dc52be1a696c9a50b0c849b0d7175f9ba73ba2506a47b0f2916354cdd9a6d1df0be019e3d22dabfa8cf707ca394a89293d277b94e4ed040d3f4c8189c38bf9009be411d03110f7ea023a2ab5eb8b32b8a6a791c7831e88ae8fce860952d54c1de68be63bfad8f8221a0fe262a0be62917165b955a3346c882031e99f0b13f1e5f1044d4389689174e310eb268833a456365b4c4cadb636d8831e9d79e8d9bd2d15e49d0ea75268e20743fd2994f1f6e8376e6d35614606e76497701f686731439f1547168c1c39f36bb2f42dc5ad73b17038f41acadb5e19d5fc8375ce49ee4969089badce3c07cf587a7ce1b2ce4256184deffeb757d321f1548a2a95d8383afda35bed4d5c11cc5287737ad6004e22b71f192ce17f3c7f971950de58b934de3db5ecb38216e15b0677085a8bcb367b73f0305503d50707657075d0edc9e52ffe5a1cba4480c1e83aa32b20aaa90ef64fbc765ca2ac30f42ea08ea07dce7ce3e52c50b1289e6eb9a3e0bf6ef0a87c381266694bde628002e38e3418ee494a3e467b0a273d9c0235f7145579a580d43ab4f05a0005da929891013fcc29cc95072fb6442c8435f233e5ce0c4ac93582fc928330b70cfddb9718c1ac42bc7f3c95dd5bce51877a31fc773a845c5761eb746caee797b2895dff3a2bacbeeac12da3998e8d5d8d7b7e37caafd824dc6f8796cc470707352f5e1deef59c5c04f3585e01b32342115c72ac8f5199f049b1c66ecfe6104c2db3a0a188ea48b42c45e81ca0caca939dc65c7eac9e9b9f4dc22eaf776ff5dfb0c31ce07cd09f03d94cd39f531c058cd78e1f943bacad1ad7cec037ee617ae7b9eb3bf07ea983a16a37165c93236489ce944e60280c00d6dfc50cc1b119687b2cfc6efa880d1f3f1abb1028aa8a732b569a0efe473d0a0517d56611439c7ffe476414c1a2e79a2fa7210e9e1e8c1e17f59657f6b03e594127d989f280288d4711572a015cca2aa36f5c6d56ebeb7b990a9a7d99c4d74f7b07532792ea92fef6a1b3c2b48d7bcfe5935319503ab103a66afc42b44b2880a52ac84bd27a79b24fed151b42901698968836ccd7e3bb46341ac83109e38461d064a3a741153fe26f85f87d48feb171bb529d7fbc0e2e8645be370fe0639b179ea4dbf300922e7c9bcad3d1f70c396f03285cecc7cf44bef34b00415a0d79bbcd442079916b15e00cc2da07fd25f3d4e6e6d12ec7a8fec72dcfbab4581156ee48861f3ba39b2035e4399f6c04170563473f7d9b149fe47c2344a3e456549ccec5ffa348d3d87a171609067fa8fcef220504e5d886bdede744efe333a9e56e0e4e7d34d3ddfe3f51783c18650af6faf1bd94f2f0c0b7633420840db2d1c66072b6acb3ec4bfcd7a8581fb353b85c33754b2a3a11b2f51b86158f651584232053a526a4b3ec10061521d1bbdce46164b9322d8279635313faf677de512addde153231167727eeddb2bf03d78dfe5201cddfb79d65275a26b8c33b004bd0cbdbec555857a2f07c62f7aa84506eb1d7a784094cd98389357e977291214a05838b75e8fde48447a8ea358c450f29b6d6c8fd6910681e7fd80521f456e21557e2ac0df3d5aceb5ba6a6156765898ba0c5a6f8b0b77;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h142da285bad2fd34ce936ec2600a1c9958e3bb98dd535adcb468d7ea46224ce18dde04f606f36f8ce5f752674ec12f458e906e9189e7c3464ab69c8000c1fb3854cb2068a5ca3a89db58b1377a4b40159b62c33580bbcdede8862d2ad37e80fdf1ab948aa031e3ea2e2cac3dec694c01a1b0037a1295b706968a042fe112e5cd7b7e59860f38c722e9c3f83677884bdbf7176c20f04308b06984d25579a6ac21ca990bb4356a6a513b54dfd959d6eec7e9c724633db0e0035c5a3b140c081272caad935dd61abc55c6d5a893cc54886947919282a5d073c468e0b78bcef108744ff39348a15cf4f75199164cb46130f6a3ef0397bfd04aa3fdd01a7354bb03fe85964df4e3534a723de2571d17b897cab5731ac618bf9ea66e599a377e50b95a6a5d48650e9f94e3a0a5d41815c2e879d0a1a6ff9448445dd707ad2358c2876fadb5a23d8319fc94f0ca5a4a78a6b1cbe951e9fcfd07da978d513cd4d3b20b79b6230968864d834709c64f424fea368b56608d6554e2ccb0f2d1c3b438a804ba4517da002c1e81b3b473a08f54377dc132032098ca95c535db3ae26fa97536d07952fedb2f8625cd45f6af00df29b4d3f81720e020956f1ea86703a5402a5e2aa8edb6609248d9e607272ce589d3dbbd15da81b5ac72a66530cf94fd91243c93e1d9a5de003e6c559d9891d3a6bbe8e171fbdec5013822282c54a1bee698881b0225faefad9fb0d3d08bdacbba80b7549dd28bddb7227789bdb6924c63b6953eb1a04583eac3ad951901c21f9f0943985457337d8d183560826fb8668a0eea7fea8d8ec40096d578a478227ff8dfc8663890f42ced072c222566740ed1abd3a82969196b43a2a6141e18bcc7ee2ee4ef91fabbb8032f3ad1205c4d68ad08fef4cf777165ea63dbd99fab432bab6afbf2ca2c284410b450774c4736976662128110b2399a7297dab6326cbbabff3412f6d9928aca65be93b5c8c9132cc1ce5497ae5b756e927d26bf235040e400ba7acf98041528fcea108b4e396ff9b0f76b36b5cad0839d39f663fd1818abf8beeb70ffa943164fb7526a607e0e7e5beb605f115ac0b76c996db423cf7ea6594681f2f6a84b353c433c3d8a8c6900e3b14c8942e6b2fc6aa028d1e28abbfb506012809074270cfc55fd09c6c51011398d6445fc3ec0d0c6141c42b79c9a2b1b9d84d5e2ab18a383fce01b29dfbfdda769387dfee9dbe2bd71ebf2e49fed5a33ba92e496d50f49ed466e9c882a080baafa1c9f3863ced1a26b8b0c00b1c58fc0f835ac1b98091341b7f5e950b0ceb6bad08d9efc843de317b06d2ac0140b583a7ea033cfdec2acef592c70a58393c1245306ee90cf445f1cf681c49a87f27e465d8c7c46c9e0e1a3b4e95f457d83e6b758e648c620adf5ff0271c3d4a8935f26a9efc0e79875e16ba8215bbe800a665f5e677dcd90817c93401864b3c7211110e92953000b27add3667898a08c84bce63c4ef4d7fb4bb37e22990bc7df48088b20007b65b38d3d0c7eaf0d9c9f951a2303d836602d7ab83420868f00a0622a8da1c47feb89a186460e1472060c2e6ea88e3d757d83b7eb168d0f4cfc99edba31b636db538592572c8220a112318ae04df0a07a785f9034b1152aa1ec1a6b4bd205617cbbc67927d39695fd5c12fb8910b62491b2466faa93cd641bcc2936f757976c1bce56fc09863f9c57031e0436c1d7913e897bbf4738e2524f2cd119b72215f026ef0d8e7dabecd469d488f87efa706a74c1eec3344698637b286029148df5430e1f413f8c82628610f0b0d35a3788fa0bd34158f18ef86653f991a2961888cc5ed69e496b3867f205919ebdf501031b972e6e8708beb033ab2187868d1d7f7e7c2187e16755444279ab692385787a6c6859a60e1ca3223127401ff9f650b0a3898079cd1587ba6fa1aa7d962918aa5aae8f748bcbb1e992da9716fd8c0d8e35403f44a8c133440530b1f853c5e56905d88886e8022d20774bd43f8c35ce56fe4a2224eabe86c6a6e797827c3775e44d248ae5dd61740d58a81886a000249a6b304a544e06663e55661fc7b247fefd86ea5fd63164287ab02543d9b1604727b88f720a977c84152a7a87f6479b1876e81df8678a47e09d662b881c33167eef7d6d4593a1562a86e1b5f4d11e7a43fe6ff4d4b2166341f54f929c3823e6dd6a601a43c157f935ebacdba6d0f673339b8afa0fca847181e7a2fcd441543119b08ba939cbe6ada0de7200cdc4de32df89511c0be6daf3f39297d89f09d017719361f3dc9454b2b805f04af8ec4e1c896b040718273b0ad2dc42d5cd75177b37dea417ed1093b3be617b0a85636062ed60091c85eecadcabe3445077bc6e13bf55e99fe465cd54fb96968b57c9b88908fd3944cee70e7eb6f280282490cf6662e41b7a7294e689800ed210d2ed58e4e03424015e45e645655d5dbe6ccb2f017b3fd2ad07c9c9729e75fde604163bc7f53adaca2fd1a4cc3922ba7606ebf66363281be8414d90ea0f1cae8b80f7babdfe92ba43b6d426d774bf0a1de10c46ecfa80a9d5763f948818034db59b7d624961f238d3f9f3af2fa7985f56067aa52b8122089865e3dfbdb92fd075b56e1cb0966e0b3f49caf81dcc6de4b5b76c01eb7c00f31feb29b041824ead946454144e3c3fad87a44be7f264eb5912a2f0f70a9824191cb5f980b338a3af5a8bfa1fdccd549ce66b2aee8a768547fc2c80926059e5f29935e6155e52ca89df6752161639160a73f7a77d782ee880247a93df504aa655e1603f47682907347e58a94bf88b5ec9c60fdb2b1ad7e5af375a4871f330c4b3d363b8ca52172f0b408ae612b51e8c0b987a036cea2f56ae85257f3854112f031a173234524302750a7a887b38fd177ad9fd78478ef5eefb46175ddfca1887d5cd6af55a9cff0e468759505c1512e99e4b2aedc085100f438e97836a0ba1ea64da003c9595fa10be4df9e2012e2c26ca0d92c5855cd6b82af93992c1cf7cf543e96f0dbc1268fe2193b36756f0ed156236a0b2b024081d981ea181bdd709a1ed25f03fc506f64499eb8aae6346a53f8c0a9750eafb1fd507212674ffefc9ef8cf58c0fde9ae95600dfe6ef38969f5a0de3c846b620b53e2b941b039094c1007f41d88c657a8b3f15ba5662a6d93a109cbffcd50f042b672cd48a8459e15dee4e185c9ff95bc425d7e11088ecd3bb8ddd3818b6bed815791e5d4b0968ce85e9c6a289050c464bfed71067a3d8e9b745ed855ef42af025031cf06b8781a623d0cb00608d3ff8be65af583d8d739fabb1d2f56702674a0fdf6bc0937726ea668698e29b90d4bcd2cca44fd267e55d95e01ee35f8c76f44f7bca9e14a74e79653d5bdce6db5147561b74126d8f32d092ddabc88434d2b344e0c5e395d22d6a4c76b528107dad09f51009f94b6c7921bbc6e73ee269f796851b911e01dcaf11caf6ad085ed31035dd580533c9a3f27b284079e56ad36b5e41d109b69e9e3169a4e04ea3932f8afb75d9a9b7ebad4eec8ed77f0cb60164eb4f6b801e97e118fa822cb79fe9d4ae6054a30344a848d6fb2b7ad216eac1ef66cd3472b4743622375fbfba62d97484e86877b827353a01618d3a203fa7dc27353eb9331bfd80fe0f9f928883f7ff07111df3de7fd27ec3b0611e0f538c202ed978dfa5391ca9980285d02e0cb86375fcfd0cbcb0da901ce4d40ed1e2fcc53a363d7af3c2553b4202c08b840d631b878ea6da87597a31bae23c057ad1119db8d359999549aefbd6b3753a03147ac4be9bdae61ba08ac5d546029cec65e1034d3d353167638ec27800c17b28bfca496d65d944437be856dbae44a9672ed3b09241d67f2e5bbdb38ae9ec960263a66f8ff21568219c729a889c321a16df36a954d8ae15207f231bbf875f6b78042b166c3317b54efe8ea6b5dcd7e86b63f49e54164d0f9a82ed95101456c0ea09ae0181add85faebc212bd7f206e2915e18b35e664d13c81115627a24a5a004fb481a26b5506a17a0e38b7bc3507a8e3840e2ce3bb440a2f4b180587d6743b46a1caf45f8cd184c8f92356a49d645edf0c579a52f8fd6cbeb912d9c767f4d585e171470420ca05377e1c29ea19347bf083409a9d74dc5105a47d34778287cc0b864fbceb1e2688bbd259f17c51a84ab5dd6bceed0cf7f750a80713270c5634257a151ea18adc16e3e0500f075f2516003db1c89c1cd3a7e74d914d8be5d3a312ff3dd2dfc76a11879c72b40568b1e7434a194d863ae74c3e319972523aaae405056802481cd594842b3428934a40f24ea0b9a44993e3dace377363587099d851d928915dfba58a99b3980b6b40f77fb0d5659e8c3e6c4238d2e26fbf47d235ccac2daac5e4bafeccfa58997459849c54e6ccfbfbc95ec54d10f85d1b50ab58a377cfafc1594b5e31ed93fce72fbd58e97797d1a4e5e229e5b16fe73e069b970c88286bd81f84090844b7afe2fe1f7ab1a7e67e993ea740080cdbdcb1e99d0a1462e571d2670a52a6dc0a8c4da543eb8d1b720dda66a61cdefb1eefb76378a570a373ff9397a1a9bac13e86b215a5b4c261e8b4d057c1c02f92e98a17fe88a1f523b34199e2421d2891f76d4ee5ac038679c901a89ee9e5fc26c95d5861d191f1c0452f6c0bffc3382fe069bdc0937c3c0f05e1e2ff03694992fe89df5960882393c0ca09307d802647a483339b749103ac51d3848f7d3b608c2d0d2c60cab85b13b6209e16eba8886e8d8ef5813f9b08b97fe3ed1a8a6694b0037e08b909282808abeb470a1cce115fc55471a763969648008642016d4688a1abde7355bfe12cac72e8b65eb2b481f509e009872893914a0e6942cba16245041a7ede78e4c847e7878cf1e188134ace2b7d6ab99beae9acdb8590b4e291ba83fb4fd1fca32cebb8da86fceff1ae87699bf45adb28261e2f59930fa3a77e080470c8c403ba979820f91ed068207a7252c933271ff5509b7c2ea6a9cd5c71deae5d85720dd710afc0e31a93ff86cf198af022e4c611aebcd476b4212bdb4606cf2b623ee4619cc9463e68816b9460c3648c60d8d76b0151df05956f2ae1198045805233736769bb1e4a0cd9fd6791965d2edc2121ac4e01658de91d5ef1107e9063497d5f4ccf274f964497a247e48bd774337f55cdd843b1504c94ae46381196715fd2fb06e76465684e1edb10b7a426e3b75330e9207131d02bc36c7670bb13b15480700b8851e7d6096b3f8a9c8753b0950906781d37a750a2b9c6a47805d61eb97efa86ed9137b312aeb46ae7ea0ff8a054f806f798d8ef8870531b81391c6d8e88a2635aabf8d31b0111efd7afb84c15a15a274c55136786ee424405ef3bf5f68f48750f5a73d59351fb76eb95ab1c734f6b98f3bc6ef62ff64c37a39ff94ceb065c4751df53a8a5990018d6f55ce09707ca135dbf3c3cdcc544c0bf723b634c3a407acecca41942402d0fd4ad4442ed41b75d72bfac4bc50f3eed6a278e86df6deb326a241a118e91e674846c4b12922c0777e5d71c0a13c8bc1ad5b0f3d05ce860bd37f3a13024ceac5dab237d738fb1ae63cdfb94b8d0e84047c35a5b36efa6c99a7836a3cf9cdd148a95ad52c156e0fd7f0ff79c7aa3d6d009782a055760625ccdd58a79f44f440b86611f13c33d9303a0ba247d8bbc21ab430ced5e64a034b45a1f881940116a272972889d4897cf8cdf3b0090da5ba27929f232f7105e1e7a6dddbdded0833c707706f4404fe9109f6ce861189c32988bb256588bc591e927bb877b098b258153f5f924bc68c7e5b3c39e8a0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha49b5f2471354c0afd606ebd451533695d75aea4f9e3d753cd2e422b11baf25196466adb2010b378a900416708efa79016e6cbeea1a71ccdb5cd93b30e904ff51275c4fc87ae1e81b545342dcf52c1a8278ff9c6435e1a7efcbced512c4991ff7d85828dcbd4ca99c898aee2ae2d4416321e0661e38df03c6ba35e221192c6000b1aaef35bf00508b551ee9dee561f38a7fd32319b47ccf11f947a31db5a0cc7b0bd72ffdfc1e8d672a27ae1bebde73e1a5716b34cc95dc41e18ebf5640852e2260593875e65cf017dda6aa295289e726abda3ce66ff7f93e717e13ee5ed2779d6f18090377921527499a995480a2c3fe779f3b52c7729903f367dab33468bbc25a46598e8ee139943be0784eb3c782fc046161c8235314eda250fe777cfdcc48007516c863402f26d5610193c2b7ede7b14d411c0c5acb6f915ab218f9cef9e83dc801edc41ac93dd285a05b85ed28e1c58b8b8a78320a3458b25df0862cbf7a84198f171ab0e69f050a524113427dfa6c5c2819e09e56cb051e966da917ac4f7e68c9fb7c548d0685d221f31ab1552d279386a88bd31bc8506e8a53b61efc7f6707e2c611ae905c3f4aa50f11710c28f59ffa194613e1db5d981fe5cc0f9193fe54c2c0897542b81ebd0bad731d49a95da7a6ea32a1a87b5f4f878017c6d0c6578c5fa21f40bf2db39116b6ba1ed08f408c97512ab614264dd3d347886196af76a51018ffc1cbd532b14019528e66b9eb1c1fd6a1efb20b5ec25efcaae20f865a3ad264b675bee8bcddadd10a1f716aea762fb6aa68392ef918c3495fe26a74fab3eee4e932cda711d46839d4600623a44be94315dcae5c0f1a85b3b9c4714975f2f43df1e4b2e28a08b0d7256aee455531520228d8f6ad17ca47487c8bbbbcfb32a1b3c50ba2f3deb37bb68c8aa84871faf49add823622570bbc2897584fdc0d57a0948f65ff577b23d7eba15da138fe19671784ebf2aa10846b3e4170b4b9f1123bc7fff0e52dfa8f87e807b46903331d654b3e37c56b25cb0965c28425ba33bdfcc159df0fae6ed2f8f9c2adba01dac6def8c66888656199146823b95fe6406747d604e6df09c8036c1e53cc8930bd3bc9944873f07190d15304cbc4b8f6d082d4dfdaa1b2df205335c94aef1d2487e795835147cac2b428f55d20cde5a6b1eec2fa3ece21475c97fe00d3a2bdb121d3c03cb9e26f70fead3c67af00506bb8df7afb233a150f95be84a9152293e9c70f0b07261f29bb7f3e7b2597978271503ce52850d7b20d72a031e1168203dc63073f1d526b2490ab047b99bf6e73a3b483cb5ac32abe5f5c8f2916eb03336e39aaab4ac292603fd77c9baeef90dd14c28e1fa261acaab12ef610660d8dd04a27b21690872f6f04fb918cf8ab8c11259be5cc2be64832f348105f067aa41df3238eec64febff786f5e315fa64d6cc371596eee0b05e446bf2de0dd605293536616cf5bf6dd1d6a2d60a1ab344c064a5402bfbf9f4c425fffde4ff41af0d0e47d311bd5dd8b2c7edfd0cd3d9d9509503bde1d181da6b07a043ec15bf4c0a60e51f2f26584ae157b66e24311416a0f359aa65d682701291bf0a5992c17db1879f03406fd46b65aa17963eb300c149d58794d57a6afe7dbecdb81e5a644f95cbaafcc5e0bab13b7034827ed77d9e4464397255ee3b6a520159add7bf4033b6f3527f2e29095281682a380609ed477292a7f3f256315c453093367898a4b23aa60bf03dfcf64a009f4eb16766e0cd33e85f73ba3730b9a1cd4acd92d2f9914ca9e8c88921e8bcf8ec430b43791885c47c919535c8d4aba97383ce4a410af375308fc49a2bf7858c4560465d9442592feb3048b14f432021d3b5ccedfd69cf7b50a1774521d3b8e265d74c3cdc544d7709c84f3bcdd533f31a5c557502b0601723272eac0efc3abb7e6e431ae8dff71539a7aea224f429039ddce18fffe54323681bdb74aca12416540b14cc15236b89c44d0b12842893b5e8ae2e92f2e556ca1fc9dd5a7541794e0e6a7971203efd4b9652e4dee2fe3353c0accdd097b2229acaaf1fc15aa07eda16f0d91ffdab2c493da1277eee11423bdd2743be01fec9a592efbb7d77b8d013f6c34bdc95f4ef87113d58a2ebbe678f13e95b38a6c6999a9e7b68e506f22344a6925b482388f7bb2c80b1fee077f2943f0c498ff5b43d89282ad7534a44d209b7c2007b8b0cc30e91485239213875964dfe9543865cdc0129a9af390ec8ae7281954cbae3f0ea1368ac60ba7b941f0ccbbde7d1d51b39f757a23916a73304aaa607b91a51e03b7a33ae566d5b30c73079257b08198b24eddec1efe73b80f2aa1a1dd57b6dc44138a6b52b15be37b4be3ec37c6be09e76415cf9a025b519e4b4bed990ce1ee5fee4584f02afce16a8922829098759773be64893e73325cb702c9cc02c5b78bfd8445ede8183b6895a94db3959c555fa7c4ca6b3662167b696dddafc1be0a8740349d3f081596cd0a2eb5ea9ebe1bed309ce8655fb7a7709b4cd4b6614987ed73ab16b41360659d931da14e7dda21a1527c8d906c07fa9ebe03d025c4cab3410a85a4de475b710568415f1e718972cb0924a1199a732a13bb150cecda2b3c572a30d9be4b58d4d58a3bf7ca12882d04099028e9e7163bd126dd3a2200e42392a0013ded77f4097d30eccc9e05c882cdf10d9f5be343010d437426103698433e0e34e0f8e2ffdfc0d20fddb86cf7c1ead6a10850b60e803c0d681ec311bb65087d0938de125f058c0d6cf3286e4b9ab56d17cc6e9bd19996b974be136fe6fd4e54f430c5e1686d546c341b9ce6e14a74408001af4ccd86977d84a370ac09f744f2dcad50e5996594e9d0aa510045e1240d6ee56c3899371cae400ab1893da28e900a32453ae3f51ee7e419448a862e73a6410deabd81005c49b123d2534cc9ceb9d7bc8d6e5368e20476d3a5be73253f24d4504b40060c763077b968b232fb34063b5b8e9eb00702bb5ee4a8c91e441461cb78abed3f5419afe0988fe2eca70860cbdd59f9480f9bd13676d9bf932f601e1243554c0456cf82b72d1c25301dc6c0927171ef7cbeee839c3f0426a2d1c16a1ac242892397444a2a3373335b9ee22bfbbf2296140f097e5a9152837c17f8993fa47d3416148444b8e9e5030970c7f9174b050ef287cbf824e5e3671226c523faa569225b384f8e9dfa19a97fddf05ec86c43aa20bc649be389e73a4a4ccf746654feab48964b38e020c8137e1fa2e463b7d20beef8e2623095537f45a2a7f6bb2269d54df688475a9b1175c2444841f160dc462645bfc63b6ab006896775826e2d6d5edaeda199158ca94abbade4f7c8887c5edd567f22f5d826114fb81069cbeb695ad5627f5b9b0e7e2a1fd35235f6c940e7bf0e34751d3941e1b9df3c7688e4a5ed556d74c37e2771e8884be4dcd7f460327d2148afa48fb4d1cb9d21bb592a5e8230f74e01378ab67116954d1238ca73584035c56d009fde9fb6d4233faa862adb7dcfe0039cc43e66431646ba666bd27244026446aebe72580502e11168ce26b2acb1a1dc72be1d163fcda5153f79fca26a5047a038ce52713cf2d7e9f4911e561bc92e9cf1d6747335c4878b3b98fa7c026b3a395b45767c2b34b0e75564f43d37ec56536f4258cb5dafad9bd7f447419804af1c73c68369c56248e657776bd4ecc1670706efc9dd9f3c90d7b609887c97bf718b9e975d05d0245a9db015c33854942bbf0b24e06abdff19bdc7b661d0d8dbda29b621c7fd0160e35862f93e37114de537dbb825828ae4d920c632c024ca75b1160f6519ef928a54f1221947c5cd00ba1a1dd646ff84a97d87003014b3751b36dcb5f353ad536c7fc8dca8daaebfe6cd63c68c858db34329a7fdf987b15ecee39a579b4c98aaa48442d20fda0e9cbf75a82691ad6e3153e55d6eb8f68aa8429f0a3b9095c168e98f6ea6b6fd9c0fc0557aff8087f55fe69160c98aa322e85723e6f6d19b1504343641c98f4c526bc166b86b13968f962d1a5807f3e712f9f9412bd8e3f85c5e0dca99ceb23d73379f2234c66c782be46ef91f86d435656560c08d37afdd85fa21a7bb9218307ca8d22117300de00f97c983e33afb52eb7b74d801b094593a9f84436677b8a0e396b63e26cff877f3b9f1402c7a88d09c35e83adee810225f11ca79653825f2d52ff3a9f646de7a7b77f70a969a11e7b3aec83a503469e7aeed1cebaf88f9d8fbb12cf36a5ee819a01052ba5ea6bc42f0b5a16a66471a80f76aec47e72eb1c8e22cab3ceb83925562efb0173cbd2661b5e36dafeff95399fe64a01861882e8229e74ce4d02e209efa638a8b4b9de7ec3ce6297b9c6042c8bbe248ec1fd269b731d23eb1dfc0d5ffdab988c9a79aa95e39a0ada39b5e83c731133d9e27f42aabbf7f135f9d7f2efcbce4b751ae051f0662698f1e7ad06d4d77bbfd72ea4801be0509bc5dfee5c316abc09042d04831bed7c039525a8870c67c81f884035f2a00ca5b3d00d02401f7a833f81f4998c8ac8fe2ff0dbaf61ff04381da8930b235333e3f3786c4d10b2a55a13622c562c4a2de6ecd3d2dd2db58da4c6fd5a736c289f83c443d0d3d6921aeb2aebc2f2d808dff2d7ebc7b0b1ceda223d6f882fa890862e38c228eeaa69dfa3fdebe77e468aa19303642a9ffac5cae74af1bf29d3722af0daa5f70ff9e87b3f1783e2aa252cd1f41adc894886efdcd338da5d665ec744c1bcab6cfd7475c2443dd7228087a1e23acb369abd69b86db402169a1b161096405450ce2ad87b733ff64b0f1c562582c9ee7cc1fc36493a9d6154e3d4dc5d6aabad59a87dbd95276624ad6b9bcdc124a9568e8df76455a0363e4c4b3e3ad2bc2fdac2ac33a5488e7cd2cf3ddad7e914ec528427a2c9adb6626aea8b1196de0d186ffaa3dab18625f025447f487df4b4e62b15d9c02c23a92ac20709463fd71f0b452565a21a26f28f33632e10385525ffdda9cda45988f24841ff182eae3ac22d1eaaa12af52b89c11497903e90840f992022ae5a930f0fd255605be6a8cd97d77f2ebfd12f066c4d790d45a5b114520931dd88d3779d4b8cad843b9d1581a82bb3078f0de423c1075a2a97230b673095733841adf2eff2e701892c9ca581cae6283dfa88bd0889cfb09a1b7059e4dd60522524c1d2ef792f71c8f25e4a46a84d2ae45f694a42954d2f906ce6544a3fd3f34ca72909ddb9c56f701da085fc826d52e6a5f2d9248b5f299b4e7687cb16dc8432e8ecd0c6997839344af13429e5397a4dc3b9aa99832d3a4cd6fa8a4a07f2050b116d0ba65025e42a7c83e584fcfa300762f5dfb7a46fc3ac2054f9c695deb8f5dafcdeed2b8798afceb63f82902b529b4e901ed6183cd51924d2ddc028d6609ac25c2432c189ff043bfa6eae9c0e6433953e7fa551c35714e547007f05de96c0fe9f58b7c9a25b7b332c6806b0ae1a2eaa86da2346e2bbfaf887eda3b83b5eb2d2ddd4667f45fdf65f3b260a4a89354b643216867f2259ea246d83f65cba0b4c5bda1c64f68b7da138e1ea0965132a4352d9371c71c0d0c0c5c8eee250a1c4c345936f49f6e3a47db75f3fecab01db63e3c7cf6d4cefd7e7d865d974a154eeee17d0ebe421ea72992b0285c5c76795ae2806392f47c496fec859c5d49ad78744ff7e5e6a562463c0c611b7c74cc645efeb0087a126977c8c442a18838bf3fc03f6dff73604f271ea3419bb2ef8e7115dfcea4f07644d9f308cb4b3f7629d823095549f101fa3e5af7b5c550c60892fb0fd38ecdca607a999a70a704b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6a1d8d5f86c53566eb4f5f5117903d59c2485a5bf577e58749b4a2007ac0a8528f8f8254c5ad27f1e816fe3a0c6cfba727d4697e55478bf17a1c3ef26c7fb3391d98ea4ddb185fb2c44e592812a72b73d49db3f4956f8b18c672afb9d2f279ec9d47afa6581bd9446a06c961a7c0f48f7d372bd3503d69b6f2ebc621ee5b8bec05aa47baf9ae6ca26fdd38a3a3828d9af1b81673651a69a89d0efac8c712dcca8fba00f9f192f4fb0ce1d04a0951d7c7edb40a20b7dd2447091dee6aeb1d45d1521669c6a8c4e5586b680aa6894d59c6811e5dc7bfb28127a41bd53c793c4e78fb1c57e20afb1aed987b952963f22234100cfc638d8d74252c1a5515ff389be66b41f00ec5e8e6acf260702c2eea4c2eff5aa94d5d87c9cf8155b47e0b3b1f48f0c4e9302410390e53d8ee904e87aa1ef057bbec595cc50189d73afdcbe57a48a0bc7f72da52c0e04d630bcfe9dd88cf56b583ed1528711d10d3854a0087028d45df666ae6ffe89691e9c79098216e0502c3da600cf3c94919ccced66403954463161dbd32e235f172690af6cb52350a2a4be128f2cacd582707473b73c59c5631941a911135c7a4b78512515f952c46ac612686e32e0d2e028a3033097eaae9d177e5d9fec6b0ffc60d43224b25fadf2915c6cbeba4549cb037b492753e153ff805e1329492b755c44b17b37e080fbfda46be620bdb47128bb3dd20183d47dba87a4def84855499a310bb30a30b832fecdd0360f7654b596754bebd087578519773d411620fb57e5ff33e8eae38e0db909547ec5b304c2aecf67116950383e0bcc818039d5ea2f1cdeb6ed22605815579b72e4b91dab824560e7e5d4d6209d5bf084fa56e0d4ad2da9ca90f86b48332110615ec029e939c6c1d369b3be402bd365fad49e69fa851451ba5ff363575322ad785f18437655475af53f6390e762a027a867f38ba1a298b18ddab2b5eb3a0651f0e202255452feb0887cc62491a12da92371de9df777b93683a9b3e64cf8253bd9481716bfe4fc4cdc41e96279dcd195398354c6d68a48b0000c758c8056f360a48a1400b8aae6c8164343676f9b5e3a1e5a6e201e0c4627fb2687e1a9d997f918301e32210e30e36eb4584919c84cf94207907d683673d9469c94b5b4c3b3fec655851d58c0dd1d10a0d7da60e9d500ee7b3c63bdabec99262699850fa82970f719bf2949373ff73607dbfdad091ed5639609bfe9371e6b6f8bafad37b3a46d94bccbeb4303bc267f7a8a243b7cf20690b122ca0af41054b502bda00a9d41421b818676c032bd5c500a343edc45b812ceae28149b86a8757dc69923bf9fce6b7295e88de79290a8f26847a5c2274f79deac96ff29aa982c101bef276d032ad6c4822fb0240578692a353341ae3a9077ac2210acab2b7fb83ef1595a484ef825548510cea8e018ffa0654ceba319a003273be10e9bd4d6c745da9f087579d0a160c058758fdf09abfed327ef1ffbb809a966e99258e5f3475690a2019401c57cb533abe7fb9aff48c1eacf6ee2f37d7ff0548697ef2245139e3bcfcd1bdc05a8b69549494e9bcaae29e1e201c3d7fad25079bfeb20fbae9cf79dc997e93e01417177ee8cd5932e849f55efcf7af4b9bb8358b8770d1fc0eb3040f50052d308b55ea309a17913964ca5c6889ec4af5a97580e71eb82e113d2928fcbee0c4cecc4fd878a38fb26f72f2535e8a6f429de0a046b6e7cfdfee000176de39461abd946cdf953893ed60a0d87c7769a09d8dc75dc152436d3b9dd34c0094fcd5a72ddb12471ffcf2f1fe6fb49e3aee53f67057ff44bbe9f287c68dcf22f91fcfeb6c35e6ab3a73ea9228834869db71705727d96b4e9d83603f6c1ffb6a1d88f854c3d19e27e5c1a4dd305cb16ef6f7bd7aa0ab05fe963489d1fb4aa74764bae033e9367d58d88042a23056bc5dbd7e7733ec653315097fdd04cf43a8745c83203be31f8a7e8cc55db468484d95cd148036970da2feb88ed49d22ce91c1a88ebab0256102e25154fd2f0198fdc7b99ce6126cad9b071c2bca1c6a5d22d2986fb4dfa24fe02fd84ed071979586097af8ec111c4d850f9ea7b56e48a90a70735c313d1ccd34acfc4014391ec06cef2f3a9cb542801072bec72a2ac03230ff3ead859d5c5f0809737ac96f6aa48f9e8a47892b1640081f08fd56ed55e9f40bb5bf9ab17255135a9c1823ccd707717665c06bf64f7196b55e8fa482a53780d0505828f8e5c070b05c3f5399220d8e7343855a3598fbc0d98c6c835a2fde706ea4ae6cab8d59920a9462d806e0765661787389f7c830e8dfc82df2f264034415353fc1e057b847f14a7c44cdd6b5344c25fec1c9e24c5981c795f3377f5746b1e1b55ac47377cb6fae2b7076a7001481bb28c8a78cd90b8528581436b727c9d15dde0b16ba743d5034775e4b036a7ec99bb282b609bc63e680d2376372712bf6392a86f5e8c3cd0b040d3002bd2e30ea26a92540f391060a3a310a114dd04f96c4d8c261eb99905f3435a64297a1f7c7ff26456b4572d55c2e9762860955edbce93a59ac22fd6830168f5eb841ab431c4cc5955621f75eda0fece7fcedd9b59f55ac4e669845a0683c696ea5e2603d8d31df1bbd94bd3c01c5306dad57289c1efff806d3797e2636dae94ea1a81c8d7d23339682ec451db5c767c3073b84c0d9a511aa2a82fa14dc4137ee95bf09cef6bf536d0c3832b6fe46d045b548988fb43d3ab9e66a04917adbb058e5fe2959f80bffd5e9333eabe54eb86394cc959623b0d0eefabdd44785c69e7ab38a041d33e3abd78af69dbb2f0e9eb5941c40052c666cf35be51b50d3c29bea1bea8513832439a6be92df60ee09a0e0cc924c63ced12dbbd7b03e5a832a7c1460ddaf73cdedd9082cd2cbfdc89ec8cb4cceaee04d877a90af2e2b7e528f282ae29ea3309e7cf6968ccd7c362247c1ece7b25987bedfff2915b5ed4e73b461771ba5f5fc55cb68e71941235ea212c0bed9f70eb1d1738e94e82e972a3f78c62097abc23d658d2699b429b2beabf19caeda380ba458d3d0b3a30f9ae348ecc09c4005fe5ac011099c0ee9318622c765217a67ec166bf426fd1425c1fc5a28f6ce5eb82d23bdf9713da8e98789edf934694a1b26381bb564ba19ca431edac87294ef00af1a9eeb882fce31c5d93113c8d3414f79129494f40e7aff2e955d999e95dae3789b53c4e72f1a7c500c250c984c295dd186e5fc609ff7e957d9dc287ff12d14f86a81ea87889653eb6552202b3682a457d94132ea3ad5905e9d34e1b94276cd2367e0150118d47a91e408137ab77cf61e37f5a23410692867b8c96bc12e2a2f4555431c9b6810979987b8fe607a6924bcbf18be96e5b0cc0ec9f5d8ce0b5d77a6d261e995c41cf83c19a6b063af3ce9814bfd424b9573d3657a7e4b7603ea21e3dc9136040a234fe48d70ad5fc9ea5f3f64b6b8cec344e6b6faf9ab206a8f6495638fdbd89907252c2603110e8b802d755c5cf9b2ddd851116da7f61b5aaf28a194d46d89c1d87b8e7b33910e308fe944d78379d2e3a16a38c3ba44d0edd682f320f074218cb0688e5ba5d63fe2f3a91b0da4f5a5ef9a39025d7a19a5bd4bae7771278c138c87ebae64b6020a37e447c934a2046832b2f4cdb5330695545915efd040add666967b71fbd17276e5981c4cc5b39b3b20c91dc033c4882418665ffad27aba4962200133e87de9eb8ad515708ca26cbacda08780470fdc3b199fef2d4380e31aea59a08a25ed27ea2af20eee34ac273ee36a29bda6de67423729321659f45ecfde9c8a50716ea3c78a8abaa5d904102ebf01cdc844cc30ba1b9ede7afaa10f31284cec17735a9f7c2f8d6744e419227594df494a5b5ac3b173c3bbc35e1f53e3a09725c5fcbc98617485df7f1ed0da377e03e653778f6744effa92da1472e54fbe9c80ab6f7d19a437614b8de47551f7db8908bbc1bd604ad5fe9fcc72a4c2b1349a2ff5c1bd977e43bb363544da31631d799ec8ade90ea7f6269e37db68331c463b89b7e99e1ef7b92cad85c603d6c1c34d8ac689b6413f211d6492749693df41879f170331d4ff49b4ae1705a87c977046cc1278dc567480f53d58198c0f3674448fd92e1e8edd8ffb304a946f57b768e9f9d2354568c37fa0ce534915245eabdf0066eb24a89b2fc6489ab405b6a59cf00b921ed06634b04af0ac0a300ffb03aef071cf51cccf43eeecd80d7a4405ed37f39b836609c6a70b0cf12583787cfb8d4bca3067cd2502f3463e851364ce602b9c6eb25458e5fac90cf920bae2a55fa34046036b3a65d65e56fa47ba0d96e856e748b2079ffa9caf3aef50b0e59476bede77b1d9d12d48d1b51f312b1f88c57636c76a27195edf458d99ec2c973151fa6181b93c3c6b38d53dfed744cac415dda47d4ef52257bf72d77218ef1f0be0346c5c0381dd27a1f4b6e3694744bf1f4f77ed92e0325bb3984e115275f5b1caf66e22a480346ccfb01620c42a8ccfe17e3853eee0e570f365bf87d94d95cc631b4615213d222a05fabc45139a29c248a61a1bf40633115dceafcdf3c8bd9446049d2296c2ffbaf90f3e8d0876a962678ffa5438fcf4b75264fa50cbcf907f5c9c0185f96dcfc5a07763f29c1ae5560cac3581c3d7f281bca9092fad29e67ca9b9f0e00f8e510d1f7825c3d342a7a754a05307db21a44409239c090e95df59c8768034c88caf5bbf2e047ab85c572b3295894d4e5a9b76fc32e3866e2a7a947264c0c5c7724c805e37d63ed230bf10f1bc736f1a2c5def3e128ed153735c54ea8dd06d31ec879ea5d977070cf9401979e2f61e1dd5d74337f6c1ca2f32a8fb74718a8808eb4837a208636eb7a026c39924253157146e14f887fb687ef16981e365c7089b502a4c5874efe78a5c2ebb918485ae1a6fbb55bb15167009696540e03a84fddbb866110aa62003dee063f3351c11a62b65b89b3e7f3a12d26df3c14574bdc24a5e9130f629170bca3323f562ac462b27c6df11042f52321e7030d1316cc38c545316a81a2a139b3629b0ddd3b163778d71c2666d03e7cb6c048ccb81db2fbce4bce3fbe5493d3903bcfaad833cfb81572157ac48830af30fdca197e6aef2761cadc05da7ff9430f342b230b0767b58d6276791929496f1707adde1af16b5da7d167fa97224a0cfff2dfd666ae3802a41ed7cfd8f09c4a920f93b00ce23aaeb27c3ebbdd62de9db6bf3df86140131780eb791c1b346181db6584d207a90a65321c6963d38b426340f07cc02c96ca33830dc38d168576c5d7494716aea77f69efddc884d247a0209b4d6d2ff0f77fb9e7ee444504321e0ff5f94fd05f921d14e62b6d07d15b8d57ec6816cb06668d3cb0afed1c31a245738679f0b8da7133c1f3797bb403e0d90076235eaecac1fc92b93e89c0cb354fc9d85a75fa4c925e59ef9537427db53e09c93d651f8802341fd63f206b54f98f828cb196b2ef7c72a274b4e1e604f8d3dfd7f2de9b5dfeb4831a076f7e0d77748c4b36f581c2ee89795174f664007542383ff7662862bb7423b9111dee40967390f5e94b1bdf38e427a9a680ee0fa54c46d625647e53ba787d5201723136c1f997e13ff7afbdfa762e7a072653781c77b9e9d492e3b3e192dffc7172ad3b5f000520aa868c2d1bcbfb30a4ffc4af0891bc94d963940dbf25cafea0956d42bc290dcbc4297a0aa80925b7be8664cfcaf40af44d07ea4ee8f0c6c6ebe072064b1e76e420cf491f9a5569ee52068e8ce982eecea7d75ed2b67cfe07e2f7f7d3e45d6ef4db4d788df0e78;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h46d6021959d5e6c5d15d9f881957b41dd2a361428ce9ed479765768d69474f71b214105f1b1df3577dacf68197339e9cb7c02930014f55085a3402678d83abdbb0c865ac7ae38e1d5f45f94147277c5edccd285adce7c73f5b359846ba51cd681bb5213d81a2ae11a37822af3c4656f101db17f564b79496327722d7528b6eadabecba55005aae2dee62205bf2d84e3c70a15fd82ac00fbe543d9c817ac8de335ef02c808800183b68bf9dcd3c6d01b30f73d4be59730679bef1d6e1d253c676f456c81c33311defeb62f70c714a0e7d8be1960936452f175e6a322541b1d1c90c34a7320dd1d493f73ef54a7ce8ba1ec94fae60164bb3dc6163af9ab2dcfb72b19e1cf1235716b02162f92df7491d1ddb5e4b8e15b543692c695b6b6d86a4282a3d9c694e7b953430f4129ce133f45b080a053ca55a56c19d54a53223972b4fc4fd3f5e38de99e85678d286b44e1245f3815adc12d37530a1d13e8445c74a27a1212d67e1237527b25f4f69703ce84a6f8e4020537f26056fbacec035709e4ad41f5d8351c944bcdbe13775c6612b9b052d9cc10ccee151b07f6e3f5386220a6664f874789d31fc7e2cd6694feb0cd5462595b3b5d72d757e81671ee3b06a33e833ccd483e95a58e28c4a82ce5795feaa30de848e2c0eaa626063d2a091c9bc82bc7ea3c701e0435a0f43c18cef51bb8e9c4cd5a7d11c7451dbb58439756c2656fb2bcfc430724395824b1e612e3b9a5d335b8c9ccc89a02aefce6d4c2f468788a36585be48285ea800987d7e97ff7691780d5d10d5f45ea0de47e431cf4c428c119ff779b61f3550690013dded55155e9ac64723c8351af88bfab7c34fa752b4fd2cef37b3c2cc493f03dfa7f450769a2859d750c5aa8d6d942706887ba8d38002585d3a069a90338a9471032b235007d596b9b2200f56a52a49fb054fd5df3825ab38cc16d12041bb922924e4564b64aa48d9408fa5f16b9dde7cafb786ca6ff93ea1f38c6e1fa82041fe4371e1719bbcd718e0326e2a2950f0681bcbfa5c23c18fe1c20fa7c96c1a8bbacd6be9501fa92f812a7f9a2d4464cfa99bc1e55a527b7ca5465547fdeca08e105b2860e630f0d366b686a77d725f37bfab328d0dc12ac0b28b3953a44d8d0e4fed2ed77a4cdf1168f5e5bc2b1d1adac6039c729a2d6f7c09930b2e9fb802d1ff309a68e80ad30081c326912da446366b4c331c0b2b706cfb67530ac8054a2c897d1516b45a6d24a1abd6ab86ddb86544c573bd16b9f983e476cfbec47d51d902fa5deab534cdacb38045a0891816c01d1ad43e80cbd62d1edacea02a8ccb750715b8ac639ec01482b2399d66635282bce6ae0b723b68dae60bc5d4b669c2286d40e5494fc3b0c6e42348975d0265543ccdbbccc613941a1fb3d9ede89e0eec3cc9272bc95b58d5c2f233c6d3d2baa6d7000a071bd7b25b68af3782ba7d9cd6f9ec4062c704144bc97cc2fcc640f7e1912b44e64dcc1d8cee098ba4c12d1fadd8da115960e5cac641e172bc51f0eba0671fe4dd7e0d9a1963dc17c1d1430a399444d2cdbd8a624188f6d4344fa5ef2fdc203dc4ff65e3aa16aa6b63914e16f5d2db553a5a937330c31e2afe428ab75618d9ab421c15eae783bde266add16f4beb4f5d583a8ca4d6f795acee8e795e5a72ee9ff75fd13c2b97af448cddc879b74a6b25342ba32293149f33df63022c6383f87657290bdaac036bd9567f702f5e7aa0c817c3322e253754fbace0f0f60f85cdfb97a682b3b8c0e93820b5ad45710df0ec57ffa5aad8a28de7f6a8ff77fc686464730f06b3c91cb2dd658a577cff9f89f5b997f4aa425e03a1abc2cd3ea034ec569bb728a3f96b7e5cede8ac78970778db6072b1a9be8ad8e41a45443f088755478d67c2aa3709dd026b16c0b83ac92f28d3ffba3500cb38a9a1efde453044802162040200e2cda7c018a4cc50f9021dcb53af3efd1c525f277913f8ba4165a5c324c32f2240f4750c666a9e5eab5236bf1118017403dc6888293fd4d711d883b42b40039523a4a3e598f9df45c1519544ef38301856af1985e6ac9bbe3ed9c8db43fcd4928d80101fdc0a104c761f2952c75ecadf57ff453cdfebefaf839a3ab9117fd7a27a1c6e7d9cefba942a310e124b87cf13855c6feb686f27d487cafd181300a570a2f1a5e8970dd0d56c45dfc93d9603cba409e998e80dffa0d25fc6a193fff10b44db304ee6ccd696641c7cf92e6ad53b8d80592b6c4252e730ba15f50f769f2aebd2a083bcde4f5abbe91d10da0d1477cce1249de2b51691f1167c1468d14cef31256352f9f8546d24dbd49c986e037f5318dea05764fff9a38de1084a3fa0c95083511becac2b5df93a42403f642ec18916c176c37889e33f8d77a7a1f233e104d74cb57f69d27d5adf4cff0775673ed597ea234650a75802bb75057d4a3b40c104830f27f9a36a1da11d548bdfa4b649ff49b89ec24b782ddcae3eabdb5fc7f5e5257fdfd0b29b9b37b38dfc5eb51cfda5ccd07c0196c458513f5d935636bda3fba047cc021a18421d9cff50e7db2a74cecb27d6a0820eb6ca64045a5d75a248a48c270a67427822e3eee3f7f21bf8bfd232327b4515a832a1ab7c903bd7f87c754e0d41bdea3c5b4122e3fb68a28986b9ef5c7570dd536b0d2d85080999501295f69271b1181b7b1af171dffdd13ac0ce68a3a22ab710583c11897dcfcb944db2ffcecf280f6b78780749ba34ee81676fcf179c56ee4644fc455337052ac013fef6dade7d683b6f672c1a48ec1b1f03efb2182fa7bffc36830a4d06c29963199b9e80c59a1dbee2ec81937e2d54b22793adcf9c6a3fdf12df9c746ab40246c8e688ff71b0950667239269764d222acf88609b513763601605237db211b6093e10840118595b7c11a057d3bddc9bf7b0dd95ddefe8a7ad019deb1a03394e058b4448bff9b45bf218007c4fd8df73f8d5aaa7bff1f6a6c04b5d3b4180c8bd23a56727a6a3fd1b2c8717b6a703378b81185a3da50ddda0a441ebbd6924d0b9206bb50f2175705d4ede816052f88aeb1d680cab7a8186b90553bfd3176c9acada25d8f67eef3f231499d7abeed5107b2baee2e6dee0be1602d1198bc94420b91e531e7c738baa0944a95191fbd237923e5ea856b3caf7e0b577d9e5049f1cb8332cf4198a075cf66da6a83072d744ae83576522d1d126cdf8fdd05f593002184d3e25ce8e6d5091d6ebc68e89cf99241eeddd6dd7bad5ff051ba13ad1809e6b101c5e37867c50dee15d042b8c7eaa85bfc7775bd0b13052fa5de937f4ac45a3471d2be1a0738467402ddc498b417273b23df87fbd638ec27ebabd30b466c9b8860660e3f68ad42e57e4304b04cb3a4682c1ed60a182587f302edecd19ba38d94de61e080eabdf43b2c58d8cc5ca7533d88f4a3ad2661d935a2c60d4549ab16295e841898c96a25eef35c0280785fc06f94996a9deaa9bc5b6c30f6ff42326c580b00758f138c92321f1e0f079c7fb21d94d62f146ad62227046de3bba68e1e887cbd3cf65c5c5b3a694499054a4abfa3d0f22badfec2d2d889cc9da382d33cfed1c3ea58ff8f561fe620f569383851a6a8447a86f86c09ea1f0651d06ce10fb0eda188ef45a0235a64d0d244d89917bcf3b8ad9fbdbc6a24cbb9439b7415f7bdb0ebe3ae9c4e6d575bbeefbfc85cb8a523c78d01983fde19f4e45c52239a9ad3b91a0fba17f034aba55701ce331615f5901185384e3bba9339fe258ca6703f99dbcf6bfb320a025cd5d998a0d3bdb849215e5e7042f52770479ba238fb87182b314d9bc90ee6b7c12be142f187ac4d101ff1185d12b8ed9288b2f4904903275be018cae23e3015188c5d2c1ce426b9f63de2447f57e520ad7a35f2b3807b9fbeeb11fb10baaf0d0e374ffd23376ce7cb91704734468b93a52e32fb4015d08cc843b4cdba5f0748685e41e4982c474c6f492eb87515608ac39d02abfadbfd84ab0eef8592029456ccd8bfcb6522bce4e0a4b41dfafc7eed24a3c0789d7f731b7e577368e3c87c2e715c536a5d3784c1ab79879e05993b17dcddc4d22ab84f72e0b8de51d84123cbf0426a3459e43b69fbdc7bec4b98a1114efe2df0c1076c4e393f992aeab7a9692d9696a982b758048cb5d672c6eaa4af0ebd75903de342d0dac4a22edb803b5614be12eede034e230f699f6044e8fae155bbb5937c92ac254a7fb74f66cd22a4ac72134f94eba5046393764d196b9c0022d6776a7eaaef7673131c287251b9d420d4569da7132557802b4b7c3320be1a45e041c5a8bcdab623443c6be0a3ae2ddf3a7b6063d9a8f8800f89e1bf9b3c3984d987af12aa6b8c5418ae29177b807b3ec6057c5f4fe8f58f8ea87816cc6910090d49cd5eb96cfafcb039123184dccd8c20a4b37fe30c91c699faabc1e58bda766d631cc6a6ee90fa4883dd89f38453e2859c3f702ccf6d8732000299774b94477aa77d58a9fbb88239f4ce4386102b9514aa519b2491d45834be7e2fc7975ec922995d3b1d6c0721049169ccc2469e00aa93c0c60cfccc492e1d5820406a1bcf0bcf36f8617d0828ec3aa77458d3107ec7409eb009cecd68f66248cc4350496ca86bd80fce4a1acc42bbe972430f3022a8e38494e15d18eea36ce5f6b9211dba8c77af57a25a860ce33c5236c3bb2b252993fdbd4a2dcf75c22dbeed25752ccfabfb39dac6bc845c4cfee10d63112a398577e26fc8f6e727508ef25f3eb968a33c1a0cf26a7ee4a260ce750ad5865a4e133884f8b7515de60ca570417d4779157e4f75bf883e8bdce7d078942ddaf909f28636818642c5c2c8e312e05a7ecbba3116b551cf016806f2d623429d560df27c845007bc1b29771361adaedf496421146b9d8d9f27ce213f32ff6167ef17eb6bef3490f9802f1b84360b819cc75e9018f28bd710e6bbf1bbde9d2f6ea46f7569d25a05f64e456a0742a978a42272228cafc1906ad17dd0564b00e09258b4b36e5380336c0765a795b6f1ad8c1781f7f45b4384e168702602f1c78828cce9c1531a7efcacca48caafda5202017c6b267310391ed87715dc174278741d6cf538bb621069465d7435ef9de609ff9e526d6e503e74ea0b277aceb6bd58a4a7c7ecf2a85681e75375e2999bfd56446007252730721e2ccda5d18babf709fdd79705ec0a0a5f9103c2e028dc00db9e612e72cded0cd00f07b315088e425e319f179000ddf69a2b161bea729ba65fef054822e7ac91c828f64b95671b2916387407ff9638b32bc7ac32d51509350fa9e3e8910f250b1f02f190fbdc09cbba8aff1a12f5dad6f895b4d80e59ec66335c875b226b992a6409ca7cb1d516c31b8a37dff8f3116a294b9e9abb97508c7f51474a5269c8c7baa1efed6897d125fe493fc46acc2cbbea27f5300cadd3aeb9fda988433c515f2cc9dd7c7b063ca974372bbd42a033c039a81c2d6b80a5b1733f612832500363f1461a8dab717b1a32c4da75bd7ad9c11381fd3e35ea857f5c5b99637ae4874531ff8bf3454e5e541acc7e8b739059c2f4a95b33308628d215a5754515c4a15407b42afb5af1f434d71671fedba70f8d503ff4805ec7bf1376fc2e5946491557282059f0edd3024e2b790d4180a8521845ca8682fcd3cb374de176d35172825d9fbcb9f5ee5b5326a9318cd9ab7f555afc22109f6caa9432139e4a18e3686f715aa5dca1e7e5332275b206f062a9095636b009aea6c948346f1d5b9b48e605c8ab95c5621c51ce70458699029d3854b4a308d1d08a08c4e686c46b77e4951457d4d470c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf930143644559a1fc9d64badb6955f7d61913f87d9b2086d548f8a68e735eda1b6e7db8147b5797cab4eee84064cca767a27aa261cbada21d0ce544884cafb62818ddce1b7a0e301e966a9a33fdf5051ec7800ac6eb637eca331ee01b53cc85220246877782e13dd2caa9d477ceb4176bb5fd8e91d87ce2de8692424e08e9d8b44b49e1b6800ab19ed50158cd842b809e447bce6743bc07b446de10607bf091c3baa64684a56faff226d5155ba573064e4b2cf0fbccf408bba9d9c7c77d2bb27fdfea02b2ee2c15b729c2b47936e81b6606fedfefc769a052528577e3f29fef1aebe7edbc92b1a5f830324d229b8b7212d04d52869d611cebf642f09b197917683f9aa0c30235a492ef5579d55a86a7b5ff03747c68ca56d9a7c8ffb06ad44eaa0e3c347ae15cb712644701f7d5f34d6c1b73637bcf9e1be9f4bb40d0696fbc10590bbcbff44fa58d8e8896426ed35f1775f009e8d6dd3e6a059cee181e2a2e45ec589bcdb630e24f47ed0d8ccf49ace51e8bbd0884be1ca30dbe645375e177bd0067dd9e94739a9f70a8679945d4fb82fd2f33b3790a8fd4b6ea98985135b638eb46d493da5cc4b4ad1e1ecb2f9d1974ec7a071406a07716dfd83926dda6035f992bbc179df2d8e30a33e821e99ee9a71558468303b6723b9736726d4dd0e65efc62970bd33eff26c91c0e126bdbf20da33ce96c287e43799d1536c721b18555ea45f9e6be9a39d937a2c081d93a792d45bb622aa70b65c9ae298851299fa278d9b2630b986227f17f7be30e1280d36061a33f0c65d70008df04215c345c32bca62c6c25aa3027b3c25f03fd9e007d265135ff880a9f0b3aa07ae4bf87551c6a5b4cc64978fd9a502dc5b54f94ec423efb41ef1e4d23a07a7dccc853ca83525282e39f29ef5176cf08b1101515037092f3ce4f01235ecae271f07c3d26617ff4294b6499ff90ef5dbb4462f7c108d7110418183e1f88776ffa2c0610b237c8bd6ce519f6c4724e1171280f755d09d705fb90829a01fb1c0bef0ea5503c0f1b4596bea5383ad7c8bb4e84acdd196f93c036eb6cbb881dd98a75197d1514b7ad8298b2712c65bcd57c1fdeaebbe949d94193950b3f194aa74b5248858f73bb0435bca1118a895cbc0f9936f5e6de6a6db5d7a2a854b5fcffd354759c7844a57c346c75f856649d75be5a4adcf48ca7db790083e52142cf2f48c2aa1141a344dd5c377b88d3d1ca4231a2ad54757e5e93a8e079d62efa4af35159063579406eaaf9e6bfde9230dfdaaf130ec917ee1f7bebc0d6f2d71341fd7d62a57fd2714fecc7f844d3523efb641f4ad096239b76274244c1d55fa6788d9c56af4d5d3822ead59e9f678388dcc130a1bb9047f164d77a28ca114a82e74c121b4aa3001a4143fd6266e3365d7d76eb154a292d0fafe213ed126a19a312512130a4549e68dabc321cad597a170865d47fb06ba9ec5f6db32873cd2cb75223afdeb26f43dff45554781d1a5398bb70385f8afa1f25a03d24911099eaf1aa00ba673110f6091c7cea2f16e68a41591b7d36ccebcc4733ab785b6922b2b1d4ebfe9aa0ca1b8becdeb7d71d07700a932275b2a8685ca55d83f3ba1b2b77a86ff81cb99dd0167cab0b157da2fe0f80d2d170e60f347d3d4e7718ca38c8bcd7a4af054b6748096179148a132e20c32c39ed782da4f9ff98a7fa5b5159033423a7a55cf4f74e30485b3382f8b8cdb4b2fa36c31afbed665daf3fdded89f5cfbbd7784eb307933bd3852748c9d24245a7dc3ba28f8692bd9d7b9f5d9a8508e33ad42a3616c2e61be765d2f399da552f95a3742607d4dec1fed8d1c68706391106de66b80a8cff3f42bd7acac04a3d7d11a68c49d2a68ac671ee5dcd92a884861edda7397c44311189b1d9e3557a30b3497532d19630659f5212647c53737bfd18ba0d5979333805b32af64f845fb93c3068073fbe939582d8390e0629b60388ee23ebf2c3959ab2ade61a10c874e6d6065e0917cba02970637f93c777ec69598f809b8502abb9fdce8f6aab695e0a0b07fa204238f3fe4613b6a903f9ee624025c62834ba4aa10bf1f39cd7dd95a04266c75b85a5055e6aa98d6f23c4c58ed61e39c613d54fccc18fc094243b2995f439eefbda623b04f9aaa71d67dbb2703d07b04d8cf20666a0e3b06252dba7af8c4746bf0985f1ab0f5e14027fbcbe5c31143754ce1d571d2b49c69d173e70d73d9e04450b843a822149c76dc4b4678de042910eb32c62413a52afbeb420f32d2dc73791fc7050067f26f89892d7f7da0b72ff89ac68e4130779a64844f0d8565b0bae86c3645a8ea89dd785209df62e39f4dcc9df3aac7f944064f9a767145e8ec4ab2b174f52984a07e52e306c9d1e350fb38faf6ed2472160155c41e3ee46d4398ff59c613bb48534f81e5bbc72678431ff92b228db28604d7624fd910775becf6ad9ac698d91b2f6ce20452da430859ab58cf08614e3d4127cbd0fc50e3d2cde3bce9624cd6cc759946c07c6640cce33cf30add074d9b36bb2931c709833417fac07ab6395638608efc41ed5c58483d334d0f88a1aa2ee1bae6ee38f140bf4e9a93fc052a4c54b86f796b91db54d15e16ab898745b4cf567f8f88935fb649ecd6e34312311908d83d69e4674c92cbabb3249442751b8175b0341f49144e2977b6fbe9787c0555694339b6a4dcaeeea357b14a529f0753a7b3fe9ee11010c307901b166981c5fd525376f3e67fe1c1dcd9babf0b94f0649a86eae27d56698f8d2c63ba96185d45ee39c2d5d09bc527ec6ea05b11aa541508f6d73c0612efc06627b346743197ee76accddd16426cb2d220f5531b2bf9bda408887b4ba546c16607ba4d6db50bd946e7b35992c6cc87e53c8854cbc729561181f718aaa68acea9aa601a042243aeacb281c635d25aee9eea9c8ec88107a0732f80cec9b571500a73c9be95b755834663825e3f757562030df4581c18c444c4d355a0f617b43516ac6adca36c1ca68446d620a9b1b20b67e2ce6bfd0f200395fd6c7df9d0d967230a1d15c582ab6291e5dc9c0d58a87dd4d5fec6431bec11a0a9df38ba68fc22eb132ec881d350a47065df1f33e933d5e72c04f1a7c40d996afa24265dc3e1079a88bc21a946d915d842e999de6c31d7c66219cfe1a612ea727977efe39a639653e71a8d9408fc34951784ec09e4c5052867cf06126b49209202d01be246fb7f224920661c6c859ebba55db987f69caa99da4c5166c1af4d1a139f0bc870385aa9806af15f44bb7ab04b9d48d46a19b8200186a55a08134a9325435cbf57e64fb88bd0b6232b015d7bfee12e7702e95d251f2de2d7b725b8c17c7bf77803bce23cb57d0c1db516b6df219eb615cc8d44faa3d5753a6d969b703b037de8c41875bc42a5dac92d969d099ed5990ebf35271b73fef8103f87e6d398f1d5e684fd725f08290684536879f0c266c2fc869d3a55721b11332bfb12792f14d1486f6ecddef2b72a5471183363b4719bac82e7bd928e773f210b94b98618be6d5406c0db6c41ce87775774987ba236aece3fd8b744d74045c581502ae096cef5d3b3fdd0f8a0498785565700933d9b8a5f1ee45c3a39811855c004d4524378710fe5b456a472e06f2a6d8a6db98c91abc0daa4416669b925e719576189faf42ea3082244dd060c35c9144ecb9879d7306fb578ac426aa8f71b20e8828bfac6461b016e95bc178b68f9d5025b15e9c3c059701c3cd137bd278b2065834a01181ff9af690be68a7d361f994a31251d70c69c001dd8733b820f3bcf6488cf760230c6af8073c8d92e940a9b876b42c1fee16a1b1ef3a6ba48dc63d1c98e1dfda2c3564f770775ca8605b7e943b982b6e478c8531bdcf5d2dafc3c413f1a9248e47ea6d45b620983a0eef224b970853e18b0b6361a10ab9cdfe12b92363455589bb469e140ee36cb990b6a7391ed5324dcdd22cfc1530ca43fd9cbaefad878849ee800295a5eb15f71bc0ae9afc370cb4c46d23c0261297abffa5a6ebf9a16e82f213039cbacaf49674d6d4e0ed2e782f842c310881e5b46500c606b3e367f5922a87bce1b98f400c51727bd7103463edcdc36657e14509d0b8783216959e00c45eed8dd8f64e8ef6b09d9002bc12c9523549b2c86b29201c8cb7550a9d0459ae5210a8d80a6a8b9ff14247daf2edb89075a9107529e8f207b4b8cbbc95c650b8ac12b315a0d86a16e2c1823e4dd5ed739adcba8b84dbb6da57a83bb1b29eba2ba76dcd25aef979758d7fd03a11478263bc00e5ae11ce3187a8aa1885a7d893845dfa6d9bb8d9e3caeaf57dd0f7cf5620da05b2b1d926662690c65f0937f64fa0322a842054aca626f47acab1ccddaf9872f3078944aae024ca0a232bf268acdb7d8b3146c01e6192d5ea7bba4cbe51b283ba030ec46da0c312f8eb686fdf3d8033b2aea5ee81ebd67c2ab936682110a79c35d59cd04c486e179f33f2667fd7065e0ae99cebd513f161a06f844037a67e16fb467ceab17ddece33898f06d534d8c2e65fe0061fc68fddeb71fcf68f9e2d2b390a0dbea9ded6cbf3f377fa025156d9cc237daf776833d5373e559ff21c8b1f6513ae84444f7bf62b2194872ee057f0bc750f8f41c39bbaed59f9a1636a83959c615caf184d17d7b0a84cda2ccb0ad87082edbc08e6b80b7b4e74224a869d5ca5d5b9e3cd2a3014bbb5a191df1ed182c3742afac2a8d3da568919e778d83e973b054c3e60faf70e631d0e6e8b8cf7b5e3041d4f3e2d7633755bae34f6182378b5d3071998f80341c5b0766708ec9ad022eb555c06aeec694ee0798136982ee2f521217b6796a1013b738a9f34475d9c7841647adb0f7fdb7a2a03a3489048c71114a97ee495733358249059299f653bc9ade9ce71a7b976a06d818ea62eefa208181e43f4c7b21bf770f78e8eda69350ec446a959df932dd3c15d752cd944fb8915988f6dfa878991e7786f539f2906bd04360bda82e3582220c24d4c577f93d27191f2e9ba70c85e2855760c6f93a915e60e7d94401422d00ad06cfa155eee3d2b8f63d3402122a3918ac56564af9c5b9187e75da539aff6e7e49349ef2b843d170447d49cdbbfc13d0f18654c68526d6413ae6f2eb4d01717e14d73bc633bfebd27bfb4e6628a44bd6c72c062abbe05d13774b242d96ceb9dfe27fa83aefc3b18b295795d218f8e470714918b03720f10135f0f31ada304902755990cf75f78e026d45fdd3cfe946301e57c041bb132f4c98d22aa0ea750551a143fb271519a5f30d0d088be561531de2b7cf304d139c30d110b8cefeece0dd6e8aa2f69ac3c82898f91a2b137471ef192d5ca517dd6f8ccc9529a9f1ebfea969354f776f654c6ddb87256ab9eec2c8e1769fe13155c7a24e74b674d3fff52908fbac21726f15142ca6c52670e053de7879edb134106ff75994cd03a3fd7ce7e040d920588990f5309cb5c0c050d640eacad6a78a8c8d933abdeb758345f0cbfc5a11a1574a57a0fa6ab2955b5fc3ad86106afff093d4a2d4ee087b3c2643d71386d44d17ade0908f0fa0920ba739a27e754bf6a755563f01117e85f977e8f6f42bb48ce167125a146909982c44c5270cf86b89cafadd75cff4c5594b08ac29d0309bc5dd795fe78243db79746b875d5d004ed066afde5176b1db529693a858f12fc07d90a33afc1486a5c5feae53964f6994d0137d8cc7205cce34bcd88007360f12e0ef7cd9e584fe1f28473ae816f0367f2d75a1f66171f28b8123bc684bc412c6893aebce8500564e5c3b6f779782bcb998a948;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h348e1e24f44e21affd8603ae6626e1547d3b484257b516fc6acd8e4f8199fe9cb5a2d71ad0af2d56d7f4f27d7e1f03b5a6849ae96832906cea10e77b0fd4813cf301d0a37d6bdd06271eb3ab331bcb287fb562571672ab1263343f3efa794360dc067d1f6883afc1225f447ebda58da671b4ef58ff203e5f4a910652e06a669c37b97b02da7b1eff3e2a8e7c68f377b7ad1f814705346406b6caa04514c7420768cb0174963f10c12f404bc7648340196637dc9634ce6f0d6b0716450178550da64c67e05a86d06be28d7e9420b0d0c67a2870c3bad04ab8e83200bff4c7d7fba74130f5ac712edee05ec5a7c2f6fbd62549f20e21f7b5788274661b21d907afbecb745394978847098d65f1c0adf757221aea4c189268598dda98882c59c4226559a942b8b75c0840e1dae6a4e25ad592a87e004e839f477a7b62a309ae44941f2bf71e956aaf18a88cffcb092b8642ed1e9de482477df1fa58abbc7e6fb9b2f8acf49464a4d5a3346e034429867bd01428d04a4c97fdeee2ebfa9be3a6d9a6d0773d14f4f9322d3b0e2fa8b7dc306c0b90577140789f0d33b95463a2530feaf428ec7fb0d5e0f5e9bbfe96f82826cb8bfa594232c339e2482a1683e4458e8ae188cbb94ba22386bb7d0af5a385f65f1b5ea43cd85add1856c31152cf6f93563ebfea87bba1e6efaeb209fe3351adabdeddc02ed0583e10389e323a7d0baa3aa0e44600070137a22917ff758962a0794aee86f9fb61a6b7d631ada906c103490bd8706c147a473d698401d1760a92e29f36b924014be4d0ab813798c272f490cec9b83112f28f225175409c1d3f3971d6789ab257bbf2ccaf9130a95876229c819c3dce826088db2e5c8400ed3b6a481ec64ee7574f29c8a195cae4231648898ab65277f9d9251258a4fdb84d521ef18b62ff66840941b824f219fc3e15d7219b031e0a87e4006cba327ed5cb58a00d31327d2d11edec4b440a8b7c7615f6c6bccd2059b074464e17d1e2eae0af686118b829e3729d678c33b6922a147ced78131017f9de64d9e06a100b1a38a4f6c300b14577508cce2eb2069bb3bc42c38c3257b3dc2c13fb3ad1ba6e918b4f480cb63fc665368231272cbc566be9ab664d1ee3375e2b52da9228c96a887d48613ca78cf17a4abaa22dd817b051418631d0f0696f8e1b9d590ae0732e65eb4e479accda4bdc7449672904c88ff1a37e65493a3e273d22519dca94aa5f5d2c7ed99c786c4b1f97baf48c414ada83584c86f4891ffad2f3d1dc6b5001a8554d49ba07842799a8cdbcbafc22a4fc3d28624a801ecee5c7e7598bdfe903a04636686b95d3e2eed5bfff2a9d2dc97d964537812da81a3d1e812e0a0225f51d3ff8ff2d39403565ce01ae21478f7cb2dfcd2e98b8f711c1a055fb7d3dcc58e21ca1f6752ae32cb480c431cf70fc80b58bbb08c8fb15f3ede89ae33e6b638dc01d928004139bbd65c0403fc7c5fc4909e76ad984e00f01dee1c9a222d97b7f088946a3580da25c931c2223baa89ca6af818be59a5ad521efbaa287aedb02386d0b02507f4a8621276cb217d757d74a9a0e96d800e4776d005d88d4b894c1c9ffbcd83b596b94011e16696dfe3515570b2ada976da7f254e02bb83796c63b85dcaf5389eacea9aa96f2719a15d6e5532c5d73fe2714ad5cb2ff1e080f0fb35b54ecb7b76cff5864592694b99b41c57e1a6cf2133e9361f0c413d4c2002f4e205c0375b3bd903c27981200d855802ff6f559d30484d2503b4e8bb6805ffb4c98fc7a602590d54accd6e531ed75f6990ba00e7cf13c51ceecf9efa24b05b7d779f563b1d07da592d715a97692349914320b7d225e618e4889e1e0bc6f333afa57860dd1a45469df938d29d2adead3277f3811ca2e0f15a0dea074827e155839701fd2e2044c4a39a2b690897a351c8cea6b43ceca7eda21d0d7d29ad92ad82a807ee40bc64c70ce941cdb441b63f994c811743c84f65f7e1b844e7f60271604eb26ab02ef0b91dc32f1555716dfd405d9fb9ef51af3db99fa1ce680f201edab04e28515e9173c5ed39aac3646988d32e6ed15c52a54c6c727368b613fd1e64b27e1c884659fb6925283d5c220ffee2df9a5535cee694ac1602c6f5c45775663b0f1d98be4940ef56936762a230962cfd4490711d4d1f544c42f9e5ab8315c0358d4fb73f426b4bb21daf57d6bbe8e4c503402d13f27c00c1b1bffe22cd11330cfe8daed33a6875798b8e8660a42fe0dc1999019d55a4cda16ba7234b51113cb9f783800d4d453742b6937e4ebe0e1b2f89fdae7babf85f49739f3d20c0a87cd11b6284037095692152fe532c3ca567991f3d38cc6f957af74778073ee38da5f833bd8d0ae683d270438680d044e6ae24290ea9dc9ace953420a648365e4877dbfba5511f42503173cbebf5224c73116eed0fb3921072d2155974f1cceba2cea152e6b817d11e317e8a997e9c1a4f62041a60dc8383942cb9315bf26f2a0af8fc89bf18e972bd3e4ede643e4eb9a056aebc568645baa7c097b01dcc8522ae1bf797745525ebde6ae68912ffc378c0ab5aa9e5e37312f0255081726196d4983e7886ed760f76062e037b1a1837c2feeb7ccfd56c7450d16012db9d66efbf41a85e22d6a647f16a8e5f4c232fd5228abcd141177131a4cead6b05d6c39b1d6828ac19667c98b64c73ac19bb9096fd5ffdacb5430e0a933c58735be6e0d272ff627b058f4369eb9176ea1fb65ab4f0ce9cb0341315100c4b69fd009d89f1aa62adaacf5034f802785d1422295312b481ffebcde54d106e1fc5b1cb0cc10efd84f5e695242857af661141685baf8f12833ca47b45c5c59c0adeb14def36454fb0e9bfd02c0cdcb2e02bf6487404b80f8489066029a3a021806622a91bba9dc05829cfc366359479e97657d9bffae82b8528f8b7eeb8a3febb6f7ba14495d99166d45ee45676512b420d42bfd050ce1ea6ecb34b0f43893568eda7a8b6ebeaeba260cb9bed61af0c8e95ddc8a9f4bcb86426fa3c318adc890e5cb23c38673910423480f4762152068cbb2b8e9f7833b0547c9ab7510be0601b536fb89b06cc95f90389371a7d15c855c655cb777f4046b797729cd616c6de01731661485469ea32af583ac888caea101e79760c011e42e0245bf4247e9e73043da4e2388e03b3f180b900e653acd3c120ee1dd34941e062f82068a8a9569280b7ba00e8ef04affb6092287c4d3bd91c864ad1445a271a365f5376ae375403dd7f003ce018be0631d6b8637ab686da67d18faf841c7af8fa2fcb93eaad7b749fbff5547c149c899504714ee8dc4d57da7bc086c5eaa6edfaa9f9955762130f5e38a4f353d84fab650134c19d1aeaf8f6a53a87f0468019f2684dbaf6f82715ce8d7786c9560e074090ff4d0e6ed6d0a9e2d9e030c5952f9c7727b1038be627bc9815aa20826c188db9643b6a1342571a9750a8ec9670991cc41aa44b735bbf27781914b0b4b4a46ce8acfaea5d29073ec383ebc40f4df107a152f3da769fd3cdb8b3bf3f4505d262ec57b835e51e6ab51fb571d9e959c190cb17c5da7db5df7ac016cb569b0e228efe6de3e1b4eed1ef81efe26dd0b5b5fbaec891db56719060cc70745ffd3c621e32e632fd61eff622d1a3f2a48246d45e9ab2783a08b78c54ced60e28dd02d40a0a3dd7bada3200a51b1a21e7de6d7e36d026017fa124f10bf2ab296304995e58f9c2aeb779aaa1c87aeb2526be19740e9edd79aa66ff5be28e51365cec89206d8e58b8b40a72b09a91004de0b5c1ff8fb79f2bd51fed4756e3d51a589b591372fd4758ae3b46e202d41f30a7b4c0822b444cf38a9ee27f49ba6848488648f930da447b3b87293069905e8f98d217f3dc505d8ca4bd27d36058634f8f8f0ffa168977d70b4d1ae44bb558ec8da5c4782760588066d9208a79dfd3b3c693ae3b5c938266534d64dde7b2f5d41d45920a60ca5eb2881657c910f89e5a259f7b767d0bc7111d606709cfc208b05fbd3a26898a6c929ca5b771208b82b842051302969d6e3a3c320bc2e660c1c51b8a765f75007ccb0961ab50c0e371199c9307a4eb2b882e375091390ce06a1ca98dbb417b5630fc50fbde9bc11aa344f97069bd7347ce7a53426fea7fbfdcfd451039628f8d7688b62834d3e7209a4e0d77995732748ae1fb6a868950f239baa2476cfe7b8f457dd87ede8263b0574553d4479fad6bc0cdfe3e22446c68c99caba003a5aa8eb1d7615244733a5ecc96044a1f6f73f8c2df80bc436df324dc5259f5a50f6eef2f0f3d5df1e2e7ff9891b955b9da33ee3e02de1eec92c7868f91d3f2ba9f2c94fa59761819701af26fa0b81b68e5afe14a8d59ee30620e9dab032957c61801fa57e41a5bb9f225b84bd8cf163c09a1984fe86d7419498dacca1e5d2b03a36fb14beaffedd06b1e6ebfe5edf20e93ea3a7012cb5fd6f12b847d62273b7818750e94c8b480cc5c8b2038461457c07cb5861ecb30df2f63e8c15b7ec71649c36b4bb69f5e2cf6f8dc33243395f58374994a8c1c66c3b37ff00b0fcaa44ea605b8c70972ea12ceb1e6453ac244b2058bd747f558f7c4b90f68d751222f750b4c2180493206caf1d367932bd9c00c528ce637d9bbbadb95c1f348a22d56fc95a79f0d2d55f0ee3d5e0d65b1991b9e1a95cefd67349c060b020c7dc3671be77bbc36b2d7bd9726e44f7c1cd9b54e7140c0cee835fd6fed211125ae30781128e10bca5edc9c1d928d5eaae0c8dd67c7738844dc60999333c55a9c94674374e20318cc56d27f330edf238b4a5cbd4b4d18d1bd48e56f657bd149388b04c2b6f60af263225ab6ca220ed97ec9e3c714482ceda4ff484996645c255366af87b539865541839ad440ea8e3537570b7bca09e757af4faa66c409ee437e64e2068d10d231906bc7d5244fbd52a77c15f80c34624b6d54d8e3dc9605fb75f29a692d7e67b65b6c1c5ffb25779ee047f4c96fc45b12c652944ee548a003f21454a630c1d1ff0f430572e7ba663bb91bb94520dc39d74f278111439ebc2d49c2e03ebc5616d0af0f2f33d4a07d9307f46b65da6834b3e54683a183b6f2f627565a5a5b26faac3647721958012e99445f74c61a31c134c5afaf84f7291c58c42de643627b1cf86742888c41fc57ee12e452a8e9ce5f5619778b5f9e652cedef167a2cac6e2c21235c3969c0be643fb9af4a25dbee7297312b97e609b746a2330954839ed2a2cae65c8ff2660675e07221bcf241d7559102020fb93354801a00b5ccfa6c3548e59f61431bde8b0f723a313f00bebbad7ea1f10ec5ae54c40c64615cbfd74083c0e4155de462a42395e236baf9d60d93f5ac50dbd7b9bf982d953b9ef4f2b7dd6fd9e9cecc44b7d8577a2b5f4a7f4474234849b5a680751ec6507dde2212c7847c833fec2c60f424587d45b910bf32d19af19b611508568983b67e5e017b17f9d515dc3762287d78da2f2d21f55152e0bcdf821dbf2ba5dd71294ab3fd1338d5188801cf6fc4643219687ef56e4a45e95fc1515e2ba24e5b586f38b80a478c2ab7aacfa4b6f2b0434e719dbff99775487fd597fc20cddcf34e1a39ab6f25bb11e0342ff5527da7aa35aae09dd85789bfa69b0dc5ea4fb5597128ed28ed26b396f9263214f38873a9bc451eedac3eeb675e1438278e6ae69793eb79da39400c3c7dec32a4dd5e201eb6c7785cdb08116d37d600e7f2d2519243001fcdcf2d317fd8af88b39047d0ac28cd229f6ee52c62102c037cfe4bd34c5b0e4dec602afb9224568f91238a42c1e37b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbc35614e359b4494a390740e49f78324a5fcc15eee849dca8a6d6356357eaac46009be412f24c77b43c79480e6194f8ac9acf0f90882239b65f6418c659adf59cee1aa8ee0c2a4a0e02652963b8d456becb851f34fde10fa9f14ac0b9b9a24f97455cf990891645797f3ffbb5209ccbec3e84ebb06dc16df21a6a5991d711d50662d4269f7de2c26eac29d248408d66ac9b1c475a0a5885cbfe6537ef2b869a582c3edf59bf7e8cf47a08046e2bbe989fe449bbaa271f3e33913e77a633cb72ca37ce9645f14171efe70efca785b2e40d250b9f5aa59f54dcd2babea9023f9ea4ae14654007b9438f260128372345a0aac9abaf30973fe7a5929ecd56c0aa22b2a56739a84464c47466be8a55316a68cce01feab884dccfce30ede7ef81e36640ce3c5050d4a5183310d51bb5b6a2e34db9e9c5ca07eb7e4b52621c5736cb8a1fd6aa4919e88020d596e714ebebd98c184f22d820e611d2bcfa1e5d85160008c17a6107a754d27f9872e42fbfc5652e37a14cedeec73c7d4d2fb402fa44186f3cace3b07203c1845d2a43a7ffd72e0f73c9c272f1f51302046bd4a249bd54cab2798c530a8739c3c5f807fe5b3f2a8416c9ff7729f46cff912ee11aacecff478d5bf8c5eda040119fa13ea3d34ddc8b5d3dc1de87fca5e52ef5b57aa61b9f40bb8044b44d122cb3de18daf4108e05b4ed7fec598d6a8847e6a39de5185844ccdfa6f952c673a4a849107893b82235989f6657634250db785ac540876aabd077f7e8e5f7ec4d76bb0fd56c3b88e034f2ab65a11febba07c413f054ff6fbb67a50b696aaf8199564ab52ba5fb3983daae72023d3ec6aa2e712cb886d09eee24fa9a43f2d0e2baed661a60233bf80b9c83697b716b704e3ae9aac657291b4ee124dedaf291fe9d29ace832c107d3124b1cc516c71f211cd47f191935e154b8657bc1c89ca435e466cc0bc2ebb9f8f88bf95c6e0f6af72e4c2f71e46f885fdcfd25d3b413e776961902a900cdb6a2e57f47c7d003eeea5f238352550b9d9ac4dbb9f3e4323069612678512fcd9756ab13f73da23694e1cd9eb339d1f89c3f1fcbb073214c9e6aec9da0ef9298c0a8afdd6c35f4b486cdfa7bbf2db5e0cead24d269bec1b07b6abb1407e5d4668b48e181a3551173d8d62d841c8bd39fc1da174291b2e090a958bb188223e85dcdf466724012da5b907eb0ae6673b885216aa39ba959a4e7cd661c29d73fc74365798d16cd637e1cfa07957e9c6ba2b70bf11eb6c15faca50f34e576482538761aeee34935b8f7f38eb7932ad8d84d2e9f1e36eb84613dade859be9bcfa45a68c3cf2badd33175499763fa3c23c69664d1aa60ac520af257667054778a793c07e2f0a916321d5df4a64e795c35063e0aba806ca58c0b5bcfdffe4b8f6a6f5eacb6c741699271c95b77ae12ce3d23c3399fb28a448fd9305690ebf91c7d1e7189ac36454c23159bf4fc270674e9447398afb6cb72de5feeea91730bf03deda66e59536e25ec035e45f4116c6869de607c97459764fcbef5f8208a699ce572c6ff7785fc0e70fccb9868bc75a70f81e35fbb7c7b968e411f688c0873e9b77286e3cae9de264b33ec79c0b8d27c180e097ec3f5ff631c21254aa3987ef9c25b6c34a6b9d819549a08022f7a15def47e99c5a7f739b3e07e75a4e389acda2e33636f5d98623ddb161b651db51c771fea8500d3c57621bb27ef166ad6e865ff21ba316e32caec62be78adff171b42a158bb64f31dc5801d5fdcf071b08fcf030687854f4ea2b475aa45f78c4ff6e750b1b9e45d6e381d533e67eda2029ba227f926ce37f77842f67946d6ab23f14312aa47aa40b87c160200ac2fb99c49f44540097e918ce9dcdaf857bc18c6a012ad056d7e7b03059a70b4c358b0fe369918994e9d99add55a527a32ccd386e6cf788c9b6494c43dffbb6dc522f972b918d44b155eb3379f975afce40da87db29998a85bb36b0f48888d4a3a9b15184a89b3c7ed15f2a532c80019ac4bde6ac467a8c7f5823cf94d92c805f935dcc70c1cb53cf39601153a4eef875cacc27ba0a8b23039a76c9de1cf225ceca431d3ee5a504fe5c8a25250d6e6adb498ccbcc1fc27f27e2bf4a7a56439e424fc68ec0c9f2942989f96051e70996f2964b297667e132d5571de0ff76db4658b04e917ec25df0078b248fae3d4a2aaf86bda4f493c9bf0a36f8a99f450efb11cdc05bfef1133e1690641c1d44503ca2d96b5ddace6280b7f1ef10363178e9d1bd388e4eff744c3e232f0b53815d6b3c74e3dd00238dccf7b30633eae6e034aeacd3a658d7cff1582863f4336924e42146aae4e960ca1c86b4414e8e2ce151a892800cd13c0e99f6e43945899662917e3789ae18c2cdd73fbb671c028375b826254d08ac5bc8fc5ae9297741a6694a66746425ffa27425d9c38450e0377c3dcbd0e3767298908dc01d904634e4981d68dc777fc80195021d9bc338c00f368b4a37cbcc47ba2c6ed5dfdcd9ae70c7bbdaad1169ddb6e7cc93792d2a8af03bb25271f08965bc83cad2a1a6a9e16dbb594654c749e332fb0135282218b0929542603c3a18556e2ae3418b0ce9b57af34971936f38337e0ae14dba0f8d55ad6951ec042c56d3da37ca744227699d952ff23e321a977c097472942c32c841538434a30fa644c26ebdd54c3fb260596ecaa2345d8db56b1690c3ea06740f7a10131a6c22b377c2d4183df38fd73f9a869e6f3d8eb84b2fa5e69e7bbff63fe587d1ded46e72c5e7a46c40e0efdf7f51b00126bcc98cf0cdecf8365df0f42ffee771bbc8e4934b9fed54fd2fe5fc974cf2c07be14b59c1938e318bff9052d730efafca58bca8710ab3d30f818fdad5d14daa2d1fa0995b383e88b093aa19bb35f42b485d1ba8edfe5b64949621079c8832b63d3d28ae2cb9a0c1603792835dd1cf563769f13a2e99bafaec018a6df6dcd0f90172eb9e683fa4abaca567ba41ced9a50571995b0df766b8b90bbc24fa3ddd98cb611613c47d72b12d5aac63db555962f1e327879d53751a25586f54c25e2114540604b323fe4b17444e7d0428fd4aa0b5fd973ddc4780b07347da04ff17c70e43f70ce865c0c4236a7cf05c8236db7d6ffdcc2d179d119d3353717810dc91293b4c12c43fd106cbbc630b483254a1b7fd0d1e68c0e6bece4fd09d50f7b7c0b21a281cd25f2ce5eccc8155371e9bdfc9556fb7567a2dd3236ba492d78eddf666f77b496ebc189c923545d32b05b4a80ccc2042d821b30258bbd539927b084e6ed60206c297eeb19172fe451ef03ba10a578a27e848937bfa2d5613deb77e15652a802180a1d106a48a7c00af79e6fac66500fa83f904d5ef94aa68d30b3a58e18303fe1ebdd3c89009add285c31b00c82c1ea28e32bdbc225729c26d7303590e21e0f25c151e8d4f0bf13f1173354e74dfe99567023841b9c1325572b751f196fa74bea497b57ad1e31a1b0fecd240873b6bf8ca6190c9173c578274182fd6bc5c4894684bafd99f29bc5a1d4bad409469286d0e05780808c6e9461169615871af6a33992ebb22b341168eba3f6fcb2ddc083033af78bfcf76d8b7dc2157df1a84945d2f2e2b90cbea32a1d5683fb4ae98ec3e9c9b37de64b0cb007863cd5a7f08e44987a9d80efc0e04096091508c137f9611a15d2b07b06efbfee86966db120e9f97d23999aaec61016ffbc8eee1f83471399724e0a34b9be9ca3b49ce7a80ae2dd95cd7a677dee3b6dcc1aa378b8898c08a61257f29dbddcc4aa2b67a9ddcdd569b137498791393c5a61669cf4811db19711621e81960f664d5e9ed73495f85cb4cf61f315650e4ba792b305ec09afebb20b9f01e3e2fb99e7c78b63154ea9240503f00d9af1a7b4b323ebac7ad8526c778ffdcbd219b05057217ed3c5f1a832f18db56509ddbee4fa3400729071d5a226add543c768c729995b87b3faa745bf3751b091a29afa6a62bb06834f58839b249136b21384315bc052865e70fd7ab48f6040ac000c3ff4fd9fe99395f7ec26c98345514f0b67d48360c0260b588af442bbff7a17172cea6a87a25c5b675097693a271abdcf30463e96414bd31476ea4488e3a48dbd4d57d47fa162683d50fab0675a41e6505201f32523dbfc4e9e094c8efe7f929044fefb2a6bbde66a21fa39f6731d0678cdf66c624e42aaeb7049aa237eec5b93e57482ac70cc249de282f25261ec46a235fd7196385c868a8b98e1bfb4be26def9bd46b3eec277e8ea413710de64e82ea7d71be8e5fa24154b5a84729cd2c5fe3173a151a880e29be93ab7bedff1ca4fdb18e0574988904784763a65e64c6ef6eafd0dc3e3a04f0d246967bc7b166fb8c74e72774ef38c60b7dd99f21bbc3fca0f746f6ef09be199549bd037bcdefef66d3a5f6e2b5c017de87401d65395e02e891b6448226bf73faec9342322e82b701765e47dac010c49eb66bacdc2d6fb5a699342f465390c718a8a9e7821e4cb4d2706c28bd3cf376492a76daf0fbbfe17db70fb6d2a4c54b88194ceb0fcc1755aa1db668f464f43f68c83c6afe0032157485ecad834e580cb753023e12f43ea5bd27fda5ee8333a04dc3a3b96ea782115a20ee96df3f7ec3071f8c16f73b7d83ac3d1b97b578f615a95b3eec671dfe6ebca733ac1661dd4bcce6079005b0d3071703a1352c6b8e7800ef1eaa8d41a24aee622296aab8ebfac20a227a6681db70a6a548db333b0a3389c1a52ec202f8448cf94d9bb21f5f1b1902dbc851e2540bcdd41eb5f092e6d6be8b0b0ea7cf706b05bb390cf38c570e6f5692a92cbd1fea8b6cd86db913d15e416165f88b4055c1020bfd7a766147047909d22edda13288b267c3ccd39d2ef8b01ebf2afadfaaf279c3bd4bd9651da81499ffe5ec30656c5184231ca6cae8fb1fd898e59f4ef8813b0f4e577aaf976cd4882b27dd8e876baa6878da40fcde186e9645c977adafd2cf19317b564e62541005df0173e93b8b83946451edefe3a42b5f1894ff83022305b0caed192211588208735bf73171d4ed7685cbea24001c0273952a3bf6fae029cc88e8e4588e766eada60424d739ca347796f9d6a7c4b84d0725a9870b01032161eae6a6539bf440fa7e86dc3699cf4ce6630d1ce40e8d633c9b899db4bf264aea7534be9aa46045220431e3ee12e2258c09f5884eea9b9b121c2f8b0e1180844709110e3c68ab321d1dfdebe945e038dba67c565c275b36dc266bcfc012b66b2ed8129dfaa606bec8722651ac51c9128678d27dc794b7b6c4207b32c73a018b5a34b39c0bb50b893915dbcebe8fa9b481095e3599997f8a374a990867df0f5087142e4d2daccf72290e7ca863b42cdc662073b1fef5bf509c22bd39aa48a01eec2f18497f267696e296904aa67236f10db1558924e8815e3ddc5bb02ae1a131b149f6a7751ae2e168c8e3383da86fae235099a7d514d1a385ca87f12856c4894cf0e71ffc61636059f2cb192ec26585e300a360fa5941f6b20b956e144c259650594713454942e1bf373cfdcfacf1bfbc408e33e7b3c3fb2059281be13229235e25158dce7c091e1f18ea232fb13fba677704e190410ac75e5c215ad7f6d186a8914eefb49488c3c4eacd284d0d138bc5d1e13dc53181f799555806136d74855a1754794479334519c88d74bcbf67f28ddae5670c09537dc67f8994fb688e27792f7c64be4cea7fde6622756b38f36d1d6b05e3cd9c51e55a3d55244e3546d697f17b1ce9ed21bed83bc24ba908054b4eceefaac84b1539e014ca0c680c1ce0446f667ee2c4b2e31c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h679c2bf8b6a19d42a587125331106135b7912e038dd438f4bcb37eb3dfaac6c1659a2eb571d1b8d472220fb491238451479892027292264c768cf1b48f9aa6934da3b26d99cd78b5cbd0aafd55bde6f7fcd285598291aa913aa727cb5ea9cabf549c204f816541db6f466e36099779206a831cfbb24f1b95ed5aa8231fdfcf6157582f91b69afdc53d389b0508f93c7a4a7f761c4b1df3e5862ead4ae4268eff934c205f7a2b95542cd04139f770f81a88e93e7b30eb101810b78b6a8b737179218fad4ec487bde213f52160edd4ad5772d7fa019f9ff9246d1bf67d74de6750b4946937099926310188636168921ffc51f5260a692808b99067ffe6b5c3328ee885dfdd820de2f6e5bd777739505ae8aaa5b5289e87a2b82e2c08cb17b352344148d1adb175f84b01c8ba9a7d927b68281df17a78a4c69f36a4699b1a507a804d7a66a097c4528e016825b7a051594a6d1ba8ccf8260f7661ef03e46d778514d97376126b6952ec5d7fb6ffc99ec0158b7b8270d15e372e642e2988921627337d040fb497ca2a14b4ecbf67cd5913ae3ab82e544671dc38724fb981dccd1fe23ae19f4b028215b68f8ce6ea10b77e7371d73473b4c49c5f904f31bd6167a66991170b50864f0d9c64a51765231947a84157a2abbb64358b27b540bd16b61cdfde1b15efa99a2971d2c2677c6fc3f3abd81c5f06be88a84cf4ef594b15548c3e6cbb1c0e7f3bf1a4067c9159d0b8e805c9a83d29a00d7f4871539c1ce69d57fe2d6606fc82ad56e2d838246aae6089fa6e39fe2bc8c44165527ffb5beeddf84249f98a9070f071b617ccd57517172878a49a3cacf2bd5e7de683b86bca78a341d6eda238cf885329466c9b9de28e5689446d87295a5c655198da1c2808e61cf38bda6e2865874eb5811cb660d442e25f58d8b010e35a7f9b86fa8d191f66d9980d757526015d41187d414d897ddddcc7bbe771f790d271777ccde42f63319f2b6dc8da39ca50bad8d13c1c43691027e5decc41d9a6b76c4586546559577b6e0aa7634cecd293c33d6dea00a0a4889a58cd100427b6e7d5602e66d41957a452db24b75e4f802b71795e1eaee87472b9b03a12cd765a2ea06ab9e12c4fbc6f3b14f765e387150791b027842beb13bcc21202c8375c29d1ceb35f4508aa07a600a9800a0d83c720fcdf38c036f3a11861713e886f5153c7954868469cdfa0d5992df6a29c1714851b91d4710597ddac71ec4227b1b2dc9b01ce8bd1615c607009a20d692dc5e9253a747862b6b6580151a340a3722fc24d05235cf4c204811159872663b3879812aa1afa68880b67c6cf19646fbb7a913d6af9547e40cbec409ce4909780f8369f1654ccd4eb8fc5b432590aac2b482ebdd483751b8bec09ba390ffadf4b4c0451f2521f7e5288fe6e192b209cecfb064ba1b902502db2404b19a638d87f232fada8b6a2bd97baef46ac543faf7f039b3d243a3fb96944e34f46bea4b723ebfcc58095a6ccfb7af55c6defbd4d9a4e2067dc36f160831f128e42f0fd14bdf2ee74b1ffb3dd06ad42c8aa0c5d68d012b9169b2aa8afd0493605c3a29f0a1ede4a4a433587cb5cb30ce2799cda2ba9229e2f4e02bb711cb13c0a4a228762fb01338c220b8a2d463e1bf51ff2f355d6b6c28ac0e74139534ea3957f05298db8dd86e4b9853f2b246415c229e5b776ad4e1244982b9815ff24885b1a34e3cc0c44aed804b5586b8e8251e950e2701d6c092d42941748cfa1eac8a13031feec8e5879648141fb3e183ea311d711e8589119efc71cc5a644b7bd2a0fd72cbfd4f6e40596243c83d5b65e85feb9ef7e78b520045783aef6bd6d7558d5a66fcb1147aa5f0c17a4ce8abc4753d8422a3cd0b24f3db954006578c01272905c43fcd3b89a328a1120131f609d3c3341f5fef11c06b327112ec0312876c4f4951895382648d97da8cf48bd62f6896c2e18e435dcdf836c426afc127b2a918fb54b6b1edde099524b5c884e3cd075a7b14fef31a0c22d83c630d41aa4d04979aa321d0afe906b4b72518d8a360acbc804e385faa32b3961401b18c1f7efca4344ffb8b76f2b6ed02167c18a9e0abd35b3c832c0eb79ea9298fdc8e7726ec14f6cd7a02244850cd94fcc249dcd18014e2d0c3335683f051cc34e05ec8948418f0b998aa2da6303241a18160d734c0c24e613158d5dd1003d6f71c2a07129032988ddbd01a4dc81fc190aad31f5ce33a41c5be6c4e1f4cded7c615aa8116412fb5d223826307806737fe250385a7ff31ab2d838f5613f77588eab7c77a7103ef6131a3e4473df772352e619e03f994635c858a7c0226b59dc8028b4ecf1e2d178f3b56e2742bab4e7e020bb155885ec2ab59c247c70fb7f0d8a3a6b18ef2a7476329c009b409fe967d478fc46dc146ff1adcb2586994f5bde0ba5ac6866ce566fc83b0163f5fded69e306b51a7ffd26faf1a0632fd57a08061f3366b56eff35c7a2d26f9c8240d0e8871cc61fd8662da7688f3c5ed7ae4ed4b82b8830e82e86ed9f9fbae700c15e353ad986595a685b2d4db80c08640dc04b071ddf7a20e15d00f20798b09cc1120028a5a19fa12c22c640ee26fe655cb9e14ed7b5a0f66b686f19e380121f9241e20b706945bf350c4d89c775958a3566c96e86fb5caea705655f261e0124a1c2a85559d7e4dc442926c0a2125bb5b55fe718a5a7e57af8c55ea4e59d0813b0309c0eebad115ffdc3d2a29366152bf8faf0c3f959d31658b83f4cb86ba886f06b9cf95d46f2cd12d55ce6706fc1f4b103a1eff8ee05f06a92399ef4567a9c8c72c52895ca7c35e6d5ad53270f9414d19a62b857fd7e215da4389bd0d77adec2af0045fc5efa1f9fed0e805c00485d9b7dacc8453a0a813f1c5dc5aa2d907088cf7f56084be4cd201d5955851609954bb5324015173959a0875ac0ec575e84294ef8774d45b2ed37530b91e98802960e3db8978e83fe4820c2022ad963582aa6b6f955498267221423cb36b562ce80af6d043738d875c144bc035f18987ec1683503ba9e7c8470322bc66448c1ddd7052ea721e90c0ad89b023a10cfd30b975f549afd075d18df0276a203c667f9f4096dbe5469d8f4b9d1d7a2720614f474d19294a576390273d7e69445f8521ba7d12d4831495e1f920bc15cdec04b6685a4959bafff6651740ab9fe73373a3e6a0ec9dca33ad020804059d046daa29e55e8d94b50918ff2b6db1f84f97fea25cfa129d2fd139964a7f0199edb98a3048e505e8879f9ed05e94c3978e28d298a76c690df1a947b9fa8f32eb8ec9ec3c3d5af442f328acc200a2a8846e67d2677e24ae231bd8d4cba06613714ed4e6523c4ec54166b40b49e28335e48665843978385b41c4dce4f0122663def31f7af9650efaf4014cbeed3c7b10e104e3a003bd682a0e90ea77cbea2bb472a9ead43fc967f352bc08eeaba897c443c5e0936a8e4a65b178e08bc2048956d7c91cfecfd8dfabc57b7b13ac3e2e207dcd425b72f19258bf196a1653b447a8aa512c2fc89f3f82a75f68a691241c7fb20ea0139e6b4d7d660ec08023956e9615761a2af1f04569c341619b5538f4fffd46754bfcfa29951031b0915e196745f9fe204f7c111a92fe947a36cdd80c1c26a5991ab507c5bef0acc99234a3945a50fb561c1e9604727e40972e1087705724a684cdbe8295d10652f5a4162fcdf1b0b9f469c720e1932019b7d919e7f3a252ed61631d2582e2c668cd3cc2e42f47cd3e44fbd3a11c821de75201a37911d2e9cad83226b24b01442ae5ae0a2b057d44819b533f7f379ad629baf0725fadb24064b2fa576de719b2ca461eacb756c81daef9b103c6be277f7e17b367253f62dbf55d273dba6a21dc61d4c0e855d24fb07b4a64582534c9d60e1f1a12ddc20dc462541dd5518896d3a3624ecb1d2d304d8d270b765e6c0aa3e34aa1010b4cc2513547b7275459f503833ed4fa83160a3f34b230e36fc6f2f7bd40bfcafb9a45220073ce5d9a04e3b66674571ffd50fe32f5c7c47cf6e8125c2f7caf869df341a4c7d914b19ce16b8cdbc945a1fa53c17c2972973fa6ddcf1f47e32481db3501b2ce498c7af8afeb333972689fb5c97b8b90bf190099dd816addae44dad474fafc9f8a2e5bdf7fcc4716ad65b08ab843683456bdb4f7baa9cea6bed5c44a9b8937b31faec5f38ac8d854c60b2f8d4e8ac945df01c1ce81ffd17c72dc8179bef666c235b2f07a040d2265e79c83db5de1bac31f49297cd7e2fe822d625dceb8ddb19f319db1011e5119f9ef12d8e4c01b53cea271397f45c94743ed2fedea14cb90ca0455063412e8f7e79e25f16d57e2ee58bfde3448c44c5a5ecc4dada07e36353e3db6df4dc4292710f7f009e4be7fa2b93b3bcb29e5ee16e23450c3d56bce5ddeae7696185c392122e1a72812e38c7cda27bcfb52cb3750855e356689115d0e1bac83b23c66a590befe640cb31a7dc4ab30151da4ff0fa39251b6256897a3dd9f341789afa42789c15f0aab64892d9307967e361bc441c7980fcef9798bdc498ad3dcd94e229025b964154a62043d2ae4ffb7666848e40f90a3483d9bf22e0fd512fd218fe412669563a69500a31e8dc1acc600c5a2d0e40c8bc8cc4c1b1f53f16a92853bea4286bc0363029e81e7b234488cbc8604ceedc1d0795c2f931a131b651e8f1596a81686e07d0a6e85ede2b87b4a41c8acae58f60135e19e9de9d9be9c6664f503d27748a0d51bfbf8e539749d6909842276e9bbc8ca1fd10b47c1ebab894a8840a41f0350543c5e762f0575cde666ce57e4f606e89754d4778b0136284dcd4939c2d6282f2b5c627f39c7b839ef32584b2b509bbbfaf465b86b0ed7688979984b54bc7345a670a8c6375ababea81c31ab71e01d21d6fc17df9ecba4c16b1263ec19e2c7b2a48b16f15bac74091c6733745ddfc08e82245b1e0faaab6760d5f73e50645d7d7a61c5a9dd577813829866bb335cad953f21459c45caee89553e142268ff85acd67c91ff5d6f0846dba7f8dc779d55f55e8c6bc05bf99b1babfa22c9267d9ec30b2fa846b537ec53ade303c3346db699c9315d5bd83613a660fa92f1f934556ec555ef8c10b3ce65b190e341fb696f1e9bd395cfdfecf778a1aeec371bf063ab577b6320c10de7d301058ba473732f6147d0c74002135a4ecae46d3e79d83781446f17dcacb5f2f6f945d2c609d090b5f0bd5a3729bb7d9f88353b7c1105cf6a88fc67daf434ef5b2cd87c6de5f9c7c368d7e66ce1f8976ddda08f6e2944eae1d4030c018154fe1e7e51ca312244142e05df974f561bb24f275113d161104615bd25317515dd001182e7653d2495b888d8a4c746bf726d47a59f523523b6846dbc267e2823398ad012d1f5d2736ff9cc28ccfd5128d146c1caf69207ddaf1a30546ddd1d7d859615b409a61a1cd714af3c787f5027f858adac26e19cb86ab86cba92e4a4fc7b6314f02dc6f468432f7636d5bea03844d9bdb40c5b8f021d4ad1ebb236a91e64bfd699becada33ae54d6aab854f179528e7b79b6efdc57ed9a818a8bd6232f3159e2b9ece1289a60c83c32d3d74e088b23d9083f007217912f8e2290417361882af397a8a1dd74b5ecd868f68b90e47df62fc717c1eeadcd1e2bf712e3f5a3f86fe87866004e64d9b74a3689813a3619fdecc8518a1546fbf801255f00e3f01d526ef5702c8699ff49aea652c7c56e9b1bc286ef8f0db0698717e19876cf8e7e0cfe5632c18fde22eb635efdf416976ede7660ed9c4365017bab7b54cb2ec646174e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hece91f9d1f8179ffb640bea9ebff0cc18fbc52532a9b2cec7b82ed568e3999a35d9c39dcb75bf3502db734aab33e3c8945c3b5e13140c7e60a65b2b71f9f65962d2f2f1856f0f7a313cd9a04ff98649e8ef2203febba73c08aaef84bb6d13d6974a3a4fefb337b96d0fd9877bb4ab9d0fd61e649cfd6782e2bd9086e500ed601f06615de16686a7796c0ff7644a5137098399767fdbf7c689747b9bd94edd7f3795375b7832559826647b44bb2ad748ec1ebbb2fc77e326492a074f698c3181168d9403fbb40758a2a24166564a340b51b5c23792728ad62c00da94eecf64fe5fe30fb018f1a9a0e2afc1d59a6b17b440ab65e2d91ce11c878b3a220344e757ab1e2da179c9eb4261f68c48564ef316df63a257eb135e167e5ab1b0acb1911725899de909e44248801cddf39dd91efba1e52e4e1e6b663a7c11b0ccf634cae31177efb0f970777b3627d90fbacf081860c2a4ff9151a9007f0f1e44053c02c57059b81cee53eae545eb5661626ffe14cfc156769353bd2505392f665b881a7822f98066fa8110219a183fccfdf4fed565b685f7295e2bf9717e570a09f41e7102ea1808ddd9e49e33cc13e226d8d31bb4a25c58f7f92e2e9dad611b23b1d24980301dee25217838852ccc9a8199b77fb2129b77d3e09023c8a61fbeacfa5e5eff3202be171b97e0e43cb2db673b5913994ee5bf43aea7da4958874dc354a26e0f843bb2dbf75ece197b8ab4e4769375107ac1be5ebd7f8bafb2e5c9b55ea96eceff285853c0d8b57ec7c62b73fa2e6715f4c07b105f49fb051dfad547806150952bb625bb44fa6365cd0ca711495b9353f3a2e41b5e532fb3ee751b588b39588f85ee85cd4258d949870924b4ac7139cad3efe1f4df89b114fac3e1421f43eb01ace02f0b31818d898b45a0d670555c1f6129001a6cd6bedf996bbe1da992c2355ef87ec08e4147808777bb1653ea42a194bfb0bbabd66e98a2da148a898d2ed2be711f3f30b54c34387775ed8c04caa13fd481eddd49f52227af6c094caa2c3874068f6ffe4418b7bfb7ebff9769e004f7998a35b96479d7bf4dbbd655988f850586ec380eba48206056e71628c3d0926d39ce97f396cca532eecf9e40d814a82d196a5c6238409395c2e12836e5e198f86d4345f9e3a4f94ad0918abb5a4ae81b4bab5f14016cb5a207d539db377dd9672341db162f391a05ac8300915be60efa90f51cbf31b019621a52024313153af027e76cc2cf8221928e344bae283bf38f793fbfa4e3e58488264ae28c444bf6afcc8501302b004ed9327ee8d40812617e15bca15820579b3500a1be5e2c03e7f7c45911b914b35c94c1ba8196d9fd041f376f80c1392d4f4f61b44f1fcd3a2b14cffdcc1d606624649511a9ebc3bf682683887edc8ee081bd44764ef838a7796ed1ca50049fb9e9144db96eabfd235f90d3881ff69e9cfbeaa5bd93666b60775236958a07d16eecf84497fc8fed564124f9abb3d123317cfd1cd1fd7da24516944d2926aaba33afe310adcab14d2406f667cb3cdb00236d249fdbbef787acd6b934f4539efd935928fe21174983cf45eb1649aa51aeda90f3d9109dc7f1cd8c8fb88ac1383f59b64814fdf25a0b91e6f925fbaa625620d2bf0dcb63d765aba2a47c1fc9fa1ef5a6142bfa153d6ad65ae45871d685f90758954ce1dd7ab1ea98b25eecba7e321cbacd01178d7045887879262d15b96c418239c692624fc1388281048f9b982d26393b6abfe91038022d37f25f9b88e7f01abd18cc359ca5294d887a0c905aa4c779bf572bac483ed99fe6a19894d52cd6331af4aa4a4b9a9370f6b8f1795a4e89e39505dc7bb73b437a5d8a2ead1579167cab584870b6a4d14d39651441453a1497adf32544c5647295fa0fc5e471d0d221650ffba3ece197554d8485c87f45d92747783e354c461ae654554585a4397076064fe7e396c610957d7cff58fcf878fa19fe3c8979b788f0ae7ce84b4d1e1dca8b145505bdfefae9695748a219aa31c1d4fa6f04d7e3ee333517f945c5cfb3aed94f5833b64047c6d70a4b6a6d0f16dcaf2e9d57c5f086ffe518f5cae52fbded68fc6fbd9a18c180ebaefe29ee68e5b63bdf7fa933965a00774a7184ded1d17ce3248f3fc1ae5d14d7be60cba30f697aaa84ffb3bdec91d46f93385095d2369a5322b0fce3828ddb336542666594b8d7c8280f2aee2ce8bde7c3152edbda5f451c086959e6702528a1fdc0777ff1483b5ba3da5aa4d92e3a2d330c7f0dbb864a49c605b242b2bd1a98e4b3e88dd99d698df812b6bb00827578ad6ef02e0e6562ce8ee4c129b762f053816104fe17e4e29daf3cbe59d977abc2906d4e113144a0b14643d1b915af46b0cab572b0e5cf9a95275b6067034376606e78d9e11a87812f4aa0b64646ce0c43bef9c40e5a9fba2e673bcd45ed8ec3bf4fee8c9054200d39990497e0e8c5872ec1c48f72b986f7c57dcfac90e7008410fd6314d8441fa90259620b27b31ae8380c9964d010325ca2e5cd8c0048807653ee47083e88e8797ebd7c007cc2100aa2c60bb777eb0b136c6ad1bdf42069e8d84a6f356d378b797a616820f523d1c4b7232ccbef3150ab1d9868aa2e5e81cd22acc0cb46012da8f74bfc0e60eec5a4af174fbf11cf21745346c065d895c5d78887f317e9956f79ef23daae139f1cb4e46ce0a21908863dd7d834b1c069f1d99c29e9a41a9011ab42cd6f7de6082429fac113ff329000a919c58c31a969527bfb78087987558f23a8a72a1d6ef8997c21efbde37cada9396d34a4f8cbf9c7e1193541ba7bdfadd466631bd69719099c7546eeed8793523d1195f74c3b0659410b1d6c3d9107b095e805c9da6f24d7a11d39c10b99d0537859464b4c72046b968b28ee1c2787fd1f35ba202fcd8fe39932926718c57f47862c1c9f6d59762447cd43d5b065f6781a667f8c7268db02972ba585cb9166a6f12b05eb9b0a8b6accf10fe6ede7e8197cf05d05de4845bc0104caa1f5438050b77eb99775bc5d2720e6bd1c04ec5ab20e4879a140154468b7604ee6df6c6b37460c05ae51f58f096d1b943c3fe1882770a26ff7207ccf0567c3dc12c1049e45c64407a8b543ca2e6e1c01d44154d83c32b18cc70a4d7aec28bd8a773ae493ff1d690c440d5efe9e40b2a9a0458012c5501c23c28900decc16602a5d1533e89dce796aa496912ee78630a581f1685c0d4a1862d20b30f9cbb0f9acac7f63fea7e64b8650b85fccadea42cda8137d50adbe30c4085c7cf18dfb1bf18cfb2bf65b997da1286f4332b0cd6be7aa6a94a76797a54a39242016d560272974f1f8edaa07f5a445f0089b8de78a90aaba4a3358ebd5dab3e1962d49c2199f73a3b300ef6d5eb91e349ff8f00d86852e13841aec2276f1c3fc842cf0f7ed3af52b8e94e472c3a32f8463ac1ff00f8403334c9cd80eed659e45a1f7fbdd84d9f0cecf2cde34683979c94e3cf419fabfe69d49120944d1342ac8fe21284c100a3d1a892fff368c9f94bcb412c912b9fa38648cb47db66a8fcc252001a07ec88b3534fefdfa58685fae4cc75e5e7f5e09ffbdb89a3dde058726c28910982674171b4c1928919d53dd64cff4e415d3b18fde6c1e0e22a2ee2ccd9fbc6dbc40036116b8f31c5eb4506fbd952c0c532692fc1d07d8b13f9fcecaf3018426e87223e0bbd3bb9aef401ad9d08d49dc89579bd3307a3cd539d88e090b61d6ffa2caa8c586f18f29e517d59c7826272ac9525ffe2ee8cc24125d12b7c3220795c2c7a33e53db410ef8d0f3de55e335c20e3876c472d61852d253d34f900f9c04e8821393d721acf7c65c7ade756e452ce120d3b3ce9d5a08241cfe6a8569dac6f154a5890ddc9b2366fde6cab4f5d45d841f81985cd260e77d8a1dd14396fe939bb75827cad129b56236d641fb29472f0e54cbe758b1862327888061636f97b913891d6ad8a9e2f8b63d2c05a64a41461596857539941bf78b25024765b1514a674e8bab27292060f2e07c0cfc3bae9eca773e06c9f6e48c0de2671c0f4dda96f41e94f41c86851b26bd062205051f0fcce8e26d9bb7b027470443d112332e5693f1141b6a55eab5c7cd6d232e143fa91ba62808f6b88efc3244799c502a45e7670f3be2a18c743c786af4b7a309acf577bed4d4c9d02e651c3ba2f134d00705c5f111ab6a91e73b445acc5c961cf915b80f44a4e4002e2695aed692f3e6888ff6e38edd37d761216baf95b1e587fabe4310203b7a62f7e9a6b1215225446d2ccd0e654b39820da8edf52b8fecfdfe2e5d2d0c4f9cc71d9ef949067d26b443c053b1649bb0a34115544e063983932f194b612f540fdb36d8507963761157951dd041176d641f454fd54036ea1ffe837d8a7b376fcc2e85fc91d45f6a1857cde80c2917320f482911b35de11b70a915f6964a098c04d17878184495d67f3d40575fff353c5607cd8b28931441f82057937e680f0d3adadd779c66a23eb552a234ac94c1c02ec53780afc2d1c383a05cf40c216164fbc03ffe2c2dade6c29488084f59565ba1e3583ef9251a6d2671f585b097fd4e5ad4db27b03f3ff0cad731b55151dbb37b035a19575600ac7bd9c262b02481133ceae8ff124ad9097f403c2d00f1b8077626e443e8c77784ba18a902e6763253efc4f16405940b6182222597558dc0db57904b1a85ab22491d03201fe95a58376a3de5dd1ea5487699de3b6557958541e6365f6269514281193145a5d811a798c092e2a0003eb81fd6abc6944fbe1e525c7585273f2859a261c0bc3c91b8f1acdb12ff95cbfb2c6b3ea4d8df52122d95b09e67cd38de14183eb53082f36d55cfcc4e6699b7b50df6a5087ad7fbc4136ca712e809ed2c4d3cb0b12a0d880b6d4b2094579680c1834d2b3a89babc74c5fde0c5d2c5d78cfe197f41fff3c4e6f7b080fb92c5c7440dd7b22151226d2bb54ca980b6dec340574459159500b7766ccfaa33733cc3844afa55f91ea1a4dac5b13a14636e8eef4a55399098725fb69849de734ffb738bd6a8b631b7718eaf99f8638162fab4f4692e2f58e32b040f79b63379231a0a49122d10ad13d0feed4681fd935160229738ea23da392f7045518a7d19a23c7a4954788ef9396bf30b6e337c798a2a548c3d0cf3166a6a11829d6238a812be217924c6fc2c34e235827306767c25eb3cb851c3adb8ad60a3854df1817ed406a87b8f3fd02285e279eda2fa4b9651941cef459fa23a0fbd804291082a69978055734350b7949f16480a27aad2c4a779c0b2e39b5337f5e48a6f42bb296d2fbf4c81b65daac60d273e5f706f820830e223d31780c5b8cec5d444f9e034ec7ce1ee2c336165b05293411617b8ad88e4a6906f55e5c6cca73a2d81b0b17bf0fb2edec2c9f5df21acd4ecfaa5440b3324df0ecb1489c1b3add5bcd0f0ff22a462466729bfb462a74507eab32dac753d27a880933ba35d3fa2135eb670759be7c94ee88e6cd8fcfbd010e900d273db68241b89227238b04dae56d9b90b19c3dbb76080953244288a2316e400baf390d1123775855db0f000751edebcf855d0e74b41b671c708dc5f1f4205119ebc6cad4de923b7895a986675ad54fbbe0625547eaf62d2e5c5f45fa386fe8c532516d96999abab7a60efdcd225efc9fb0b3eb71134b53e8a15debd674dcdb62933a889c350fcb8bbb52985b0c0140c6b1806f69b96b56ededeaa5390edaf535f982cffe65495d7dfe4e5b9f7f1a2f7b976d63d1e2881c00ec5c4ca45da91458daac9e7853d5c280928214b215927e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6344ce95df30bd35935c18137591d592764a0af21be363f7d5d92f2ed529b36e68b15053bb295e1b13ecb5f2c0c5aafaf7c091918cf41f312b460b07979cf9f21f1bfd1e57f3074f53afbcec4d4339a65fcf147afedfe945dccb590b2974bcb15312536f667683460932d176c42615c4fc1a42e1ee5631aae5d0ac440d7b4701921f613844379d811faacca9992d8b50cdfd0b5be0b6767ca265fb5024d1b850ee53c85a2f6158c61de5dfce80a01427513c2fa050b44e46c463bdd39fe6fbc589e8e112621f8b5c56eb266ba62beeae48019a317d52e0ce0e8b2f8a851f31e6283be68cd71cd576032f589c927ac76afa90cab79ddc4faac8ccbd2f2ee2e535ec4a227f152c17f14e930a18ca131f5afb689c2b2221e5c42e9644697bc95f6967b1426e7a8257e7f314bf51bdf613248733839ffdb643eb0aee229f4bd2726058dd14ecace11260c87bb960c64059f88eba792bcf5eca45243a7b6f5b4da1aa1749aaf04eed717f0057ec0f51b1dbf588e7f273e088d5c67a44a5530fdb69629cd600a321d3a52ac02c15fa31f79291aff478131f1ff1f3ab52e4f742195bf29bd5589641e858488c86976ffba2797e74c269a67046fa82a83f353bf057c08c35a11b7e187e8337e35b5975b0cd770e3de932127bc9b4b7b9c459b7e058576b3a2636bc8d4aa9efebd0ca9c86f30f97070b9eafa115bba0ef75c72052e912bef968ec3b20b3edce339d3173eee8c495af67a028f55926a8855d2aa83732c844c78f5311b124c8b5bca9c4e16dc4e98ec3b117958ceffac2ed51c5ab921c84bcaf7db179dbe704727200544f74e3e42ddde0437872dd0ea6b7c8ac2dd0a44d3b97bcc6f4353b665cf830dee9129b5280237f5ccd4736bfac6aaf372e0dbe02635c77237b484b0d837b876cf7f42860fcc6b94a210d4036c1f7e5ae38ca488186a9917e87e541e7814b4d81278cb8b783abe45399bb38ed835845e89fe2beeefb1d16b82b091e43b79a7dd2f5edda21258f40aeb448ae9fbbeabf450d9abae13fded031c64c4554a92bc8a5161a7268b0342aefa25084832550d503b355c4f56e5ea72ca6443730fc34e63a71e931bd55fce795f08c33d4ff37d940668eb29d48786df22e7f63334d2f6627e4bb9182ccac95bbb81c718194b1df4206fe5001dfdfa0bcc6efda36db6ea717d892332184a55876224ce458f72603e74705cf324346823d2504515bfd5b35acc535e9afaffd6d170ad89a053d5860cddae889d4d96a606ff80ce2471a243318db4fd7b163ffca05475a729618a51c17f9bd8f8a9bce4e432df9baf7281848e98a49c1181a04a6a0435e0e1eeb5bc11cdcfd720da1758dcc91f836f3f73786386803aaaa9263387822a452c4eb80c819e9cb3088f6552952f347aeb31b141a94cd139315d911e26739f98373ede9990a3c147c2b6c35e2409b63e94b5c92dbbed94707eb57d3487b33c2d69b58268cd140f9d1d9b9a5b8d7d34e28893da46cd1c6daaa4df057447ab5af85e780b441e886afb62a44ea7d1ad8013a2961befc80659f361c870cd76888d41c7e329b7791363da03f9eb1853291346cb83f0510739f3d018724847df01aecbdc50d3b721f7297ea607a7828e53db706245cdc3bd755d5d29fcbad8ad946c2f788744d93a2043f431f9adc763ca5e76b58bc2d321f2ec86af125dfbfb2fee5b2b1dde31e22626cc2bdfdc8fd9d7668f99e561074b84932446a6faca23b62e15963ffaa74b62fae508f71a801422d1d71dacaa666035e6883e2a8dc81536bf531a95ffa116dca2148183cacb7776e91eed9137a9b775082d1da89549e75b175f20b927510493a853a64ed1b538fc3aba2668987ac18c92161a7caa91a254ecafd965417435f13f771a4ef6bae5f0c3b5e1c30e7041b5e4d538a8de277dbfe6ac0182cba0d3361bcd8bb556c5990dc03d5cd12bcb2dabf1ba2a3f90e9e3e3247fcfa889564950666de4116cb03ee4924c75867ae3df80e3dd1e1911f7af9a6008110dda311bc9ae89eb69eceb1c371671875bafa42c130d72e4e1fc7e4dfdb5872687902d5485c36971f09b723cbed1348b1d79462731e099957389e5f52e077aa59bc7cbe53dd34d21af09cf0c63cdbb950c9f7b1c03ad5ab48bd0d53500a73fed2e1bd958e1d28aac9f6a60110ac90008aa48596185056158d66cc09e08b7ba83f21acb51cc494d53f46bfbb2de61b4b5b3c2851e302f090549e756e236be6026d8109b8bb050b93c90876bf5226fc626750405be2718271d12b0c24377e1a6cdd3b50110551d1e196002e110cbdddfee254653904d15e0f24a3d42a4cb2657e3fc376bf0e8cbda27d201e6620b34858c0233020cc29376fb4dbd85ab813a9bd843c82e3ba9edc79b56eef59590f15ba1a3029f3bc3befbf2230876a533e74e9aca8d27861505cd816790aa6122403698b904cf3ddf07bf1dab9c41f3985d406344202358e1da559a5fc7e66fe233498181ae6dc7f4e6586d0c8d65af36423097cce531b602cb6ca1f78c7435d639a4a8f4c8885232753c6d32809947dccf77cb163d0e99194d99344de042acc4b12c7a49b0de70fef90bbc766f444fa47563b699c1180b9cae0205bb2528c409a181689422688bc0187160fbe2e1d7400068d4a250d98e747ae87e505abf530f1d190927a28eba06a9c273b45534ac23c8433b8c782f4bdfaf755f62cd911e148a897512bdb20e79574e54aefc3248bbca10ce15b49abe79bda82d0b4aeff19da6eb92de191dc3ebfe126a6894bab7620826a9bb3e17bc60cbfc734012eaafca25cd385b1193db09401f8648f124656f7eb3501a81080fe652e9bd729879276d000f6852798c0a157fe32fcd12e7335d091a7e18065bbce929f20ee31f0d8f4f19c07cf718d49a75afb11fd052dcacebfde46ef5cfc8a43d575ffd95a82bdd70ee2704755302fa952a7b12ad668874f19c6ae4c66d3f3ca1bfcdad200157bb04a7de7c6ae4747111ac16376ccc1de4fea7cd59645c9a76a7a1d1bb18df2a3232a0567e1384d5bab05c989d3a0fe52c978c40fc0ac23fdcdb447f447949479201c601a9c7b18339747db8be5e2e6bb061cb0e878f03c1a78f7e7d7d4d359195d5df9b0be6dc640cd37efc99d55c03c07eeb57f44381cb1c7bf1d6b8348ea35fc105a5abf4aee303eb22046c208a5256b237457ad8d2f1637e44a2589f044b9692f9e5cc447d92bc396fe0eff0458f6b103e551953abe63863b860e55650edbb73d82cdc61e2ff9f97be54e130fdc09922be9738ad80c42b4c32d36d2c9b0b3c7c21e8d870e7b99a8803d5a569349857e0c55b9df696375dc5c77ce8ba3433afcc7a46a8898eb837d56834e9fda1944af6eb080ad4c4151bfe468c390ecf7376938675f58b933c3824f08247a8721683ffdf065a5fc7b02180e5a938453b4a289df7a62ae82c8e2a4b10710b25ab5c07bcd104760ad2573081cd8b37d640783830c60ac9b3a1ec06d9427af662ecdd1310849b2a486bba66dac83101be1799936fea28e73309ed4e0b74af7ef8d94795c6fc0d98c8b55fe7e07a03039a7c9c1aa06c575a09f036c2106438ad6c994d9044b2a0ed9c8aefe0315ca855073b1281375a0453873eadab5ecb9aa0d9eaa84a0a59df494fc177ae81159f34ac294f02f9a5fe51997e7e803d4a48c1e8af9606961667506b129f2e58e7c3eabcf633377167771159304cd7151da76835cfc96d5ee50239fe780f68ace2ea38a8042d771d39786decc52d88d1668662c956aeec6e36987b1a993562119bc389ed86854eb4bf4ce2c7a4d06b9dfd74664cd3526c68e46744896a6309778c1b578b25f05a7ba3536d3b46988c7c5c91742e23410a342f7e65269a3a4e7450a43b7b536d4359ad67986747abcfe411ae958cc3b2c50b1fb90c9b0967ef76d48cc79db603dd2226f3bcf97fff88a061da8945670be93a2c3e05373651960c6bed6467e26b4498969708be12d4338655fa18ba9da612e67fc86705d24baeb41ae394dc901b565e1bad734b4422019355cb8d4750e3a2052bc1e08d24bd276308e85b37683c37360bcf5b110e93a5ef80bf384f473c92226824405879feff244c35e81265009c36537816e382ca18310a864b3c1975670afa8a3019d1856db0af6c80abeb65f4912f3d841099e4af1ade46a839e84de69a82324be194e3cafc1d95d2c9eb9360b0e8161eef49c8c08592cf34ca456d380fe9238374acf7d99d57ce185a2016bce7d0c77d35df4e57949044d24113223794fcadb9da3047b3e5d9f103709aa9ee51b31ad8db6e0115e28dea80d000f47c7fb128b0ac4daa2004005d166054bdf069d2d8c0bd00e0d0bccb8f34a26030c147331db3b070b88a8795d67e240cc1b688d9c6601efe1c0ef5e41f1f561bfe7c863b28f8be1e64b937298717e16268d89123592f35f59733af0c01368eff61e4b34388739fef287e937cffa92cdad58e887d70bcb28ef81c17f3774835758acacb00e8eefbd216cf3bc9ff1805d317587c16effedb97f940be9b08d09896c44445049c82df2c3498ece953f7e7923ea74fa1d860e82233079d2e371b99d84fb6b621f6adcaf44f66b4132f8e0b37bbfb186c469982c2099eacae96731b9759f1db214986abac0a7617c7e687d5d07212fb82f851bbf2f46798f3cc9fe17506bb9102a977b52d5b5d763aedf3d72dba775a459543e31c8e6de1a70aa020463c25f0b912ecbae75debf64c031d2d5d82af6aef27da016be985b4aa5c00746681d6e443478f1a7e2f19ec7ef4604b09bf539f87455cc42902412f80a7c19003893b7bd92e38990c7af0937c14e86ac3b4f61e0c44eff9541b7bfedadfa1dcded2733794bc290b434483a3cf28fca307f0ce1ab9c1b330b52ec5188b2e05bba89b9be09168218b8fda8753f806b85629415b42a051211c5a0c54a4424f483df5fa523eb0a5cc4be8583f5bdf929d8b2e979b87919cb308f7e8ee2ec1dc246890fe8db7859a400a323ef7370cd900a1f5c5871ffa2fb3c45febb3dbe287273b5d315c88588557ca1773101a9195c3dba5e142817bbae5f86f2f335a27348232455c8ac7026f21d5ed0d2290506b793f795843823374951b6cf2c147a6f11b12f85994ebf3c85269d564b1e82d040b7fcbf3a847df698de8acaf9d6af4fe99d6a06ccf7e252a8c3eb69d880c29f3bd758a24579bfd661aed5c25a93a78e8f337fd4d10cec9f56b022f16d72d6b126c5e0cbefb411ca6678d1426e04c0e2d774b74c3e30d86090b282b8f7c6426c9f63786a9f5540f98fe032ad1a13c0aa986c63b0b6fc9d66c10457b3278f8387affcec08123e22819e629e38dfdd2e0170c82f66b5b0d54adb41c910221592a5e7a50a2fbb1ffd96d1272d1f445852c64a5eb562f2aed160cd658c47bcc367fa6cb8742d6aa3c1de2590062b54dab74fdaf9c2e9f9b5d6dcd5f951e358c029c7850de931ba805d8e0ae9f9a573e12bf6453f6449e13612f5b3019b198811b86188c7db2ed07b59e22c7f81d734b5208ae095c1bd3029f84eae49cc3eb02193e8fb700e3a0dfc33c5e71a2497a4e950f766bf3d063a2ec4a53673880732b17973c686280d120130f2dff863ceaf2cf6fc93ebf395b82728f23ddca45abddf595af7afa1a4b20a2ce0f920ca8a592eb705eac83baca3f4e999ec663e3a0475aa2e31ac693dca05d21c9dd6a7550f0584bd423c4090b5c163e15ba927c06f60a692c0b6abf0c57287147921743f92231aaacfd20b289eea94b00111f068738a5242da2f56;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6395a503e7b895b888b695e10bb117714ce2e47a26da99b843fe89a2e861194594bdecc5d36882947d6a2753fbed24a4375a1bd913e383054e03c454024a36562a8d9c91c0c1f6d88b133c97d100a420f7bb42e05089afff967a2e4d48c6dd45d6377147bd430caa2dd8274638e63ed33ca187207808874acd45ce004d21419538def7b674a622332bd95e0c5074a786a3aeb0b45fbf02565851c0f425136c58d740cea30ec93b86c06c49bb0907d9a519f1cc1412e4867ff7b5468622d99c8756ec06f3f2350326b64b8aafb143da2889b21e69423e16ffda75aa7175a37e7b9707032919601bcd0acbbc5d106118f3247acd305c9a3b4defe9ef314acd8391c75a519ff4a89e91a2a338a06c8d883735646c5a91f44f9b064017b107404dacc56d1e4688b9a2367ab036a0be1ce1f5c8e27a431af009071304e24c4b73fcb6445e2d6e717500dc65e5393f54f5804452ba2b42f9a6eeeb5b2cd3ae91d2be5fc705ea6ad41361023a6ca43853ed39e4094ea1cb7b85c38102890f62d895dd3617421c1cd1545fc259a6ca1e283eb6c2724bb771f83bfae6c7784de76299e10b5f37d99b4128a6857213fbce8e7ab9bdd98a4db97b0f6a5bc737ae447b2b15b9f2ef646b0a9b43e3610941436f64c0d61f48a7bfa04648ab7c1d1b5b48ef242d5ac770efde8890d863886f7f5b09de1c138a82b39685ab9967a16a95b3bf8e44eae750e5771646ce2a2fa0c2b336783381e5bef40e375295ee921f7b0a0d5c148648ec0b40e531795f46809950be0dd7510080905eae4abf084cf93993feef12b631940072d7e5145275590a891bd8aadfe69cb2657f95b4650f51c69e1ba382c6b773ca0fca95e12e0f5e7ef7816047c747c9c4c1fa609b2eeb150c9f421398600b55acd13e2cc48f5d7192aaf1597c52958def24596cde38fed2535dee57b7a4496ee92ae49ccfc6bcb92ac499b6326e7207f7e03531cf22fd47551e20ddcfc1af8cd5a0de51b599dcd71b48944d610780194d8e9e9032497f58400703e6456e025a7338973fe4df9f04ed4760d031c7847b9494f3512a8394aee41cecdfe458d832a53d38142843b2a75a64c52ec7702d6fc1dd8475b03cf0896d6a45275e81c199f0bf738b99200cec0a0ffa13b320ef54622dbcfc1c33c0f0b5ca90bc749af18efbb61f50338cd504bdac574a16cdd0a205d8d33b8befe17b6d139e61b20d911856f74baa6cc59970d5d004133ce6e4ee1058a0edd574a66e6347e182047bcdd27f46430d9868546145f8b132d534d0a5a8f76d363863b3b7a6de050c89412b558b288cc85b31482a32d072706e9d0a9a2a164001050e7b5c73e3d89a8b984221d26dff008580249df2f77c73a1154f512e3941fed6c090b5269c54b5487cebaf27223822686d581b71ede525861b5a9d3e36d267682d35a0d45b2f9ac4c1216c010a2687f9de42a0579da48e8e53db6cdd68e02430f88c6ee99860594276880bcd3444aa85b89e80eaf0c48dcc4de20b5c7bcf201a940caf76023a155b5f274b70ef8621dd954ac2d4776b0456623b49767ce05808d3b9e6ac1b8c78018a61e5d30a7c3e538ac9f2c2f12b8249014964d213d08da1a7ddb6f641d6b6a7326285ab3b6ef6e7d7667bfe37b52924af029ec3082de6af911f719057cba1f62948ea2219354b6786d4dfbc20ab431b8a3480ad4a7d23804e020734a5ab64929d9be303831ca4bf3735f53dc3001a48baf36a7a06ad105392da50b8eebfbaca84c6e6cdcd6a1d81b73ffadb5df8b3031433730f31f59405d1e41c046adb9b8e4c80601ff35a89e118ce37cf1843d6f187961f7bd1c8080a194f742e4b939ffcd26e0d35b923569d4bbe67107deabfb1d99656489d81aca0c6e4f6b9b6e80b32ae1680a49900110f2eca727cd3ce45148fe48c7ef03d1520768ce03d07369cf6d502ca7389aaf8b23c66e71f79d614556e0291902beb220bca194d65a237ab9930db1ee00bd69dbc051a5f31a324dc91207f29cd361380f185f3377bffea15b8af5178b82e7a5a5374c1f74efab85687dff71b2386545ea4f501983188e6926e211c0e46074b464dd6638a0808ab94b4ed7b9ebc3c5b960f7499c3ba55862ed3a15f5988fc2a698e919a4f115aefddda7cb0a5b1ecbb559c6cd714f05256b4f77c713b0305976d04177758bf526ea55c0ae2c5a14262a6425c7044a10d682ad0673e4a389c715575898d9a714a95d272e42f26ea51c08545550aec155f1a69b09c95ca6d649b18dcae30932c7483222f5d856efbc8b6bc085ba912384af59b0c8ed1a0fd7b786f336cbc318c52eb156d7561dd85d212be18125c330449f8262ec9d82da82325940367804074b19652818410d1ad61d007e26d8c6a761fde15697a19b88e49c3181753572e03d278fd07008be7f3db63698f8b8ed4ef653af3fb6922861273b33dbcc4a84c5c81530131fad6575a6e719a638a9493b7eb5b9b1d19058f4439347e5b929bdefdbbfec356d4546294509b969c7599c50239310a5fe70509aa989a1fdc1670892126bc11442ad94881c806fb38c92a0fe7f4787d5c9acb3304a8e6b818f67fc131ea517986573de6371c13fd9db03185c72f62e4706e3f531c77768de43efaf104d1a451969a4227973388937cd2986e63cadb37d5e8a46448b49651dddcd52d0c8b04c0170828afea5f3c9b64a604c05d5ccd399f6975c107503136285f6e3ac28d66ca0a5556a0c641359a60b15a883943fab5bb3eb75d461d7b279dc19ba9996ed92619d4a59f6c01f236b8ebd83f17d407748053b5da334a50ef1b92cfd0b274b0b7b41b8feff3cb6b3d32dd2a573a1e778b5329c6f94f3b2fa5cb85c58356ffdccb956abdd3758f95cc70b56d9b5e2214f667c7850e9e1faccbf504e6b2ba9647566c512df87d65983c254520012468c1fce0e72db8a3f3ec130224f8b39e90fe2e0b4a33f86bd6b590111326c4c609956e25c6ff930c818960538cdde9f12d6f54b132240ca2f4a67f8a4d1bc09e38db5b93dfaba5db8332d0eafd572f0e7c6df7c5926c7b41b4aee75b575c0cffc876d9d3a64df0cd879042998ca4af30889e209f3057fcf7a068d496065e30d2078c6aeed8d6b5bd0fe7bd4d8ad0370dad80f7f5adc53003f7dcd1d250dededae1388dd713b0a7a79cddd2dc4729f9295b2af6feb100d580866672cc0700abee2b34dd18c8a640e999b5ac3bd2680a8aaac314c48c9dc22de0a7638e6f332b7cc81ad20422b65a08ddff93fe412c254382d511c94f5384603ac27bbabb0db3cf2f8abfde5b56ffdd7ceb27221ea0c0dd0fae6633a791f6a2f2159e8ca108b78d5fc890a511c57c9ac8eb94d58ae9f491c5ac097320b2eff3b49b480ab158c5ce84d88b8d608e8afb711205e5f35a7afc7715cb02a4acf7f9268a92dbca5f23e59527f72fbb96aba035e52733662ca2d3e74fd443ede87734e670c0e7d77248f57345ba4dc7b81ff1165263fb7455fabf66133021f6ad1d3b667f6c91688181c0cb50a878c7daf262a30dfb1c4740546d856290dfffdebc7aaa343d46798aad186a8799103b315912209b8a0d2ecd5145ba3334e955cdae8cc4a38374cd439eaf84afd932bd3a7877c011bcae10812f76378e6756bec4f8312a839a58221c26b323340da7f8115c20de5c524ffd75fa3aa06dc00619606e49d926678aac8dbb17f3e6fe3529d95607e8e77e4f3951197713794b55bccb998def5aa9bf32dbca958ee15f368f9110563669299a818692c208b8e7c665ea3d97527366a07784c90e08f9b424e10d547754fb5c244c2902ec89fec4b1d4d66fd1812340082d778e9bdd976db3efa25843e81ceff208808c66af93750f7dc90d43a9a800054ec32cba8c6d4908e7abcf892b8228abf0b3f2aa3b7e44c2389ce818ccd36d3175d9881d4fb4f334207674ec93bfe65b916f53d7d2443c16c2997d1a0867d5610f86b454b8287269eece483d1dfede03e8fd0b504b1405c4eb7d0db1c5f35c81af100a3b4f8c3e4fe0079e188d2b7e6ea404414400bd86fd04e18607f7553b3b1e8eba6edb786e1675ab5d6bdfc41ffc85406f23725a2a606e8da32f37598f9cd2be1d18ccb59485e49c15f0b2b91ca9484d68c7011269e29faba11976faed21987efae4ae17a9f86a3e661817e1ac36bb7472ff898a0ace7a1128961a7b3b965447b931e2eff9d5666e294faddefdaff889e9d98caee8201f50b79af37cb72594d4671f04745e87b189e3423e10797de016c4f762525919c46b2660ba41b526e161388a91d5df94d32eb576762e57eb509764b6366a479483b4074627eb4111de65457050f53b8bee8e4025a90709dc7397479786ba1a4fbe75e57463dea57451125a30bfb33fe00929b2455c21c904a9feec3a54e056d6a17c3babc3fde542b054d4c017c477b1ec4875a43c22be250419dbefe2db9936f8838a4d024cbe8a5ca93c965116510e9115246bf6b8bece7f2743dda2cb169b382b4d9f0ed88f174175d501c42e64fbf1fa24cfdedb63b6543830a3af4072fbf715e76e14dbe340d7698d17fa829ee82d6692f3438e925d3f439924c4eb0f63d52a2adad31b394399a08c6ca9f90e83f5bfa170c80221d210a389fd5ed6851d6864e9394e6139f4121bf026f6de44859da030c14ea13f14e41d3485f4d3b86d63d067277fd457cc4703540d101734c0cbffa2db0818de7a1e0736a31f68dcaee600e966910846441aa651a65225e2bf0ae13947e8c935a112c323026bf5070817ae6355b02809eb7c018391ea82127d061965ebb8bec0eef2560e3d6e3f1033ab88c7c9ecf7c9793b54408ad5226bee0602e280cfc89092c72fd33834c06831f25fc509910f6b6a0782fbef5f706aa6fe01106929f8afb47cb56ec982d1fb9b039a5d3bb99444032653795c5ba79bedd7673954ac36d906c5c21f259a1b0c8fcb3dd3c370d536ce2ab15a80aea55b9d8de5422d44f4c0e99103d4431e59d74a8e1899401c526e0610e48be1d5c2a27144165ba72245b10208017238a81ab84c810773ae61d20d80c47c4125a0cb65f1f36ff283ba3d94d20119682cc968d92535800cee6a4eaa96a1b0b3f51461a9d853e5ecd512ab79f2019e126bfc4e0ac49e2602ce8a7c1fa1701384343a353111c69c13b3eddc8dbfdade7e7c1fe390cc96df453c71c8c2af29c5d4ab79fae9e5aaf52c273da5ea106d4537aca217d4c46949950aa475e204ffb70b10d8c0693d0bb7d9ca7b72dae8a1e0e94af7759f0814814b33812e63891cdf1f4bf760419c48bc712d328135fa4d1adb7e09f413f4a695eafa2e0ffe9085ddf9a79739a652099ed8cd5b19fca7db0b558a33f2b4daeabed65c89d9f2e41d171707b0275dfe8689a6ff0f8bead77bbd8bb085493a3a90dc7e210c8c0df58f49540488a82581778b8b7d50e65a0f31b691ec7e65deaf65b8c5b0a75a0ec7e553d40217f62760d05c91b3029425f4d4bad00e4112d6e129caae5b1e68b04d771f69ff29d58432aa8642da13abc803bf72ad746b46b81e1fc55518bd9ae8d9a7734033366db361b7ba586a6e6a78744eb07d730bc35ce2ef78eeeb32da910b2966be20bd88ca50eed33bb5b3ed218347d0ed7934deca85986a7098c838666737270dea8c0a1621184f44bf7ff896f1dcb3108b7990b492acf98fd031292fc65fea1b8e3fe39767b440c6cf25b7d8de6bc40a3ed6aef7a1bf655f53c585eb57f1c8e3a090dfe1804b93ad055bbd94d79faa22843367cf431c13e0d42772d4cc2f1a37d18374d243;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h2aeca720462ffc8f0ef8f4ec4f703cec17a4341dac0332e06ad37501726c5518960ee33198e6c20b8ef175ad397094d58864b56c5a203857e94d7e18dc05b59aa5cb28b40ed30adc53eef4ee55ca542df669f21820f8d146117d3f9dbe546d401c5d890b00b1eda8abef443ad5023d7b1e9190816ae1e85152a001a96c6212b32a65c4403c46e00e2e7d064bac7ae3a388be975282a75155d1710e61b50b72a8f6b035fee9d52b5db159e7e4358f2ede1beac99f42f5e36f33d0241054ceef94c3b73ca96b864a3d218968d69dcd29a05d7c1449d903e4558db51000f2cb25cdf3b49f717690b77e7efdeeff6519827f29a9a6bd9c8760cfaffc758a463686cceed48ba43375e62092e20df53d1a4357e27fab1bd2dfdc0a76034ed2421d7048772f08364954858517167b5a7c51ea0f1fc7689894c12be4547a70d4c7d90858167dd1a4374b875b8466c0974b5cc455ae5b9ec19cd039da69c2ced14fed54a852219f1548826c871d9424047ee0f5eaba3e949c3a832e54e551b9995857ac8abcc11c8b4b3206feecf11e782c62c92264125592916c181a2c28ab02cd65865587eaf5264c663dc637307750e6025290382459eb8543a53507fef5a94b188d7d855b03d9585f05829870e0388eb1e7a48f9a248ef14f1060038fdf991aaa400f0a5a5d67e53eb5e6015c173f6dac57692a41d1e32c843cc601f6ee16a72876a18866a89da623c29c2d0ada4a54252b7b5b402059668aa7a35b8b821e2eb4b837ac2f590dba4504935c02ffe8a5425dd9ac643b21fc20a67a1ffc633ff4a0387acc44f4104c4f59e6a84f16f579f85fa78a5f24253cb6502fd0867f57ef58107d4d21e86e2eb53a818633731315be9326c34003d10d3f5e2c0b6aa9407c2548cbc7e9c76f64eefe5f3dde27cce0a34763caa357655485c9a7c6cd2c20acf0f50b0da09efb112bb52f9e906c43fb524b053acfa3e9132cd61c0526cfbd70367274fd688433d4ca624a27d391da81c0cb174480ce312dbc6887033d1fabd4e9c2c8fdb396b17f28d5d33a4a429b008cdd1aa6f63e20d9dc8c711eaae238236a0fb80a99807cf0136fecf5377232a80a0fae6290fc101b3d39991b2062b653e89ae7b4eaf9a9c7c32697e645e72a31d9a1d37a3e17bdbade23fc457e826a6c46b9eb9727a5b9b6f71c17c44ad65f5c8adc0274b60cc359ba9ab39c11fde7220ed0a1e9515ab03b16deb9c402146a00948ede3d642ee887db37c9604af92053d4fd65ae13abf6a7142564cf8027d02d87bc14423567545cbe10fb265d46d798a07d4e7745a2019880543ecfca15f355396897c150fb44ec71a641398698c07c545e80e394ff39865c1596bb7da137789489eac752853a40f9cbc775817caeb4a99a54a259f2f6592ba46415bf3e0da0e85542fd5024b3a543d8237ea6f751ff57fe04b74cfcb4ffe796b3c550761b8500eaa37403c175f7771b5a15cd09f0a4da7aeb900677a932baa6cd208d8839ad65cddf5524babac4133b72f2491e723d4429cf43122edb0a7942cfade9ddfb94d30f25e0a4393667cb042675635418d5db390030cc60373be5992aceef6f11a2d25b4f7c1e2f251905cf9413c424f62eeb1aa4b06135cd4df116812015b59bbe1a408f50fce0b1d9f5c0c70dc0fb103e516459e2f410adf4b448b16c027359ee1bcecd7bb7c8e3c530c88430c980c96fcc292e035c42c200842eed918ba34f55616523cb1041c080dd7e3da879249da3c206fb3e237d72fde996cf35da710cfc012b271858a9d58e3e4850ab99386747eac5e222a7543997477e2b6d92c3dedfdf242985646c571efede75f464b529d51172749eda5f862533a93e2cacce7041d6f01fc064524bbf08c4c462aa16b956b1da7de9ae5850bf2796d9a0294691153fbf4a1ff30e5e9a813fec8e54b357cf6e36a02d02a2aaf713506eb061256afa774fef977b0e49b6f00c4b04f474e497c254e1c6c6ec3bba4e770ea8841cc152b347abdde6e376c31d0f878aa2fd56571091c60898679c6e2654c147343e983bc92bf821611576c96e5e7ad5f1a2beb47d5c65e87f68ce7714bd0aee87e9aee1317b7359e7bf0af3bef8b70119c21efd03a28fed35a866404c83a9ae96b99e996f9088e69c32b0c9877c571272919fcd8e1f70c59042deb88ad791e7b0fd954648b1c6049d651f5074892bf57dec59010678f7382bd15839e00dc9c00d5de2333c01900fe452fb3f9884482dad997d467263b386d90d22cef8000ff51ae970f856f5f3d26b35714208c05bb1030cb01110cb48d8f2975b7db6aa04890014a1efdb2e6cd3301b41594b82f813c1d2fcf5dd26a2ac100acd2b7d5d9e449b2d675ee36fb12e0c36a2a7957613bf61ea60b637f2ecd7e45aaa9f17b3f17519e9fdafcad854b1c5658f543f39aff91baa2cdb3b2e4caa597b642768c2ce55c330de3413cc21f81fa5d33d178225d65a6ce29463383e3c3c171b8f5b06c2a8547d5cce9cfbe2ca104d258f7134bb7ec51b56544e9a441092bf9187844988826a5f8a2eccb0d7596088dae283c725de4268793fe13f2e0adb121b509413d230452eaecd3f767b1433650ad9690c1a215d1974f321e8cc928232de0ffd9d6fe7cedd18ff9bc2456d6d83a1ba4c98b67e7992f0414e9aa9a4dd629d67a699460b2fd2531233be07c7669a8492a47043e67b0ba3dc222e8529ac1654c79916fa584c0b8fbbf51c3ddc27e697adab5fdf95ac68e1797a42637685e71f42075b478f5f35f630eac2f37117838cc069ff77b4066bd12e82955e307a4e33c79cd94ce9128b8d47ad524e4562994e012069afd727625ec153157c7e3b386f388e9b5336f891c39c69cceefb814543347d59fa044f6ba79ecb6cb1640bb7fa8b088909c80fca03d6f49eabe7d5c820a658e7f7ea3f2546c16667a001c9c28b190470d8352ee3c07071a8a55fc0d9f98854755e48b1241c6c984eead5ba295deeec6e582ee7ac7ea48216fbe386188e0dc1871fe1b8b67bb2a9aea37e43fb29f16c944d438e52e38e2a4158d592aa67376d5bb921618b16775ca597d5deac8b90f329d8b2258b45144c5222f9e2548a244d61810181838cd9f3a4dc88697ef4bb42e9e1d7e6160276e46e87453c0af22d876783508919a9839e51878d6af62d1d556c835abac7bd82842fd2a72d3b22d48abc1f5e2217f74eb23e54ffcc643c275b273658d6074aa53715a0f2af256c93b51cc09e002653056d7195c37783db9d8f968dc1fb1ebbc10ba8ed21c82491529be4e493e5666135c0b61178167881f1b891e062b052339a5c5862385071b771f96590a2aa7bd17f8ca5095bb1349451bc2fd98a392848d267813df3d8431c0f93412c571d15ce6b7b74fa3de988e008c74de541660b811707b88abafe998aa8cb3da836875c4c7863db9364be52158f93301eb5bf912b6a705f024079939893a99102fd21853839c6aac44879dd106ecb3b971da5b99c6f11101ab783c6c657ab393b2ce5781cf02f8045360e02ab59af7567577aa53e758d395498f95adf708b6f67b07a711ade36c9c9b2fd33e84b1dcc5f29035982b82563c9ba9b7f21ee1c9113a991a010cf80f560c575c8515db5eba66b364aef590b7c282ee9769950b1eff4e1839b1de65bbf5e83352f0b46f8ff48d2ebb63cb53f133557c3bb7e2875b90a14971bfe78274def8cb42f785df6925a7582cc0f964a2bc18cc5540bf53e2461d9197927f49f300ec7fe74db087222874b10c97ecc14f8612247da0bde05b4f8d0ff6d606a9be49ea771aa493807f7d2546deaaf9a0a584282dcae86af8bd81fd42b8c327df83f224701dc30510074ebd5721ab2106d36892a160d7217e1597ae0a836941395a2541933aab90c0eacfe99b6dc9c42b1293e636cd313c3e3d477be8bcf1c7fbc0f112f2f3164498bcf4d45400290b7e54503ac199097aa19dd9913437a5708aa69386d4be148f453c29db53c7fdfac3f453660d2d09d9562cff10565bd99810ba53639e5cc30ca4a19ee3cf6ce8818a5322c208bf378b7184bbb8c3a4644a06bea42ae57c2fe1c35741191e5d97e0e04b64cd1b84d8cb29f35c1917017f2f35ee73a3e2bfc02cbc8e8544a513881af1ecb33dd46c2fefd0384dfedb49a3e7370c45ade2dd3f630ebdaead77735db4e8de7969d4375e21549b073d3a79b54e25b05834816056af0a24a974da9584e77c2482718293b51a407b46c3c51b490853991c9ad97adc1775789c4d8637d812bf8077aebfbb688980b21ebeccb49acb123e943a0206ed1a6416983812e4ece1ae7e5af888af5f630bc6ca361c76f4afe066e6fe2841e3f6b6a32b5d0033283be828349649f2875d72e2fc151bdf7ce22af8152664bb576a5175a85a28664b406ca2d17b2e6288a95eb4b3ba3f5340a3a86e2a249ab4cd2411a11ce434585ca6577bbb83febbb41ce5c2dd3856ef7e4a982a0eb73da5c2b229d41b4abbec5f3280826fb530d2b454f1928cdd1b78b723d6586d595d49bd2cf74d1b24d0597ee51fcad45cdf4de7038fbd324d31125637180c47cb255773c7a918c63cd0a94a9a3f91bfcdaa029a47d4d29f531b7ba383f57a97317c691e29d6f6c5a07b7d1c51a4943aac095723c94a6ec2f99271297564389685e84b312b5fc315a0e8d58afbdaddf999a86a652940b57535c0f492a8a4f12ab32af225793e13a3025461eea00e2d129f5c55de31323882659d88032ee2b4bc868427fb9e5fdb7f7f14853f897239a85e81e888186b48b087569b0dbb33b2bf1a92bad0cd510b0bc84f76884be8549ac5142c3a24300b22fc0269a3a88c537782a6a36aada92cfa709e2210dd9517b6f3182da352326a9abb65f1d6bc8a0bdd6706e5d7f3f295643bc1a3bc5bcfb20843f6c9f6e4bef31b8389d4079632ab29de458f87163a92ce960b24727431d1d0090e7b6a1b32b5302b1583edfb136ab1011e025d0893fdc294f76951c1bbf4e7f779a7f06cf107ccf3af51e5633bab4bef330fd9800a90ed71ae5149409478ad9a41c62b101923c60fd2bc2e453145530faf56d33e78565acd4de4c3b2748f23d47b7b79402df885694d98ea136b891dc8a1ae9f4320db40e1d039dcdb6ad19fa1ea460f3f92282c36ef7d30059d930f06286bbe23a249277dfdd75e5c070e6606f39d3da0be6051892b96c22b4833d72cc1955adf96d31ed8c3c3deac85df7938058f372ad4781e0b2ba7f081ec6362d49c22cb7997101cb57c983afa2682093cc28167f9dcf7bd8a39518e0f94e368228d0d5d904f52e1ec0fe94fec3ce1c74ee337c4b8210ffcf3efe381748a147f8cad13bb72674225fa3bf3a8be9252f15a06b02d3f67f418e0b548043f9622244d8b10a338f4c2ab20bbcdb3e36017a76b230a1ef720a96894ca78fbed86ca48bbea901d92161651404a26c4e22f81a0a64affcbfeace07659fc36cebc45afb8a75c01c2b3816b7bb771edd85dc173b2554cf41d158c64e4cf99132df4ae95a620a6692e4b269035f97621d675176a08181e130e3cef3c4ce6f3efce674b183a199a54fac590080b7c3954e147008f018ce76762f01084b380ef44c44369532ced1ea48a2f75c3c4a69bdcd1082af7d847aec5b3ff902ceca364d923c58a749fafe391e0203d8492674abe9565e00712a712a1ed33a4b7ae102e1f316cde47f312ea12d50fb35af7d43356717d36bbcc08546bd2162283a5e713630d8dc8a75a8b835ec2323bbd99d096fe73d5048e518f4ccd52c71dc87502338a543e73a0b88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7439033928ebc69be5bd33aeaa0ccadb5904556958256130d6c9e0fc510b66d443e3a437ad906dc781b0c6879d7e1670d1d948b1208f49c44f4f945c4503da5e9a31cd95cbadb7025f8e3065d3d7d815091c14ac207e00fa0cec509a08afe6d06da82ef899bd6b6f8b74f3f0b184948d973f558fe1c6d14f4e148a7436608ff8bbc1d8ab4555ce935702bbf3530c3963c7ed553501867990701e1fe1d4229d25702f313b13a6d9e17a2db475b2928f547d82e38ab0e359b992faa62eeee36af7b8c5febc3562ed0c1593a575b12ac493b023a7591ee99823b694b457e8752d32ebd3812f72f68d0ce3e517297a9838c577a96f4e7707bbb01bbc251ce26653d36a43ae63e9958da74cc950fa41d084249f12b1b071854c99c60bb2fd75846bf0b61d929700c39572d8fc6cfb6d8f45dae9931ba311249efb29478e3ce0db5032df1b942c222a6cd1c44884395f9e4c7a16ae2ad59003ccc036016912181481e5bf19dcb1df0371d7dda2b70f3b8813557db0d308a14d62f03639b8aafc450ae0ada7a734ee80fdeb3ad3c99aa05cce550857b50797049d5e17a53cf94590eba2876a528451ba2823f584ef5ec2ad5b32f7e35ddf410dfd9eeb2285067310c0f6b857df4546b76855c63ef4069c9a91c738cfc5170035e6075ee3c479d61e387aae808bdd90242b65637d8ca39413586561836747faacc2852b53c6ac93869a3e3982e91ebde289715dd186c0bde616b4c5fa5c08568701b88d4c00af13a57805b1fe6e3024493b017c1f2ad6d3ab7af30d396004b6468d5cfdd8085066ecd1722e961fb1fb9a0571b3e22647baa876414efb8ddcb4a6f2f2a0f5d3e41cbbe00c30e892490a39f330b11be55d6426dfd9b0a7948e30bde4c16abca2a136d41ac8f0e3b7c123c0ed9898ab7ee7cba835389990267b373dabffa60664a3de08cd36c3fdb59234ef43841e40b9c5c4c19364a6c430ed8e92f51c6c301c723220a2222aae703ec8175ae275163bd2199ea37f39ef0960bdd6b02c4a7bee1ea28b85e5a6a94d6e14b4be6947a4ac62b03118189b31052b863a661f7d57560cbd95c4cd97fb2ec5ad5d56b0f0547ee45de93191245ad8b4fcdb010d0e4ece51db95dba8829f3a6de5de59e8fd97ddc8bbd1e623b507f50c9417d9fc7c5a6d6c91bc77e11c08f65cd4ca29670352b4e23ba5d2efb2a61003ac1f37cbbdeecbbfd92c6718b3c1eeb07cdd9711c16a0bfe7653dd167fe3e908cb3267016e1884129f641263d2b8259c3b74a7d1a0cf2016eb6790632baee4db1cac92583e1f872c5f5e0499ec1a1ab20ef888da6cb68dcdca66430385fd2da6f1ec95bc08b1acbeab4aaddb19e168910bc362439dd52be67014b29b5e4d31aca9149ab5089ad797302eeaedcc2ac4f9bf12406238ca63e5882764bf59c68b876e02de9cf539730b7d89a22edd6854cba74ff2945f65504f85a6420a398d41e2081ff817e4ce3b33c0b892bf95d1e5e8bc87bf69caabd5912d937157591ba28c19cca079f8182dacef8411d17d92b22c908500abbc101118187c1e8bebfc5d9d680d18aa834c8fe2132b378d32dda311acdd3a47d3bb59647cee3491ee25f10f2a2b3537e61b70a913f5dfc20e36ff0c44470aca59c2ce7b1096bc2498c8123e10af0d99053c46d43985d7a7833f7b18deeef4ed63a5f8e03db1b6d10749b63d12d9aa32a9a7df4b3a0032897ffaf8028d4533eb20fbd9979adbf14fb1ac0d9b4597b5769a3284cbb28f377b5569e7665950c029c2d87f9cce3cb28cfddd5795d40437c083332e58cd0566016f75fa269f1451e85e761300118c5b4f6b82fbfe722cfd6b2ce8e7ec889a6c65d1262aae987b8f69aa4eddda15e2fbe6b0d4c0a02f44aa555e933e7b21e7b62adeb28369fc2f63004ffc5c80e618a961a82dcacc4c4b9b22f8d71ff0e5488b45aec48f44c0c5fdf0bd8c498d3a89a696292e4ce07ecd14b4382e479361d7d130a4dab89a8c44b95b79f3ac6f246896794cf91aa7c60c763994f8dfaaeaee883c02b0abfcce7b1eccc989cc6d4a66dd604948a25e8440fda2136e0ce479154a559e0cdad015b67788d624ba2e57fe81aa0c355bac30af2e20eb6a21667eefc25ded89f2db62f5477db77a7c7ff467aecadda448354af1c991cff5c9ac76a931361bcf30ade653761eb65e28702fc6713cd4bc3b13d376a5704495b042ffe570dd321981cc4574d0c35f001d2ee954216753b9da02a23a8196070888d0b11d04ee6fb75109b1a83192debfd0e598819d95a310898fea228f654cc0155addacc5e161dfdff03cfa3fa2f17d50362e3526c6131f60133a51d63c632c725c482d05dd16889d4e7d3e55fdea5630797624fb653e649c1a13c502f32426a1f1ccc1c7de89c1eb5360eca415c1a5c50b13e18944ccda86e7c6939965730a609ebf1fe4fa59aefe5c4dd8c4b969416420d6b01d9503680b7f3f4514d9f85c46da51ed5dea11c075c099ff6a0a06bbf1e8fbc24598798a4b405819f67561374d9572e2f680dfc8cef651ddd80885f993836cdd07db752ae7a8e50bcc96aa647201d872da15790b634a96e027fc1b35dc094058b56ad7dac0e8ba1f42c7e08ec0b4a49da91d6216f2531ace55c57caf2922f5a660677ae58acde4eb57a9559915a5b70798e9b60642a68fb13256bc16e18713436162c83ac57cd17d69d60a0c02cf09ef4cecad0ec1f803378eb90f4fcb51c30fcdc14b88974dfb413a697fd717d253207230ca62f41bb6bff476da476c442e3fe28db88ac5f81c099a128a25dcdce2eca6b3d545129c0f81ef1ec9fcf164396318df574cbbabf3749eaa9590fad9f35501702186f79e866ec5e55d93ce01ead9d702e92cb1f914544bb992d700ff497884f6b321d74c90710c37333c16124f342c3b1518638fa1be1a6464b6876f752c62a851861f43f8912e218e5cad5868c733e7e1feb4abf9ff618487d7a04b51256a5a7f2b4b9450ae97df7aac7bef2bea097eb5e5cf82a206e14f60e584a11533d440151a7057140fcc3bf0c44cb5e5052b8ef06dd2fefcb2240d7b1b2e7aedb7abb372ee19d3b81436e8490ca32317f5d34008bea8c6186a583b8eeaf99dba5cec5c5d9c29e2b5881e04e3205589c7b63c5c83c75e16d8211e8d4d5398d52b35c3c5f3c4fd0244cb33eecdc3b94bde6e72d4b07fb02f4be40ebbcc84371deb56828933fdb70f76dbea1d893b4a83e46a5d72f71455ece8c9ba0a0901bf8a21a3233457d0d6bfad36281f7c026f04d52a5c71f5fc60f6e547cf4b283268825a8d3418afdef16ee3d5f8f7bed51784655dda120496399596c0f836084a002061c4cbd44140d1c82540128a07b72a914a77eeec3e48ea12d2787a1c31691982b8fc3058fa0224cca2247c123770afe42a4f3a0f6e97a97768f75ace3153f5787dd4dd5da3265d65e29e9430650bc60b83a36005a6e7718e568b577332404c0033a999ab3a87df487090defccf2a157df62ce628d5a6ddf3488eb299788b7e028215409f298d3d520e658efd8c63e26c1df6c530f711facda68fdce47fbac6907c8f4408f094d250cab0847532170aff2909375ff3b668708721d7319525a3d2506bff8660e38d945c234b654dcdd343a86e201241789f61964ade1d4bc728a9de3ef14650e5475496cfdf43b483e9725f92e6efda646bd49aa411c53eba15d04b97001428c48a2d62ec137ca1e0d738e8716da2d903ad9a636d958799e3c94746fe3cb97fef6deda221a2f20c8c5a0559f002dbad98b066083237aa41b77ed8acff220d387b32f3bff6b19ea2d44fe47b841fde2561b1b45236e41b6f2ccf00515ca6a667837f9dcf00fa1a1ec9f2b8615750e2adc50d03a26d13d8a94eeec2b70ba535aca5e6b51b82e895bea0a0ac07782c3b28fab7e1d6f17ffdfd0b8a7239902abfafe84721813f884e05ff4d49f1dbae78ecc68b2cfb2427f59efd7de570d104800231c3481cf21dcdf227153db0d384eaf43f9365441d1f58de200f8e757a89b6cfaf7c935e0fb0cfaba4afaf508c65f9b80d20b33fc700e37d1a159e2bc75d92e007c4b8ddc4b0edd18fd258d07b17bc2e6d3fea426fd3d4de362793eba2827b9e263d2a247ed569956ee3d73cbaa0d52462a3a901eb86710f05ecdaba9bbd5aa25cc2fa9d32853ed568588049bc53097f2ce1b484ef7e28ba2108bde58ee0f1f7d6edfacefbf648edc22b031728689cf57d074872cfe1c4b5459fdae5cf335aa7e485ca8306e54f360631a1c6adff497970caddc493e56b39db683112d0cecbb0cdb30db8fa7cebafcc85bfdfd560d3059e205bff0af7c5606d9f5518e6a4a84b3ce6a3c5bad0874256453b2e380c862c0845c6ce0e81236f65755e60fdc06ce73dc60b4c3166f268426293f397af122a4664e2c65c3d8cf8ede21c012bd22264d99f9e96ebd7fb13681ba324302cfb2b26263d8abd83d7b33f967b217e8cf2097fd178886cc5818357574a36f57c44d953566dc432868130d91ce569b8db3d9f431c09a180178727685e2dd9c4af40c4ab3904ca1bb23f2844c1df32f694a3f8531134bf5c469196ec9bbdfadce7d57ded5800081c6ed18ee7a1b061aef3d623a0d7b2c503a8b59149ab74584e148b72aa8908253802966149e09ebd1c10b8c553d14976b38267a9ba2b6b26c73c42e178dbc2c14629a93177ceb24ae343f75d10c825d015507925fe687bb42c7c7d5061d57267341abcf0288cb2276b530b33ebb6f28e75c73339641d7fc74ac0c38dfa507e69a3b5ad711ab2db946787b66b15348bb18ac5939025e2cc09c3dc1123164020d386292ce6c920a692dde5a6ad6eadaf7a94287711fafcf6cda02abdc52426ead73c4d14b81c2f954ecb746ff51cf45bd6bb92bda0f3ad0729a0dcd42ba3e6466c9d18b0b6501dddcf43d6529041c5b86db742c2c65c46e271d35b37adfe57b02a9d3bc538e62fa58cee6e0e2ac65f61ad716511fbd2a87c1611cde49c4c4d35912fca78a668fa0196e2ec05f028592e784d2256ca3b5842b76bd94d31662fc45ab0db17015f7901bdba70e343c1f79565f4a9b87da65ba98567b4c4af218364cf8a6e7cb2b4b9fa151a93e37d568bc203bc6422b391b0b6f4a0aff57a2a4ceb4cb4d125ab76280ae3c74d1f3a6f85ac5889c222ab01c6d4f816c25a41a5e65a0fb75543b63a0a9c05a707f933761158c934dcba8f2ed0cdec3233e7ae2c672caa83769e59330ec50849b263835666c5f5df8daa344b194294133c7d97aee67df684105fa1aaa6d2e7dce80229e180da85b961eaf446067c1cf9cfc76dab5eaa09c6d7838177c81de2361480fb014748d674386473b0fee925eb7cc383121c1d44727d6f5ea1303e9e625334c37d0fffbdd7586c6388695db43a7fb5fae20d56d395c271eec758f374c774a4596f2dacd2fc2b4460f36a8a12dfcd1323ebcc6981e48537841e2da019d19ecf86cb82e36cbd04023c5ade6b3baca6055390af6f4d992f60c24b8391d403d72ed2b7f8aa57177745244d9b48af3d3c19a463b05e1c38e0226c35bc61069d231fe19cf12295c908f2adc3fbe6df53ba95971a3592fa7b1bc6ebcbcf39801363d22339c785449e517eca445b198b946de8454fc1ce534a291d41f356d3773d4e85b54486e709ff11c881968e1afe85354972ec232b80372c92b7e59b53856effbc37b01b17effc87934ba0bf529f108b2df8f2feb4e453a6796b3cda68bf458810072330d32f6d0f733b2b897c682fb566c600c7c11e2b1e75f0b6d505e3f8633e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7043eebdf1c3eba23818e9e94f6e562b47999cb8236385fba477a98e7c5f154fae4398a3fe406dc93ed887cc6d8f01ea4d9615d1d0053423af07bf2cb681d4b6860e4f1deb18f5c8c9afcec96eba6e057d7b694be31cc3d10ed846a1e169cb1bda1ee82f4b05d684446e421fa475316a722cc63630260d9fb912cb5a96510f780ed5ec4545bd77872082d34f8f613c13a2f90a395b7abf4c627523cd920c5352d13cb99d66f243488624ccc7939da098bcfad21cfb5b1a0a665854318f9c08ef637b9cbe8240ed47ac7570854e9c147c4e3affac128738b1cf9f241dca8616292d030946efae89bc32dc3d756c84d79dcd0fa3ab73dad9f8150a0674924fe444f67f4cfcba17d08667fcca7c63f61de27d88736be7eb04a91da78c4a4332df2eec40a8060166248dff0c246bacd716ab11541866dbabcf6d838eb72464f008b6e2938358290df6ec89f76ca2c96b23b04ec430ac2870524d3fb17ac9858a5c3f83ac1b7a4fa9c5c5ed07c49c5d7cba14a504f3df597593e1c3c7220d6bfe5c3c3afc218b22823474b7ec12509f42bd079fc51b87210a9a42bd5f9dd6b49f8727656ca63a5ef5df51f77be27e6bb94219f2390461c0d9434586e37d0f8f87045f0ebda19cfc29f52f5ce7df81353a0c6a00d89ccebb0d9b4f760e9a945ffeb4456fbade00797314ef238cfdbc9db18a62dd8c9e3583b01baa18ddb209a4f0c72d7f451d3a5cd0b633ee6331e4815d3eed273a150c31e1174424547ef83c451319040bc6f906f1f6a188ff90c355d41546c446bf95078f24e0576c16bc528884e817a4d16b802961442a57f559fb6a6ac1f843b6d2ed27cf18a3a47965f67485c77dbea178ac58be7dcf8ff8157699cbdc715c2c1dc198b14b037faeb11564be78b9f3e397675e7d9a1bb5235312aa32cac8e3ffe5a69b8d147f6f58376149bc059a138f9620c322912ecdb6d6ff4aecf5700dde6dcd0b5b554374e718e184149b7fe527648b09f772e9a5914194020546f80b235211662bc54dc4d2834408c49af68c4e50fc3f36cdaeb1cea943c63562c47e1dd39e4933ff5ac9f8829f84cbd3888b6857c12dfc8f357edd70672677ad2749481aa6786a41b681e60bfe6e3e2074984c2fff9ae7b571fed195dc8025100712a3a650b10d77510cf5c1a424787cb7f2a8436e418b8eb82cacebd600c0e2e82b5083b6b465257f3fc57f124c1ac7549d840f120428eab004bb397726f3a903852890a85c9ca127fd49d453cf8d19874f163102a287366e2b5bbeda910abaf236efed4800be838a324af1739c0d6fc345517fd797ea16b8a699678737fb926cfac5840edc7a3b66a7c6375281479e6a048f6adb65df1e28915b4b08bae86e80040ba7f3d45fc5a9396399f69b78635b0d7a3df20c8d41816e56e31328b4702101c71aaad2d23beae46635ace6bcc4393b062292452ec9b1531563d58154cb41129a04577bd142100850f45dad688040a0e137028898d005807cd4b9ea44d7152ec7f8bf856f2c9aa262a5a713ee254a806f7ad327b26061a9409771c6a749055e277713edf32c0cf9a7d565edf667d4779ab5f8e41df647cf5dcba028c1276544ce1201dcffbed175c8fc5ca7427415a607ff5110360e572ad56fdcc3c20be624f6aaf0a2f33afd421ca1c0ebec093a7bc2b23640579043328a05e746319dd01e2b47bff50fc26ab8e47669917b880277280f56dde627f6bbdf503ef2b829500f03b1e33e18d45d8c6ea8a9a02a8f25a625659efe4ecadbaa6d20124daa67244447e7a4badd377367b0070cae4ed006999d7a9e0f12af1bdbdcc66ec1b91bdfca2c51dd3f0d0977a1b1ff4da1fe9fcd9974dffe04ad2f7faa72b362e210fa0164ea4a33c84615cc0a9bde5af25aef4beba72a520ff19194e3654cf8382c620f501ba4dc2548f305b96d72118e1043658f0b7bc923f923c602565f11afce3fcaf8cbca8b4573aa9f545340fd0bc664c56f5c1b5945e87f14992b4bd4b52c359057ed4c94d2d0d5b255bc00321de2f7774455c0f96e29e82d7517debe081dc695e679496d7accaa6567867febc6185061f2496a4fa685009b8864d7a9d5b7415725e3832d5966c409348b1c902134d672d3f84a50c69ce8a985b22100c9383b70c13723f3165b3056196f36625abcb7bc12065ec345ca5f99b69f923fcd8a04038e8e79b588a02219057c69f8765166449be467b81fc5c74a3846aed295503aa0a877ab1d219dea2134b9ad9700e9f68899edc676290e9020d774afd485d00e02f7fa8dab81340a2f4e10b895563eee961109edd53c1e5f0dbeaec60a92e3d471eba47380c0532495d94463a56fb383b6a6ae544d2dc24f783b37683209e4c4dbf35f533e30998bce297c294fcb9fa47049724b54b71264c611651bb7660134144fa0e1cbe6265e23848f34cef546cb4dd467cefe4068e099058d690fbebd8ef09f111325df84a80e6ad87baa380e883aaef685fdb191a4caefa1f743347deabe1be148722223456c6fade25df54e55dca60d8f4d5555c367b6fc495b8ea4f3a0ac176f5dc31baf583cb0f121347a7a8a76cb1c26759f689d3f941be80ffaa430226a98e88d865abda521c2704de2ed164312ddf6c922fb2ed07a90609f6759b6f8f37c5adb7aff109355a2e603df2a750fd44a1878692f6b182c3bd75e8fc593981c1f5f172e2b5039ab37f65d4e9ecb0317d0fa0dd9289d48334f01b88de4c953cb4af0f0e949ea6572675e9aa2ffcecddc6b28e2d5d342cade2079f96409dc069b04cf02187ca1b583df46661109c78b63610b89e0f397343dfd0344d14ede53e69f1c558f82b2f18ff3fd8bf8f279ed42c27c60fd3c2dd6e0d87fac35988f3a6af5412b22b7a52cff8e1920925ea7fbce29ed1853be524a8d8bb37fe6fad1b7b31c4b28f5f50084a7690b883ac3bd2893c25fcf370887d21d6258be06ba1bc923f186b36de0013e53351b9e70f5ed32969592e2d7171a26b28b42080ac3a8485f37da8b845ec1b7fad429b3dec27d668aed1fb7f9b156b9a4d429e7e8cf11ac883da13ec58a8ed7bcad9ec243ca12ebabd8aab537c4689376058769f6ac09147f74835da6c807ed6e5f2979772f50a37ed326e572d425bde61fce7cac3566ac724ca1432c5eaeade31f2fec758f631414d5720ad9081ac18cc6e2a1b729c7eccb0f9a722d6efb83a1fb61f441ebf81cc1ef2c8067159b396c145c667dc7cb4f8494f712f3263f52ff7fde267ac6a392731e4c241ab739a4d46fd5eb0c634c6e4085a2641602695440bb31b2e94473676b793ada75671ca97c7a7a627e491a1f593fc8e56f7709d20d85bfe22bedb3bd28767d2b3800889f65f70f980d0fe009cbbb19f2e1d1224873d892066b4dc9a14fe9075fbdf179a55f7bd13af932f95308ed843080f3fe0c479b02df0ad7e5ca5f19d18009b0ce1d8ed91bdd89765add84e9e20685932af37f11c4f226684172688cac13c917d8df26a558dd69380404597edcda5c4329905cd9f8d4f34043ecab1eee3cc557a2a719a0321de72be2028b895b94c8a495622e67d0948e7c2ab3706a35dc7f88fdd7265bea9378a34dcb71e0d5198601da2afc6bf263ef24b0a62e6aa846e4a798d945dd4d57c7e6a3cc8cb1cf0d8b696fd76907315ac2f33fc682cf54c74927175f94b3bb90f4645234fd79f42ec294f73d22eb75d4b9514237615c79833195d3e978936e47aadb81cffb7ac58955a7edc8ce3916e05355346bfe15fff567fbb6dabc4181c77565dd13e4da62e1842543ca861894520325a568ee26126cf49781ab568bd1476bbfd5edaa8a1752dc3ffd153d36de4e29d63f57b66fab9b3df0084efba82b62d32022167c278818187f0c6f126dd971666d2b06480036cf460370e5d8f6e8f9604ae22842e623aa6a3e599a1730afb424cb5c80f00815b702d12a7aad014360b0e7ef8e6bdae0a740151740f0aadd5ac68496f96a0510117a1ee89928f60111de22c5f363d5798a76433ff651d35007df4ac6175937786ac992d71144fd2136a415256f3809d3b4ab4dfa2a177f02b1001399369ba37ec91e7b02b2adad32becdbe6818ebe64e58f8c8d3f363cf5a5cb8c2359c331871a1f56715d94e2020ae59539de389bf33295e01d3e231ed9902feed37d41bcd10144b13e62edb7ae0b1f19c7d71c0745542f5a8f78a373b1430a0f957e5b1f6785015ce97e2ee5c565ec5f6b1f882722f308f6dc138ab2448c53545b930a4f0c83cb726032cd407742d4aee70717055b31ab6fb0149695764bdc9d0e7d3c6ae4495b0a73cf3a09799f5df37934e5df9408fb1be619f4718180744ff186d6892bb1350f9fff7cfe8ecd9130e02d169f93a556dbebfdc75c3d40240aeaeec4c58bf7297c9a46bba0f71c7df261440c56c5a205f4858bac9928ec7c81b66439fbf14a2cd46b6f19e3fa5beadb1d77586a98a3e31452ee67bc539959cfe3945a783ca895d3f314e8adde7527d640a833ecf46f6e09191e6e438abc72395f9c8e1f3513fbd4aa474f647fcc73af40b6e74b05cd32071498c5380ed087e57860709960577bcfee8783193714760f80c6cdfa9374b20a9688ca319bc10bbf0d8f0f4783223cb4a5c4b748f9c0f263f48e3a8a60f2b780e6f4df2097f88042a4cf9aa6f82ad5bb04a2a3bd28edb9d1fdbbe0d2f2118f4b105bf2cd58901ecef868771f5ff2c9ab5b5d51060a0acbeb4c3a0903633649ca814b8648cfb0e2e4fd738b216ae5a68ee0b4eaae1cc0c08b145567a66f798091df6d88f2af195c581b7338678c0eda1fef6fc8b6cc7f7a0d28bfaaa7b2bb77ffd168cfb891c69cc089d6ed58ee4949c4b8d217a219ee944a0182df99a0ff8b243d0cc6a869897e28e8ccecc3951f24cb16cd6cdaa6fa0ea624a5bffe40213cc5baadd97d46b483c19a850e0719aa4ea8488535d805f1fbc61778ede4f5596a3388ffaa72dbba6a4368b4f86de8f96daf335688ef063a8ff5999fb53643ffee3576b94e2855d180a04ca0dca7eadabece876c6671d6f133c82c7a53ce72b3f5e76512c997bf93da7c5efee36bfc4009846fc4b9fef148b7642533f2892615fbd5bbbe2169a7d7d4fe927cc2c1b172cb9c0fa60a9c9be5878bdfc40152c07e49358be9ff7aee1219aafe502ab257b3ecb7a4e5c4471ecc8b4a4e2cd261543f37f7a27348a94f6b4de4da55337c0b260e3815115f33aba62aebde73ea3103f85851c3b754f80bceb7a0efaef02504932b048e5b2ebb5ffd2c25e070b419ca4e1351645cf6bc8dc89105677e4172daa83cd3fc3afd820b560f0401a9b28c28a0772ef06b3fb8a64594751e94d50fb6a316ac131931dfb8f103c60a753d2bd3fc3db855faa11e4ff191c61cf1a6b4759c7744d7cdd6cdb8c308bd12e2ef5655b369e61e1f315362c64ae3a5f80caadd197427ae3b1d18310ed0665ea864b179bfe8f2ccf6474ac0f5753cb3c07be4a24cde249e5b35481f4b08dc8d0894333fb1a6f118e2e454a55c064c2c7c4b903915f94a8bb6738a70089ca522aebcf3832d8f9ac696d101bd07ca59fa0cb5037431bb94fdb407c3b8c3f515642b43ce52012734e0f0638a2ebe99d17d82aac2b668dca9333f6d9937c928d3b1285d494c697cbd9a7b321e62117ba524a1f0ec643633bb5b81a3f248179f22a4051ea3b0e26ed498000e9fec3d2455177401c70fde85f213503b7757f0085ceb3c157d01344ecb4dceaa1e81b243bc74a6e2d77f92091634a3854ca46e9c452536895d5b8bfebcd33a54d167b701e44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9528b1cb5afeedfa1cd173145f733755566ee38ca23cec153696373a45b4c94585ac6b4ca1c628e7558fb3b1a66ae075c5c365761cc97dc3577050658b64df05bc1c8b06c0f91d415d93c35ba2c1c88cff879829a446a08df4d6188b8f8f3bfac021fef98bcfa91e6e9432409c9e07c3467b1a545ff0bde28c7ca02b75a06b364a7460332b3c7039203ad271b7ca64c7062de701c7d722afe055b112122b76d3856b31ece5bb9ea847dd26fee3677e5a859ae078798ba20dfb006b7ad72660a140ce8844cc0b247789fa9264f2f699f0c37ad6b519f9715dc40c56abf6c7448aa86b95b2ac9a7c81a737d5f3aefacd692fa85188eedfa68692856ddd6caff8b5d11510d66a2e01fa05ee49954be62e09c7c850403fd095ea68afd69d1057e3200cc068359b2814981ecf77c3a64cfb347d654868ae676572ed959b7ea73ebd98849840e63bea7782c8ce51670f7501dea34bf577e2f78ca97c5dd3c033d9531fcc0b0f9b07d59b902648439993342e1f6fafb22ce85314448025c9668d6b11838b4fc8412716cc6ae4d0be133bf1ad3f360158e85c35b86b6c5634f419ee4c52af191cdf38859753f4d22cd94b442f29ee964518ebcfaba290237976994543bb6ce36d28185a28d2d55f868969993a7395a743ce69c609d76e2c295426becd3217e1c47ff8857c7bfb379f53d507c49fadd9accd7ee1d30bb38befd170cb4cda43467c5dec31d6171943ef48c8276ae79e8b0956da32a43b708e0cadc6e59c29d18880d8dc89feff79d1235db78318d0ebe9f18826ab14a117cafe44b846388c57061606661bfcc8e246ffb8724721d353587fd5e5a0d2332633b70e08c7433f777d8071231adac6aba3be8ed43b79536f959fdc69dabd757e16b649a912ce8480694467ff1adae97ea19d1da9c37e3f6963b2dedb83e90313d73a2bc331a39972e23f6472aaab65182b192155e99b0ef318cd714fb9015e27da70fa566b59b73aedabf3a45fb1fd9869e8eba49b7f50ae2208f5e2f98643d2f223196bca8c9a4ddf1500146e43b3af02a2d510deb28abe091546ff34018045b172344a341a50e7bf5fb84df1b6bdd08a841c527e98f2f1d164e0ca068cebcef17268eabd1fff5c69a1018efb7405c4de7f1b1e03a6f470e64fae4f1698a6366e4592df050919143280f350e3229d014eee2eb856e1e08daa011892322562f8891238087f6ee6f0361b7e27e0e990706248bb2c7de53e0994187d5e09e022d705c7e101b96df2cdaadf27d44c76505552336a903986d914c587a989413628b8b489d27d6be1117a47318a89818639296e9da1b6f45301c2c5a285fb0c4b7044bca2dd0483b0d8466adda597ee0c02cc34a2776ba88d85a014e26cc4276924c99f41481e05a2d05b59f5dcb6a6f4896ba2c0e50a4a50efec7b0687019a2a2baf90aa353c82f2f618ea69b04002ed12dc2adc412abf9351dd363b736ef6ee97767d5d3658204ee9569dd408038d4bfc897d31ad2cfcbd5b53f3ab9ce134b13970e0f279f98445a819e4b0b7f12b778178796e010b3bea1009da3c0cdf9754fc097bc5107d6221469f8a04ea7520bd3fe8c88e15aa6baed271730aae482f9a0e4ac6d65744f5b40eed99e96542900c96b00e9e6d69ee9eb362afd48d35ba0c38e5df91fc90a8ecbea481a11c406dc10abe0b4b3f32c1f4930f4f7a3386e6802d3ce7b3262331dfa8922e9b3c4b015eabb4716a94ecbb8f857e5c95a78f71b06fa63704137e2c3d35e910f71cdc2497d9ef3fb139fda443b7432f0df20fc0e95173daf0fd6e9b3f59ab764045586e57f71e8abe21805a053b195cc438e29134caa417924c2a67fc59faeb8c547745c2398dae23101d1ac38b6f92b83cc61cd36ea2bb3d1ae6e14927729d3cb19503bd360c3203b1a24ef6e03b2e0b7142cee77edde9eed29146ded937621d6c8ac19da9c700b363bdd63f9e1bee817146d77652cf5b0965e54a122137356e8bf893166accc2b3b1a6f0e8f23ce8fb0f126553884f00d99a3d07ad9321f06ae4f454e7557c245eb6cc8a0e7ba3937225ee4d02dffaf53f364607b3be6fec18a10920fc87dd0d55625c7ae6e982b61ed702fb835c5eebee7a1f6b058740d8f5f3a317d08f2da2be6c9a9cff99618eb588cd394c4dc3c11d3074601af0cf17383ed2c129b5a091b65ea81b6b90aa9224cb2c0c3c36e6ee8c0b450372555c5fe71750dd1a6c6fc5ae30a390300a928926b01e71da76c9ca0e07d52feba792910cf3589a6b4fb42842c6ab704c05464fed2a431c6cfb0abdff8b588973448cd4038436a7062bdd86b1ded7ec327bc4ee2fdd2541691556d881a5c335b1b79e60663d4fdeb355e45cfa47cbe6a0fdd61655aa1fcb9cd7eb43af2944c7a99ed5a64fee7aff2c517ecd2fc2eedee8f9605f2de57f71372c89561136e0362d81240c21024bfc674d865192884db79c19997593be1ac89f5786751b3c2feff7766ee4eaa03731bedc84491242cdaf38f699a2583e62f3066d7eadf5282a2bb4eb1c614fde9ebdab1dfed84bc74d29b9d3eff95463f68799ebb73879ae4a2169e5cfa86f666f6617891ac5b08e6438749e114d49cd77a6ca05cf78cab3ab0ca8d5465f401f9eeda2e60d8ddf2e7bfb238c5c3b4c9c42b757953c18cf65beb932b7ba9bdc7659f9b13148ce42509e9ec5907ed53b5cf8f9c101a58b6049cd4f4db84cf60c7d7866c53e97a6276eca5393cce2d4bd7fced9dfcf4e871934d5f1c04cd634d9564d9f1f0edd3cb117479036e088bd4b11803149a2f603997989ef57ae0ecf5f45ca045e67f6c17d7ede9489cefbb72c8b1f098536c05d1f7dd4d039ce66c8970540e90efecfe5565157605629a4b07ae0ac23894f1cd7db36a68ff8771381806855cf9d8897c2f4baad19415c7bed36a25acce726b46a44ea9fbcadd6d6247b8007e4b684408afe766223709878f072e8e4723fada04aea67b4c9c4ac85711b02e2f920f4622cf39a394847859f742b6df7143a6375017a3aa0fa6364229fc086e931dbb339f6b27f8a524c72a1fac4643e3f47347cf60d3af6346f6e1be4ac37d208420f76fc267bcee55976e58aeab960d323268067d102eb27ac18ca78584fd0b75ebb8d18c9e7ce15bab16b4fc6af07d389d10f11fc0214bd1bfee965c3d3dc5c18adfb2b07acb176f56d0047fbf401378d3326742af716d37512199b3e20e4d4bf2a9036fbebaef08671174b7b32a61eee17c4a4014dae1c2b806219c84a43bbb3e689ea40589b9a049f600a987c9a7b1e52de8ae2ded62d042ce99401c48821c1ebe0deb31a8bdeecedece7f2f234b38028f23eedb9f0e62081b4785a5a07813b98126e42441ab38b9d40d1e1447b0c9d3ef1e80a94a16eed204104f9465b2d07f2f2064f545bf0006bd82b0768bb523a8186a402df97ca73520e9e7dd27967f00931ef9d2c66aa65f29f1278826a7bf2baa7b8a025b4c582c507ce788b315620366dbbb60f722840b95f49944b2139af020c8ec6799804182c032dc9e30b1c9a77e399448bf7b116c61717d3c7a629d606b6b260895dad064eb405aac4a6d76e773d5062ef4b5c4038657dbec3ab08b242e9d641b898062added5a84e8127f0ebb2b88dc56c1d82cc5961c62abd93c36e1c71ba5eec18f817bfbba41153ae7c2fa201a98fe4c2c8420ccc64b8b21cad6bf2fc1a0daec50de26bccb69b1f73cb26540d5f89f44e1866f38f2b9446d5ae4753be585bcbfaed35c9382b72d1a6b8360c56da25ee3687d67e1a96fba6935b43d38bfd4d2aa56e246cd4cea4dd01911819ba861ec02f141567c8b7fe645c3c5ce1fa0e642f2c7c8e378424d3ba79a7a90a488dc400da84f5a276dc6ac34d78e3be0426b7131aef44fe122267420e423c8ace9f8cca1a358a526a00fec444209df30e5832964b67e724a8c3746e1f41827723e797e78deac0f4bbfa8576faad01930b693808add63e017a6c8eb1bdd8439749b380fea823c0406b2bbb58ce31b254ea04104a7dc6af80b4a37f890c8ac754dd2e4d5a8966bc7c34271c194921431a39d6453bcb18bd33680c220411fcfd5ee75e31b56e1fa69b7b49e7c477c1b5fadd2ed51bfd07b4ffc40e044fb1abb5cf8254582305f51404b47b3de00bee12cc4af4b965de9a4bc672156276d5363e05e5ddd6cdf09a49c1abd7119a93a90504c81c64fe123f21185837ac0b1fe3a1fd6254ad2fe5fae8613aa4992d23a78e6818f69308aacd8bdb55b5698ee02ad81530f81ab4ef84a608e7b684164ab4637198e162e9dd757b3ee790527631b921f0d1651b2b3203752410afde055eb859b3bae5f932a99dec65a0b90eaede0f9eebc5f24139ebfcc818daaa456c4f7173ff6a1dfbcb871542f3e75f8d98b6276018def9ad338cc3b03a4e3884944e052b9657856ab79e95d3e8f71b5dd5ad89e249a12fde8d7a4d2dc0ca95c7eb4032e19b56b93e0b5966980f1ef0e408665e59a4bb7f7ef8463c7bd05e21737bc14c6cf4776371f0ebb950d073179f883b06f65f5c85a44079c1650cde42473b8cbd66fdb5a4478bcf45f52be0ed51f3150ed6643c59cbe03f0ae129ad0316450360aea50eae9b28ab27a98f9623c16526cd9ad213aab66077419399dd9c7acf5d5821272d3f464088a1988b1b421ff126611a0529ec01b603a0f38dff0702b4c9e5351f8bde5a7316371dcb4c80aadc38324c3e794e0df5e41d1ef46e8e0c6209c5fa10013f54517ffd5b1e99f3c1b2160ee3dcce6987d0270d27dbba73225c6565eb1690e4099eaa5049337f7ed52ea5c2d6c54e5cb57a5cec88acad253dd88fc3df365eb9a8138d7e3b19a6bb6959c25d6b7578d4bc0cb8030a4b80cddf40e1845d8984faf6a2a38428643041f968f11cd40378fc8e8001fde66df951b1f9e99efe73fe1d79ce4f5e15405f8d0ff8cc05bd5eb673d66ef7acf3ae430da16fc591b68240a45b36b9236539f900ed585477e26b308828603569bdac7547337b18075e03016ebe5ac16aec174379b5ca213e72f0ac55d989c0ee0fbade1027cd0bc71f34428e485aa97797d2553f01ddf0fb994f06e60606034fd8c183214434c6b2a8fb7bb4b9193389cbdb868917f183529debe013705a8ef86f6153376c4733d7ee651d60506d5eddc4926508a42dcbda8ca3b21ec393abc199124412fbdb28782df6897f4372fde803dea9f00ac1d69a8d0bbc36b4f42134af95531e8d8d23ece36fb39d43740a99c6b8424fb3e0a63cb5609e5f4db1203ecd5208e2d86fc99466573bd99160ffbfe8290e677ad489d5f3c2c4c8f200ecb2515e5213185b410f99ae8a3dc4d8bf4f1d2a40bbe6c7d230b6a966dbf769cbc34d2f98fab0e58288d263d3ad60d3282a1955aa3e2121c122eabf04fa2168f10b3c520c7bee4e5e04764bd18c5b43902bd1f2d9dbcd3329d54a0d68d5610662588a29c96d0a1e8fcb6d0a1da082b4f6af3babb3eb72e0dea3a9d79fd3772c19a55ee1e37c25aaef840db95c06653bdd0160a14136564f29f85bcc9554b2211dd1dd23871046f89492b33b50c053c377bd65b015f4f523bb5ac1a9c74775161c50e11b522b958c9fd550bcb007813a865dd4e352829b50d987b4c11ad135933017bc28cf9f4e7a13180be85512957af639f7c74c2c4f267e6e948a6baf6acb527105e89fb310091ba50dc1532702167dcd530f1747bdb0ceeb587d28b7d1892417c273b5c5b4db2e34c9f7735f1a43659e671d4988fb12b6426c386792a7747a0d217e519b1d18bbe49f7639d5c64aa2bb6e2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h70a210de0cde6f582b7f7a57486e8fcfc62a7666aa60a7f56d76d0ffe6eb1ea7e590ce2141014aad1ca2da6f98e543f9d8e2115e4ab26746397f32a3c930cf807bc87839daebd0a60295c320083afbee44a4afe6d7f10026afa9a96f5f06350c7a2dceab3906965e4b2ce8c17922b4e7ffd94bd6fc9356720c54f46f36f3eebc477a2c99646cbe43ec13044fcec822a31fafb10ba0d0bc33c393c54c99867a15fa48508980ed0fef9f2bf8fd77f16f8fd3429ead2fc668183c6bde3a54febc2adb926e24078b6d9253712d0eff25afb68e3774e81f5c518c18bbaeb09b82ef93f81384426edeac78a5a12a6aaf87396d0a46a439f9f4abb433c5967e5d5611dc9b007d01a0d9f24ea14caa4156f0b9cb88e67275755944edd314e182c120d9e2458b0c51c22bd4d5f035b435497afa456267654de3823a99ea71835f364a782f13df0ce63097a8fbd982e80287bb273fe0a69baf156f057db8562800c5f7402944c2159f01a186f20bad2d1bf963661e444159a9d1d1379c78c391d4630aed83980fc362b264d79e4c3af2840381398bad9187160c7a301d4fab5db83441815df69efa0666c4b16d0f958fd326331cf881857aa6cdbfa4262a875e5c21bcb79ecd561bfaa4372a04ddeeb377e288bb10f00587a79cb3746df723453997fd164e88696645faf2d76c73968e38eb8de6ad3060afc31ebffa346d1e2eb8f4927db9089a9e3d36ee1be4fa15e88be3a28df8b3ea4468b5e2c340ea70208a1a4e95c8d2ef730cf29c428f64fed9a37929fabfc4a65b61349aa9bd554174bdc930d9718024f0f9976cb5f893864b78357e60a6e53d2a673fc8ef4677daf3f68d613b713ea3bed39d0a6a084fe73eb30cc434224e34bfe91a51822df5343fe63a649d52b4a9b5f1851ab4e811a58cff591b1c3e73a3df0ec3b5ba1631c2f9e7b5c1099977679e3eafd7b2537f5574ea79adddea3feb6b37ce3d056f0dfe43e880dedcdfb67938acb7c3e8fb27929bd3cdb6d2f1e24a390b5b7680dde8cc463e2f9fe6d03cccdf5761a2712d03a750d50a8826cc202cea6f4e508ae06de584488b79fd105aa373f8d1c3e9307ed257f71dee9513adbd5d56ad44ccf28fad7cdb1556e1d97cf80ff33000b684b4e2c23bcec459e5723de82c7d37254013419e810d3e33da7e8dc559ad01c84101d0176b5ea0a8f18d2815a4bff4ff1e85e47367396dac2d02c67e265086a459719d7b669f68fef74e8b601a56a4321552cebdb69229f78069ac037b538b8a57ac746afad2dda19e676f24410f1f07a46dbfc508f3187fd90396584612a82d58cc3fd160acaad6dc094157a9c377d9f57a8ee00d94fc12aee01b9970aa6ce2c57af7d18ec8eae3579838dcf2c28903d7ff89d4c85da6fc5c72f6537cd18dfd5d17cd8653320c6c35ce42fc9bf1f582d17a76b49b9fbca5d61b18663f1289b403ab8e78dbdaca75a59518c536253f442d55062c758f6f35d53ba0e208d232879d128d071f180e532ef3b78f28dc52b25d27418fa2f2f6113cb02ef9a8d16b971c7211fd8698d585f870dfaa85b6834686a9fa49ede297ce851fc4841973e6850d174c3a63e1a3c13c1d5414740ac52c547da20c5bce4dd04cdbf53e0b80bd143260e5111629ebfc5b36c4b3f332fc6e47868e64837246bf01855f1713855d9bc4c367495ce13872ac3729bfa0fa1ac1ae30bb7ebec696c64b1b775c10f4dd0915ef3ab69cee189fc0dfbe55ed4a4b8116f4d3058d96c1b3731429e8722fdb4a9e35341b6499eecd43056f90abdf8fb1569879f523d42e9a445abe51e342ed908283d22bf6a0d3f5a3729809bbad6f8f81484a7a76ce4e14856730c0ae23650b0e881e7b57bdb51e27ff5363226d7721042396ff205b5cfc412f69f03576310136e3c8075f337bcf3e98ccb2ae816649a31b1a167cce821d4089cbeee6a1e3deed3af02dbd3dc94f7dea42a0ba61edb1516622baf0cd86329b125a0d2005469ef8fbbf86168ee4028d7946d38fc8bb5537a18676e15000edc1a070d189435b129aa7ce64634896d51e03515210b9f44680e03b09fc28f30806c3833f27e137e132cb5f116b1a667a74f9a115745474a274e8530718978bd7960d603809b75e1ebf8526c47ea7cca0356adea1bae45328e91968a789e54de9a6fd26f1786e390a74016f10b56e53d1380c1694924fe41b7fe430739afa00bccbecbb1bc3cbf3a0d89cde1e7b35099ed00dfc3d5d28677db482523990930be3f9979f8cd6fafe3ee748da9c0aa537a6411a8d42b4bd760cddf9b0448823d870d7998851b9eefbdae6483b12b3ef34ac69371a187f3c2629a8ea71cca36ebd9695b0a5d0230f621545ee5d6627bdc5a088e1a30d6483e54c616b9213e44cecc53b066bce97f6fb94c21568b591db29577df1e2a408d37cf0c1aa2057ed55db338d9b3fc6252e32b1a6b538567eb26fedd2d2f837a2c158f4f5b43ffafa7542b3161eb03abd63f17cc7e8b262637c06c777dc21b453f850ab659c6c561a0335596e5024effdace8681c269569d5cb25dbf6db5e5eec9de936f8fed2334e5dd64adca7a31704f4f22167af301ac24cf14553428fd85fd1ffe275d49e1be34a23deadc0aeffb8970b74965ff7f656d2e368f8bc756300ceb62a801aac808aee7caf4545a4d5cf0c60128f2a8b598b8886067d48778f3ec00d15d0dac1ee1c4d3dea2157b7d1385efb5e2341e2b02513503786a467ed7d2ca4bce0a1decc3d22403e66077f21d92fe627f79106fbcf936c4d14539ba1fd83d45dab4d9dcea7228bbb3399967f621c371c67b00844d2fb69b71b1781e78e9969c2eebdaacbe84107b1ac6533193e296f346e16f61fd23db39db5111c28a3ab385227feaef6d6113302ac4d20566a730189530ba544de3d7edd86ae4203e19a10b45ef647484490d7e48d1e07ec97a42cf98ebf76d70246b18a6b1ad36de75fdde1fd3c5d68f184e10397fdc13aa82ec8c2b8383c0f65e8576d5203034d4f8c6850dfd653bccfed3dadd47f97f49c404ded88f7837bb1ff2ec642fb3c86e4f33c86015326ea0b674d0a2e59e6282bb715019ac43f1d4de58e3b8962fe003a5b171b6179597f46b75661dc6537430ae270175303e97042239b908fcf0a89b7fb2dc226533ed5e33bef7340cafcffc3a525e8158b0859181023d722225e65a25c32630f6e31a67be158a63d8de3b39dd6ed7a2af977b2b316814383e137b6f0d3f4ec5ad748acff9818891ce8c55a8f8c48833dceec5ee54ef95abc6c3af72d04e505919a12611cadba7462c953b97937da589f35e3c276851ff629858ca4fea6aa9397248ba456893c86d24abd846dfa5382431dc3366001bbf86f13e0eb181642aaf5d47e845e6be49ad15767691a321a2b9b6257c1db5940c83081cbb20691811bf06cab791972541839c1f4778b9d83c900be099264efd87e9d38eaac786991f10f4b25102436b9d25ab4e0cef95e733069d7980c81bbf03e80d8354eaba848784b16b5e585dc215fb66655a86cd17ab688e987ed9561b2628a8ee742a4537ae3ecd0afcccf371148301ec409184940910f523e2b402dee599524bc5b8554415ed5733002b395c48baf52a2cd68defe454c1f9f8be1415e41a3ba4722357771d238f28cf46aea31c9a0d8cc881bb543658e88c369f09d3352ffc96f6997b960fa6fa570103fa5b3e65e6417dc464c433d517f3cee044aafb97723e5f924202ddf6a6bf90e7df5be79031071ad3e30acc256f9c557732fd69f1e045c4411e962bc15a7bb4952fdc423f99ffb507a1143322a708313791156e4ccb0e7b45f429418f0249cc4b2b232b8a88cd8e3787789463f087359716080614fba89af5d81608cee3dd7d1ab2004d053a810d8f14e0f38574bf870c2058a5dc9c1e69406e901567afaf6d6f0faa2c08bb06752e1a9cdb7c1edea66fee75a74b1801d42fd3d8d75a1a7a8d0a6999eceda1fec31d14184692c5ae802ebb38de4fb2150eb7a42650470aad97e5f99efead43ed64b61e652c90d871caf22ce0e6d7c716d5600766338b014073a06006de0652893cc104d09aaf1c748184de4482cc91ad2506571488658a5271a730ced85ed2d15c99016c8e17fa41cbe76c4538037267d114178ee4d3402b558151eb51a33a8f39595f480775ee17916cf4bbe19f13e92021d83855ca8adadd999e3046061d2b94a499854227a2378c4331d3de20d4633505757c3135c0fdcf02c77a0afa50391b6e690bfd5014e8e371136f09f093bac08b14c0879b6ec7cae1bfd48d5d800e2b161de42e5c06be33377f0d89e5363b875c49b8fc5c7071f91c5f29a9e0e85d28f19db5214a60dcad3986111827ddbc1e03a93e695bb8a12a12a29d5211c381f2108467938e3571df8c669e191c8af4555d263daefd59520e1906c764c727c63c1793f347cfeb0bf24e0986defd3ff2f79e7d663aa6c4bea0831704ccdf92fc4a76bf17297f9ee3f8f851054d2eaaf36267cef29924744cf47883fd30109d6d12f0d2a2b5a65d2017af177ff351d020398b7f71cb5ff8c8411a7e51315d7d9ef54116caaef9192d43285b1efcb557967cdb6a6f4f1f64fa00e07ec71c7cf640ae208d4c427067e12224701e89a1bbcd7b7fbc6d595ac55aa7ee4fd3bc4a94953c4af87d0eece1ffbfb0e7b2681ebd9748301baaff6cfd09c82eca4a14edc36f8379751ea6890bc5256cd2ec9926303af298e9bceebb95af4385df78272b06facdead26eb9ddb247571c4fa65923d9959d647bd183b92dc072bf53d4a279ee7915ef8965d074e6add7a11bf273f3d48710f111f60d8b36a170c357571abd706c6aa3fc924bb83e79cce90f02eb42125bf1c0ab37189a926aafc4c5870bde2e60291155299a21b30d4ea2ceffec5b392ad988c5ad8b95e7fd014df58ebbb92433c2174cc80efd569e570cc531a998d989f4847cde5ef4fb8cc0afba3f9c7bb739fd7ff8606f8f11a66f2b1b5f702f0e013e1df449a01d35324645b3603ac5f2b080c57769402e00ebb7bf5aedf188d90c3d62d44a53398418f28d20e3fba588fc889239751ff2a8cd30538b2ddba9b21508efc51cb6eac04de713b9b2eb5a955760c6eb4607a2b6bf6d3af8f1a4944057895d054e4dbeb43f9b32e936e5817464122daee6b7df1d149c3ba124c03673f0e958d75c1173a4dbe6ef186dc1aa24bea12691cbf13b039ee54735ff61464d0d731d5486e9cbda5714454ab1abbd2ff50e58e5343fafe3789ad4a76afed1859049ebbc67b99da11873745619a4005d9da64628ba718a6ce7d81f9866ecf1338d67f69cfbfafaa4958fe5f9fd16dab3fcce59857dcbabb8ef359333b9cac4e8caea4835d19d00367141c18ebd833e0281ab8516f9f691c6d75991047849afa3ef340771e8e731016b56fb4f0c34fa91ec78c3d184d585c4f727c73b2cda8cd63f5714263936e20e9c5746db9b06b1111c4dc21a93b7f02e101a8855c772eef76a67d133d56dafb40470a4a52b1465607c66ce582a6ea1867231f0254ebe29e25f5e19404347f5e79db5b7ae8741c6aa22b76a9b68688e810237804e3d46ed59a9e02caf0e2e4e0735e5083fdb071f35bb303c1915407f45a2925d207ab6782c0790dcb43b5d65d48711dfae8e5415bca57682cb98db82d976f83318fe17d3b35842af60740ad375dc93dc62eb34718f46c81786bba8ff7807d711c3fdc7cb035eb18f4388754756ffa26341f9114d54e182791032b24f31a565be17e0549aab686929b5b43f37440211904dad9c218;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hcd7c089228cc0c8f8129419b42052d9b6aa1bc2abdc6806d843ce05dec82cbc219b1696cc39766b80df9bd1ddfcd3d79af2cd66f16c76416f6af6d08a81b9b7423576c37082bf61de9a1963b6d9ce868a8f02044bc503e2ffd03aca09f90b115b58f2f7e9372f0339f8add2c8af30134f6848558190b65b556a7a8babcfcd0a7e6931c6072ed629557f9fd17bc65c061721103f8c26bb3a1b514c7c7363391045a6b99b760d82dc733017f8325812c36ada54c3fbca071a344bf1388ad78fd4f47677a72753928a7015065e64d5c42940a9056b0c8a1e8afc4773a81cbfc6854b1f0ab132f7d9c657bb2b3e7dd6d949c49692682ba163965cb4016225ab85490cbc0d666767508fd5c6566e4b22771725178bb70b34b9a5753fab73acefb53b5cea6be7f158f48b1cea7c85a6d60e9e2fdc0946cf6d97d3a9428beac8348d53c91405695683c992cee4ecc06c2e88db0fab7da003c9c7589d8010d083e36b74d8ed9d5ce7e9b2ebe7e2863d89e444742e24d33b75f864d74543daf725e784f3d2c2380e3641678d9ff7c587c8a61090834e7b7a4c0349b6e97cebb47393171c06c38cbee9170bab8c63916e6e77a6a040ef3b13e6e4b21d7c65aa5b26b138d8d981312258a69ce81b2c20fea12c12f923b268cb73e0525d54859ddb83cea38e66ed35d604712140b75fa30e73905014c9e51e2a7ced1b61f6a8b036216f21bcda2215bb5c8b4ac8849d4e1f01f3012f93cae40897b85d8e8468a0c78a8f81176cb82e1667f2b4c49aa97bcb577f043d07a0c176bfe2c574ef67c7bbab0f647cdf787324036932b1a5fd76817ddd1e0a9dbc3798639fba0b40fcbb732062261b9701e488bd1ed641400e87c816cd4dc97fec0a706e59c329f5c2da918a8b58438e4f225a1720b2704d6512c61d8a1c374796828cb6377c3e17e3c9a2452016c3d05610668b2ae267762594eee732cdfe98c710294fd33b2b3ed5e1c1efff2312abc31f7c9a838b3486f8007b29d83e95530b29314b21e4016ca7dfe0096d3bed1821f46f1860716a24f35176a06fba4f216014614c8bb96e690a5c81c3e4dc5c2158e95a3c5bad1932460d59aa997d24f9c57cd0b251f2c4b5800e822b34742d55bede10a014906f525a2efe7fd66cc0ed206f9b12b90688d7cfdb08bcd98be9444ec234c1168751ebe8010f2691b8a7d9ebfdcc2b101322469653a29340d03a42e8f8af699b4dd951cae836db5e3edbc0421e1cf5af5888af18ce963d4baea63dec3f1f1e625aba05fbcfdf31b39362ca0c5c2fc83dd4613fffcfea7476cfd0179f630798a10d5c840392a957c0ed5a159bd262db553d5c7058ca1d460138c475627ca6cfb608edc3c02fd1892433609b520a090d999400cb9435724120663e33a4f5af471eb8869f6030ce10cf9f2cdd02fab4ebe26b9a506713aad29b5f4a97e5c52ffea34b611a67ce665a55be61577fe0ea3b6a9f0977640e8102248f902a4a254aefe13aad01ebe13dd8a49a51d695db91b39c504512577613d34c77ffa127177f751c3a379d5027573700388f0fa71b7d39b242bc9cb5c6d63943c9f42582047caec47ebea2a660a7c69f9601c60292e4a5f9d2d53474ebda5723bb16bfddff841aebba60b5db661bab97112bbedbf705b710760e3e7e750ccaaeea1f0c79c89e93b373a16e84628b4b002d7fbf2f6a37edf648223b7bf00a2352d59a84f664b9d4de95bf34c8ceeea89918309c31f33b82e37159ff2b7a2baf194b0032407021fcfd52e890fff960ebfe258df2736ae525d7facbd878ff79c15afcbc4bdfbf040026a48825272366f3d4743e30ae7fb6f494b34226e71524fdfa1f339c1bb074f29c785db670d16ec4fc6f1820de0b002af02270744840e55b4ab96d5f3f596112365417c54c6570c7badbc87dea72a388b824f173013af64a85533c0241c54fdb3e827a38b86fad4d4306618f76f834e4e7843dbbff2fa72df21a6710685619399460e76a4515bcef52e6944b764933d24f0c399a2306c3a5377061b97ad225bb05d273413270d5a515f1588329b87278beae418123a25ea710b4a6e89ada0c038e9ff94f5e3c17a45fae2fce81d4db9839bc1c5c3505bce07e514124c7c117c9458d1b1b960f5ed0bd63f437f310632becc2f3cf68f4096838beb5189280f9a2e0d19b08fb3adc96b7d1f9d4c2442f69f373d358c08082efc2617dec1866e0087fa06c5880077ed34f49c03ce6cea27e1df6d1bcf0388219b5ad91defd0e45441fecec5e164daaa440c721635d19afdaac3d80bd50bd88254452b80987ec7b48588e36f827a4621c9477d893ccbcfa5d30e7a28edb3af806dc1369085fb618bad5c036ad86a5528270f47f1cb7be26405643d189453cb84c0d2f86fb9b4134a9e4e93fd9f28e69251ed38e76d684e4feec45073f76a03054c26850d385437a731439c38f745ec56c1fae1153492f250ffecfc67e2c65bf3b0e3509a6072d402d8cf1bd213cb0473b6f1c248d7126f77c1ae2aa5bc23d68a864daec9c4c7e51e97794d8ce56135e90b25a31922e3d2dcccfe67f936358db422ee6b5a86716e81965d79cf6bd4f31603ec390e92f2bce0ee55d23eed39b8abc4aa27ad25029112f6c540701af714e270a79c657e11e0f74d392d3e0585cab44cd79795ba9a507da490ea89d954064983712806f747e5be90f9722cb0149621ccf29b7ae03633b3a7dd3bc1afe01d8aba519087eafded0f428c8a1317f1617eeb233696d1bcff100512fef15b692737736b00c09db6339b7978f69ba7b56e7e0e76568f3ac100022ff223123e8beda84e07813bcb2c530742bfbb966d5384b5446564974ca6e0c5dad1d37b5e1794573328be4d41ddd8d76fcfcfb4664878c579bf68a866ad1f8f5ffdbb5d202acba606cc9509aa9f1ae87a623d0526471d193e674a3ab686287a92c747aac4c47e42a3347478fee82143063632c6f31f70be03b7c29ce762ace7e22b16fbdff697d8e69b6a7289fc7dea7c18fed7cbaff82fcbd3185c7bea76b0830949a87696168f6bc97b83a5b2552c6cfff510b6374adbd9121c219d1a144cebbf8517cd36d9faa2419d468a60840ee8285761b842053e6ba9acb7db272ef8c14b0fea958c776c65dd7bb8951294bca52817b48bf9f0762c05f0a5829ccf1e776c59de593c0b6074335166d4b3b9072bd5bba135326ffa689cfe1a1ffb95e16e86f5711962434b70c3c06b359cebe4defee796abce09eba503c4a801e6a91a4efd61b054bf46393eda686f902dab60fba1f8eaf1606aae5acf66b56e45aed0ae53744e5b60b0183c25641e0500240c4fb15a1c1185c10ea54e3d050585442af267d06a7c0c2e824468ca6eacb6dfc02faf7354cc0222522a0798b17e81481f9e6fa25f225af52645d422238852adcfec4e8fb6ae4bdfeffa93920c4b9042d6bcd195eeb07f0ffae966314fabcf3bdf8c483dc0bbf85070322ee4a7ddcaebdea8b053481e77ab65bab9d18e475c88b6d30fc669c579eb2b4e54aecb5da73e0ac36c8f30ed22e25ed0319bafaada5395032276751ebb6a5cafeea12d7dbe48d031b7129efb7fd3a51c6bd4c736105013173de700aa8ba565b57559b8441fca8a1e5a69f7eb31d53a5e86d7958176f264100678e79843f93085244f86cc536dd2a08970f587c82901d71d632f6cb33e01c1c858eda4622bdc8a84973d2ea7c05e3a33d63767b1b78ee56c6f90d88c91cb4c9f5d1913b28c0be7168a818c83375acc7a22d808faaad38a1c103c3896b5e55583d43c4be31cbc1f6322efc340888f7f3d1f39c921beb55de1124b66c3cebb87e374b7dc9daaa8450c014af920e4af7c850bde13c22a9288ceca5a77660d668755a07b18f406efb2540ee5213787f63df9add3d0ea97271398ad2ce1934d61ada6fdc511e32837a3b06d373f333a6fe40e2c11278ea61e8b71a6228022d9196bfa74327ebdcf7360ef17ead5bc0ec424b6ba30ad52f46e9a1fdf834a1641e52b2b55b02e66e0fb02a9d9958ddd0d7901eb3f9b6808bcc8eea8d8af602138dff94f3b992664adb866514ea76b5a43d1485ba1a301d207f26c43cc1a3bbe17f9e4eb6294018ac224daa9231e760adc3f546f0a562eb63870ba2cc5718f564894d1fb8efd6208a17931428ad954541f93deafe063e04009871ade79f2c4bf17605db5ed02ecc6eef00435891fda22792f29db4add172db3cd790d5ec51ea6b60979681e94c11ba10388785efb95f7c76dc09f01f54382b067ca118b5f526acd7ada76626feba767cdca802c800c94d2321ef854dbff4bead0e5bd2575493dac9323260fccdc9a89d1bc4d74558b0c8042001d7c0423a532e6a0d0848f4a1001c55d43178da812be9e70599771779ffc57466cd9720aa20795a1b16c75d7a7322b68656259603c686fad3720619d1569a4de50b80f9c07eb60b13d31512cccbb9ab5bdf8ceb136266cf5311b5063d5deb481bb5555e05be983f09143a2750862fc4644f264ddd94ebd2becce4837ef38f727c8deb213f0321646437bc2718b3c97dd5bdbe0dfde75d151ceed2f814a1ca81f9db8ed8ea0e069d303fb3b78296f7072ab9cba0c5ad1c311154b206760bad7654cf8470e9294515c4df10bed7fc39b0480ddb8f1f73a44e28d67f820001de5fe55ec0f5c010410a0a7cd523e16e3334b54b56d062e48e084e69c126f5654a679f32d61c2072ff2fb737a429a0e9be5c76758e8ceda0d7b98ffb9ef5014fe0144aec7a904f231b02487ac08b8dfc1957f2a547d181c3a6d8568fff9e3b702e559ffb14acd106a60a14b120a210341a1e657039511a8b718c6a06fcb97f0eb5d48898442e04b0a0e3f8a03e9014280537895d6c95b810259f33fc90f4e831d5d4fd88035b781d778f8b254dc432153b9a41b053585599638e2a4b8d3a740c9282e123662db48f27c6d4cf6554177b979aa0d989e441e517856126be0bc69d251fa5dbd10c94247402b4b5544f89b33308a348766bb3834274cee48820b09a386dcdc9e4a5de58fc0d4cae09de1f9c049d3443f4ca8594a9434eafc8b82acafb30f55df405e30902f4e3ac81f79ca68b9d912daa108e86a041656610c0e1d8b227b55159140a297421c19e69a84e3ab8a52d1a60f69da0fe4277a2647d963a78c585595137f92a4bba06626b658197e6647e94cb5d4aae64960abea5c2b2b1f9d1f9eaeba50ea9a2d3c6365eefcfc3fb5a7d3741e8d9108691aba818e9f2211f071203c78aed0d56718dd658a1465d23b17c5128aacea0eb15e2228d7f345a53b93896acc467ac0fd9fe4a51ee197c1347d25ac54181a5636dbaf6828fd2f6857b81b4a256f952fce63b1ef68fc3c820c2dde0c2060f68c92177127926b2b57fcb1ea1e593c2776ec8b230a67fe138378b3406bb3bebcd11ce84c168d22b709b12d8b0431733147f9314b570a576c61997ec95740309f14b8ae2f09c9e7645bff84fc2907c177bbd77a14417f8cb890f0cf4c1e43b044e15cd4c332f5b158495c657ecbfc260075f397b6393ae4a945f1059a5fbe26fe0021d241adcd82f7f4f15c5917c3494648a3179a0adabb43008268daf10b150180880904eaffec9f91b2ba011efaf976486f67b83be128ba9c8458e27216a3364068e1a0eb020e8fee4802dfad05c1028bc5323334205ec3ecd913c083bc64db9b9a2f0de75c60ede616176557b6f236039461405be5a0089738739b93e42c8ecbefbb68ce4bb0c06916d80ed89e0b845ff663a1503f2f0a785d3e940d304e4807a927206a4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h2c147943e43ee27bd4fd8ad775f128b3fceaf4541c12f313e8efbdd96a76b473c368df2b852349a6d3ab4c6c97caa28c1b985c64085988b0d6c58d8f2b833ae976f99974d2312adf2b769775d91805ec77f69f9fa9e20af356d2b0c55937e929833c0e5e95a91aa0504cd4de9fdeb8c6059333efd2234a9abb7bbd0c895c2b886371b2461994367bc46d0e27041991450942a8d878a1fbbb2346d5f8f030f6eef8fa5fbb7eb3eb3c3a597d014d0b15eb47f087016f874e1ad318a1f9c8bd9747369d869c6ded2072c1428e744542e7dbbc27074d7e250a4773c60ca5fb9b2c82e43844693192449444b52ab7b50536930d656b1ba0fc5e02b538fdbeb73160bae790ab98a949e0d637fdbf26fb5e5729a9f9dca928121113ffeadb90ecd4dddd8abe14bde0b956c7fb00476af5ea159f2a85e8874f4056d53a24311c3e85641db7cb21b7dbc4906c1dd2119248a8025873df2d75c4ca56e19f4c11077cae40469cf51850ec540ec58136bdb5ab2a43eaf4351a5ff8e514a4464521e933c75e1d78456096f65e6d1fdcb783b1a34140b30c94b6cfc806d0d757832242527c172ef49b1614289a18e07f5158edaadbe0691ebf4a5971ce226ca05e8f0c37150a7d209d627fef1e292d01d8d9e0f15c9c2a2ee7b4c8cd2424815903edd8b13189cc6db543fdc5cb0e57987c0c6ee12a540a3c2a92cb92ced3418177b88fe549cf7a723e28b5bb93a81fe122046d6125ded683886530a4fbd20114a25b2c9f2a3641fd1af8c0da497a4a9bcbdccd8fa9932de62f87721be9fd5d94928ec42d2f62cf7bd2d836e32eeab7b22f4a997ab829a861223c778ae706e233f4f35f28066f2388bcea2cd899e901a4b1be023478fe7f1ed678c26ac1bcf743d4ab36045772b32719985da4f4f5657e03b2bec8d40fe066ddafd63b140bd3d51c123fe45656f605b9e84b204675c892416640203173fb59fcb45d7de8f308469ce772e74b6268988b7f3c30ae5cd1916c44b34d6c8c507cd2dbdb02e0e4d08e010910549e7cea84be6ec76b880b13ce2c3134a4c4adb677e02027d2be7f452b27498bc9018b92799e8ee71c84939bd391ef3608c2fe3e2b02a2cf27d2e15c623f8b75a157118c390f615b6cf2aecd7d4a79a8110461a5adc943ec7a7277e78c94dc0d9ce62d3171293cd24ab0ec72f68250319dadce531283c066b2fd74e9616a2d778a56140aa1ecca524e805f5c3449a717a43d5282f49f9d1840829f06d778748ce19ef79102e62e0c0773f754c02af6b08d1187835420df4fbff1317f80b3132e62e6ab539c48b427367debbe7031db773025d192c30ef09408f5a67dd9d5c170d25fe94c6f6a8ce9f0c69b3794bc766e04cf202169111af33cb633233c2f266df49596251eb404317053d2fb669298e34b01f2f8368eb2e3216c55dd3be9f8aec1029bc9adc1be0fdbb24b9ebbd8a08f3c68527b6a4849234abfcd0a2dc7445371fe46fe716cd35bdd3f4a9eb549ebfea4a400b68fb9321b872ede349e8f420407c2fb1ffe2fd85fc4dab0957a95bbb22a2d82c6f3626f40211e756f85838d53407582ab5b970d761f75f6698a5e0b7bdafdbb8642fb1715cd1f140e4f53400d027491ff7daec72fa98b95e7b02a8eb9a960806be8d53d95d8f0373f3400b4e8040b5caa2ec50e0935462f677d597237d96b811e7353dfa3e36b39ad8f6be0a04da64f2376c91d87e4210a7a904666bd807f0fe1380b3045368dd7e4cf5e13c9c309a5d7aafa62f6ce39d89d9b75829d59162c5f044d58719e48315a5ec9db942da67fa348461a89e4d118ba351d9823ddc39be0b1ce680dad6c418e5472d4cb11fb8025f13d70ef80e9ce0a7affd6d0df04447cd993eb2e52cad55742c0314411287af5577f4fac7a79aebd9aeddbf399d8fcbe1ca92c6166dbdef14b79447af206aefdf5087489d95046b0cdcf57890c1ac53b6f93a688860ece95743fa946645aa198621fe4393fd4e3e7b181c3fdbf8c31f5bf329d14ff0369a8e4eaa2bde350fe8108df43be01b6594f0c4469aecfd20a35b4b960294e9af6c4d38d1a33c6811ca75ef488875fe3102117e4edcf0a40f682daff274c5b6310d05c8242f7790e54c8b2c14767cb49936f312bf6976812a375bd6caa38f903981ced4332feeeb8a218e08fc0d3ed68668f52e0339fb00317731ea3ca620b4c634a59affc52fe5f1a20af18f7f4c51cc2cc0983a1f5f2562a921e1900600340034cf917fa19dce35f1aa3bfcbaaf66c40ad354974a22b29abe581512bd1fdc18f62f9e3cd64e2cd751312e5a7dfe9d9b3564a178d4c5127ce061ea22c3f735b17766750078118422f3155a9d1bfc8d115f4e9ecce3600aa45a5a51cb607f36143ea8493fea770d3855387d6c5e74ed08d535f2ebc81e97cbb6a6a486ea9a3e74cb0faf814f9b2d468757778de66205c59a5a0001c4a1de0f9c09a1f424ca48f8943b951db7f973cb50b5f5a92d73be02092bb07f8a6c13f71bc995b2dd5071ab88154b98446dd38292974c98b0514334a45bc0b1b395a379374c7ac6e0f7a905347f11c48f2c1d78d2a57c5244155b2eb20c70b1e71c93cdc773b1ea53c5adba9da71e387173ba603baf5b4d2726690f210e5b011b2036f188a21a06ccb3b6a4c6259b716f5732d9a641494947443264780c374d267de8450ae156a736c7bc9a0304f528fd61c8a3129148d9117602d962830aecaec71bcffd7181b8d23bc34336320e72d45bc095404b0a0220b73a88c532f89c530a699f24c32a2f8af24cfbb25a085f43326f0c2dfb3b9971d09fa41b86eaad01ca0ba264bdae676eeec5b240d9ec6293d5b60ea3f7ce4f128b5b6c8f06b3332d68dd530409e73649866ed3296ee2737f5b15763efe010ab209fd3ff43ce2734c889a3ad6893d4d15e05627ac00c2d2381548310fb84170cb5ab2c9d768c2b3ab800d5c26d0588b7ff330b825fbd92239e14c19fa5a4ebda36782aa94af6b0f8a6bea4bd5c89f0c77e729f9eed7395e4853fb7ef85cd8c8be007749c4dba1db1d5028dd567ceb61be6bd11d113e7b32453a785276899d7734bb0b4e8d2c65a30f5ea2f2bcf82e2a4949dc9b1971d6c5dcea2c985574531677ab1d5e995dd814b89ae5ad418b02d49e0e36a64645db78ab1e884146ca5e6fa06093e8bfa0dc6b28723bdcec681ae41e23c00144f1185ec6d6807fc316cad30a2162a00e21b8db1e6d96c8120042b2d05225415c096aae8da38b1cdf44bc569db635dafaa2c51ea4536ad3bd8f4f6b859c807ca18b61db2eb0ca207bd59862eccfa62690ea7a51fd3f6e6cef2cd972814a837b8f6bd433cb59599773f1673c57673740f6d9b217db8ae6ece949920c97c5245868560b7efba69fbb39d819972f164b48579ee9f3585f341753a1f272655416c25369f9421b4a334a920fe9546caa2840ca47c47c15ff33356b9395f42aa228c367eaba01957b74461ec9334241396b453c6391773c53b129fa9e50c13d6df0481a9766fb018ffcf93f117ae940cb910e481c8eb15b3c638408609758d0a16d685b2bf898e5a7aa410fc87402ab1c7ab4ae74a8009d7dee08398fbe214d2d1a9510973a5f1eba0f2d89f0004dd48e4a3d8e5bb32d3d528e43a7c29b9bcd2a9db04d8255b35031b14d1848851a981157c97daa9de193c9d3117489b39191424e774f88a4f8fdf047ef67be2e1b7f59749fde0ab8e16b3add54267318f2956b58f94128e5f12991945ef76aab101e7f1e74c28a066e40525f5a0cbd0fffbe0d53be7e40f8ef89c327278f13c09acb2ec42d61b5e6979788560c52ea7ecec41ba570dd4b051b017c3b58a51a0ef0e1f8e252a3c3f72144b8b03f0015c4db26054923acea934d7d4c0a9e826297db0172225b53da3af9a4614bccb4315341313b1e69bd2aac734228b4e116cc2aff1972f8dc0cb715ab37b71d86b3c5a46acf19c3b3e5270013d3362d664c31d81ecd477ccc6a23390043cceec0a07db3d116b129a9fbaba5b714de1b7a211bc4444f41e1a4274e946114eeadd6615820186991a6ad7f7c7ad36fb1c2853375426cee59c7f528d89a0a2132f893a125ca65ad65320567eb519607b6ff0a1e2afac5fe090d8921cbed952616892b5b6ce5a934e831636342d666d2ba50cbbf1f48e6fe0f1925047e344ef70549da52e03695ccfaf1c26add404ae67f82049c09c2dea99fd335682f14066d0f9fddcf2c6ae6fb28c9569b6b5b74c1495ef3a30fb439604d1194acf3086ae90c2333482218cac1cafd96428140ba0793a3731825c992c8bffcdbbdb6bcfb55c3eb4b1c30f25b061f9bcbc0e9795940093e3f2ca516d9845dff6edc9cec4a7137a6c73f31ab3722683b00753a8d16e4bde7ea77b78faeab6804630742e99b5b96c8ef4332d5a8538f0f881803afaa63d4809afd2881bf0b0ca4988dc7bef59a26857ef389a19b44f3987d487d9addc87574eaa0504504eeba10ee2db21a75cbe2b98fd74decff9ce64736d5b2d9d666133122e34b32061368fa21b0f81f86bd174a1c4b684a7c6a78781d601acc0a42b31e504b657660394b0c7c69dd4ccb10524e9b9d5e6b59c528a7d0a88c300b0fe05b320f3b499a3c10985ab20335e424c2e9e01f62bb5ca0b9aa1c6814e9646116fa80d224c9c39a09b3f733b5cd9c8e236f76c121f50724194bbe29b42aa2e2e6cd78775f238fab7a738a03f906e8fbc9d688ddf092e08f6e261ae842b9f3396a92ed4ec4f7c66215ce473bdc94ee50b60673c281f16a466eabbde0a0087bebb3c38720480831a79191eaa67e6fe88c99e21b2abb1cec194a459f90bb0e4ae9878106d9fd66b17bc882641a6e788448b7f45855816ab2b8665e9728ab27b4794f00d4046acaaee73eb9703855979bcd8928653039defa6c588b875708bcc0b87ab61936c7f9f375505f51ce5168cc7561d97def3079120016c6a18f46ac5e93eae0c858c7f02437dd2ace096c2453a3980972158a83d0b03acb2ec09c239cba95947b6961d69c677569125c333abeef0863665b2ce81d02a6b1eb784088bda02b63cac7ff0ce2c499de15be1ea137606bdff8a00e3dec417827419c18ef1fee44321c0165c2dc2ea5ae652ba2975c9560f9802452ff78aa684b83e60ea61b5def71ed34fdcf08960374f140443473c2235959180bb6844bcdc8cfa0893bdd5c8be9223f67ca07e6d563e49e53d6aa1b430765dd9debf28d8f40f8ce54eca0221e76cbf48c8108df7ad562b8a143853a0fe144b493fd5696e67888bedb34d98cf81b7937584a49c8abf0a086d7afe70f5dced907fe9db2c895d265ffbe310fa96b929a6602e51e25155281348de5c398eae4680b4e03c62488d6ffba74f875004a056075a4aa03d8c04081a32e29305661c2a011739f1d2dadd4da6d1f3456bc2547814b9a1e121ad036d4fd5efda9eff28700878fdd72c68c10d3c49b8ee9d488a5a0ce58c7cf1c9416fab16510ba84a7a7053f4003873658694174c0e2f88260f0ebccb9366843587588ede3b3d76ba95d9806d66be852579c517d2f715361b26f6cd2ad26700ad5dd7a7fdc8a52572dffd30d1d21d9484fc8625e142016c7d1d94420fa02b90d03d87ba36f02e3a805e3977aea699f88b7918ed538c1de0c74b5b8cbf661db8c5a16c64a9dd69699bd50dd5cd564c7b6737831ea5e2f64fcc930e635b95d54c361996cf105a1acf9f5dfa04025b4217dfa021422dd3b55490c7791373fdd8f45990c676cbff03c8c8a17afc045e03c8f70131676d8f2df40f9424ab80;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd9890c690f288f3fb8be1df8e70723b469e3dc941b4c039d3cc5036ae8b27a0bca625cb92c37ceb1ef9d7662af25982658134db6a48bc18e5dace6f4e5b68812e3ff4eb6a1ac50193b4c33d6bbed08660ef3f623d311124311c3d5e380fa37ea4f6ba8438b4e1947d4ab3a7336238c3701b8e4ae680b95c03af779db5710b0a9499738a290fc356c72ed3099433c3af123c68076e3a7e868ba4abcffcc2ce28d483db53df9fd743c1e7b27705ceb6a2bf6e389e7400bab81c9f7a21f67991ad63d34b550bb7290cf58f78f0836c576013bd88f0daf0a8736f5671f53565d86e130a2362861ecfed67db172b52fbc55097689e851b93dafaf76730b984b6e8456306da5dc48acb956fd0a22d009002cd111416d331be142be7d9f12ef5c674d6a05eb194ccb4f073bfbd8e3efcdd12c74a97ee760de8ec763c2286b10d75c7d4e8142f6f19727cc9f5a48310f93a9975af19877391b0af66d21b3852ad9109e4e6f686e1f0b894e915fd050e25f3e517fc2af289f7098a60003e8a700102390605a2138d97d493ce0e7d8b5f0dbe6222c4836a5ae7f47236da3731e94f6fd72f7cf8ed6959ac68737a742e47ab27a936468f0b0de2926ea458336c5410de971e9ee39a78386c4e51758f38d18291b4a199eff7974a0c5b4fa8e3b31430202a38fc67a90a0ad230a9d262ec7321aa4dc111801248f70d6f98590c2e521673b9375c8e6764809c0cc23e151afa45c12bc5e13f48ee37bf6fca7da830394c314a1d6548250a6dc8b39de02678166ac49f383eeb81668c34bfeb188dd2c94d022b72238613d8c17a0c143802636b4ee140110b806e1baa75c6b25654ad47c75e711ec95022cca3c8e62162f7801affc87e035c915fb5582074e3d60c8fa66bd0c576595e7e3c683e5b4e051530ce871736c6af52fe81baa6ff636ed5880cb6067387db82b4746f8889249f8a5cccafdaef93842b72ee4ca86a8b536e271057bf48ac322496f2bb8c70f3d99503d4687f8e977a8ef308ffcf66cfde68e0c2a6221a3a3f91d5192659f0fb568d54ab6ea3be25234c516a0ec2819bca782b14fb1b4b7a3e92198e46b15c4dd6b880cf5eda27fb5a4c97df71b7eebcc8acadfa745319d4ab10b1599e2f1ac43f62232741f9d77f40c9b8438bd80afd04de8a80c7d78d08f27eaf43a4debad3e403a55e7cae98fc56b60ecad3b5fcd29c9e3472ec75333959774b824069b6b206ed62cc6b30a03a5a75ad8655119189a8fde6a222534cadd275b524e265104e4052fa0f3d6add402ac0b939b6a138407fcbf5ebbbc9250a9d36fc81b535b42950119bd2a5f3141e93ab420b1dc31d02387be2dbc29049a162be7359f3bacf4ac605a89b3622fcb7afa906b91d0bc5efe616ecc8e8f73b6ae0a9e96ae21c284d44ea46bc9aef600c04d5260e07815805ca1cfbf5f7c4c6e0a80366349288e46f175218fee1e91eae3c83002afc71e7338ecf1d5c87655c3fca29de52277c0a0464e59e3c4e011f69a6270a35e993bb0e17ee5b6e4ce9d4c470d4661152c7d0d392fbbea6e10a68c423747fe91d6a685f24f1f120e074f31a8d01c5ada6362ce7a0ad49cdab98f28f6140f4a0a505b2e84f46254ef0b29225d511e24c24851b863128a3a3c2badb60b5527fcef4aeae6057e5e835e0784b341828a3fb89b5423aba52b43ee8034ef979560967cd43602fbf01c3b0f8f3f13caeaa62e2b50290fc9cc95de027d667acbc2ba58042ecf3e98f56a3716e6fa089314c8d7c8b36592eea9aefd691aa6f2055d05540b80941d3bf0f5c681b26ad499261e1c97ba4322634c9213714c79ca89d2cbf0fbbfc13209120fa09da837aae3d71580477f33999fdc8ecf70fa04de947675c731c540d713699457aa2f2499b9df3bcafa888432438604febd454d6625a5529a2df4da54f147a94fdbb3bfcfd5248706e727cd97ae873907cd989deb16f16a22c59839d607a602d52db33d31556a6fbb3048145893f2bf51b588f37458f29300ea171eaccc752aaf885e0b00d165a6308e9a117c711fffe3383f2240142408bee691fce99a275b1a33eebd2330286a9cb5f9e82c94a2fbca2093b82adf626f1a75ca2894136aa32175968ef7c6f70ffde58bdaef4918f022f2e1d2b99b04ee0cd7f5cc85d51daf197981ecfd0f012cda593c58eae649a312f1c6e5d109e7ebde02438e3c3e28971554f4a2a12ff3d1b1f4d21b786a41c87429ca74ab363e6ad21258a40b63f30eb09ce16073a8ca8975ad60f910f6e294df2599caf296e6d25812eb9e30da94e1e6da646c54607cf731144513acfcdc11b01f4adc047563b776dfbb017cb94512632df1c3a97a1f061d9787afa3fa8ee8d8b0989ef22796dd176303ec7735f5a19311b367b420b213135c5e7d1c7bb20a4eb84a7ed9edaa56e268103641fdb77f30e0f326728ee6b2a00a511e1c73958705534deafe4e89558b93d4e79901c62e5f17824176803942122179bcd0820deda8aa977f5b3f5f88284ce781fb520241d8a9b688b5ff587907897a20dafc6903f24daf56e3f87cf421054d514ed022f65ed21ea4d6a51bec04d1f2ab2f522453a613cde38b351f6277dbd36c1304293ab6a6ea5d73eb5d4662671fc2c7bbf1318b1f1eed470d7dda004b619841c8ae05ae3c17085518929c38bd8d5de2260b0d447971f7f4ee1c51862715c690a8d32f5bb535ada642a4f34308c5097cb76b128c9f026c75cca709f0e3ab3ffa9634546a57881e836c4fba4eea8b107bccd7a2bad73dadf0f9089a1dd7e26725375ff388aa1acfdf38f053ca7ad20eef1b818906c48735bfaceccbf8f34b2d97a60e3dcae0b0c38b6a399ba8c801b79acc83e44ee7a70ab4b72f0c8afa7f7c5b4f2fe63557db7eec172441572d6d788ed1ac99b5f1f660b8aefea7d327c27b6974f00087d1f3d54ff32ccb7d554d100469c6d3adf20eb3ad66d5b21fe59ad3a866e764f4c63468c2c1dc9de91d5d6e9f7c52539c8b04a7e53ce7044027be1bc0ab1a03071558d7d659d8001d6b777b2c437d965ae605173508d7db6aabd331d377b8337831b232b11c3126a397d1d3349fb22e0c5b931db85ced1d1e96a931e87c83b79f47180343f215898fb29751ff8ac940d9d90adf4e1bd49f70af02e88709458a6c8133989098e8df15abda950f3e01e39316fcd876e5f39b93ec1233cfe02b5a7c66e99be1f49484b86e16444b96c0d2d79e006337c815af2fb97f3b627a1b5b03505d89e31e6f20f2ee8026a64e6801e4b60ccfe9f405ae68311123ef05373e3fd667c3a175d1a1831605b04350770eaed9f138697e01ca2a27d2ead0fb0ba3d3f455823d5d05f9333437d34b8aed531a3ea58e7e8f03c9554841dad574fda1b5a4c0e7286f8b546a40f894b537d1593696f57b52e8a1a695ee85e17155744fdbb6669223c4180c45142fffd977456e3ca9d21abd49c33cabae44e69d2e5a0cbaabc9c43fe7ef19125edab46fee1f0007c572b549e9b41b1a678584263eeea8d344ef0b2e0775c97e380488689923d09e36f5f4cdac4479680267c7d6d22dfd3a6895213653489006778667de4c0c1fc4fe61588d0ec964345f8abb8e0d4ea6889cc389c313759e84688db45cc58e2b8f1a2b0bc10b6761f6c4bec4265efcd850df9c6be653ae8ff8716f2d394a90e9790f6dc60a5138ca762d5125b032f4d81921e2fe542d55f8a61f6e5e9f2db9760edad1db10b9bcd7762e94fe2189c96dc2e092645fc1200c8993f482f3b15045f40873d4d3190aee91a7f1b63377da35436cc246267dd0ac7d8d102b5f442fbf658f2e1fe806ba566055d133751c5e2df72b81fe48558eb7d0e582f926ba6158e7744115da0c01e783b32104e035588cb6164446985fb198f2d02bda12bff22663abb549d955079aefdf89d4c11867dd484a5eb710f55147d1c95633abd362d62024d20e976569379048c59e68547f0e8d2d8dbbf6086e90834f9d1cb0aab20cc468bb51cb23f764a8f2d1fbc00e5b14e0d52511e296c727f5292443961360180b0d872952a40ecc0c4d165cb917eabbabd4779730e874ffa94882ad78d4a99a63e3bbea89e1574c5e3de3d8a0d3acbabd0ba092c1e26758c50342b82efd699a2c9e543d95b975321f3cecf859701521759735a0438df2c6888e4a56f740c2d905f84c927a54f859910c135eee65218869e8f7930d682ce83faeaf5ae6b695e8f8d1acccc498570f6567b02f38052d5a8607750dcbfb074b7c697e64196f8ccbeb90ea67c9031a6da8e1a780b762c0a20b805a0e5837ccdc3a95893ca0fa98d2a34eff55eff5090e7bdb1b4594588e8250c8e84660da84ac0f33a03d6847849508a688fda011e9e7ef50570766f03a37e6282dd6992d782c8638806c7527cba4d1f68aa66a61fc8a9f6ddb74999551f0de83e7aefe747efc99fcd2b9de7fd2894a3f6b7f3862a557c09da523362b27943a1a5aeaf7e61676855b4f0c8603135c984e5806c4f2529535937f2565b161fe450386ab9e1072c354769052ad4ae00ba6c78b7ba5d23dfa9d2dac0ce9f362e333cb1930676278700f5d681186e3db14313d09970453b6dbdf6518f3ead238d80fbe34b12be63f5e7d5cd434af3e553760052db2c8076605f796be9bb3c5c30fd4bbc347fc028b48985764d3e63f771b8c8d3c0027a1099141da0edf27b25b19aa818ce7914354dddba1005b823585fa862a19e3a7b2b406fa8dda517a63770ddee3e95c06f78b99c324a51b83c4daed8286643d43416ded89fe43de49a699d2684e8f9b358c80360e9d2085c8599236ea124cbed105da8045602a04865969cd31e69937c5c5310600c19e8e4257c9bbaef4a201e5d2d7c4eb51b206cfa2374e43dbb68761938960f1bf4c5b0881a84cce8b725d1f5a1f4dc2560962899154161986aaa8491ffff03753183de47db364275e6ac4d119c7d253bc5311f8768b3ccd585de58b4ca9997201b1a2d2963cbcf9b774a6952b08c2464794ebb2c2f54baeed4592e64a9f57a0dab2e26cd22f3f034c14356b8c58c7f5a0cac1f529856ad1574143491aa61ca2dbe5c4992a1e91e63eb2129e31c3190f3f8bba1f2d56252b5092f6087f8f1697f35638b8e2507cdfe8858028f1619efab886eac2d871a243fb5bec2d8ec1d3a7952286b6c8face81501112f2172d1fd6762eddfcfee298876ac14383f03e8d405ef487874c469776bc7f5dfebb769c652c1588d32f2bf760c94c0682bda31d2e1fea42340502db28abfc4ecf8c5e8a6ba39b75636ceb051a0fadeeb606cca4f86fc2c26843623c2fbe86d225921965e3d93bff29d0195be471ecc923a50d8e732782c745fa71830a099ee87c5e2c098cd1b09890a620fb5e6226ebd1e67830a128c41f4dd4261bc06acd2b0ffd53b1dc52d5268de1db774d737f311502ed472d81bd8d34d01acba4acb79bf423b4222f0b1f3f7631abdeb356d01d35b9fd2f5dd44d86978eae1f8968df75811b18fc9f613f8173271045eac8630ce69adb18b9df80afff85b0621de2837b6248fe0d91fbb00b377fbff3aeef922ded36c496706574389e83bc17d285df6a327b32b1d873909a9491b5cb4c0ad65b74915f06c9e8a79d9dcc7ffb6f04b95ca3272a26bd8298810cbeb23fac44ee6a9728e0c4e0c08033c9d92f70cfc9ba90c9bcc5869491a1bb2b5a7a901ebb18179b2d4ccb9c82f236cc035c8a1693d4318b5194baeea46640a77562f441aa327e9f045afce8a5840f84991def47e2e50f60d9e159a7c4ab39018712d0ef4228d1bf88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h96738e440ab9d0bbb1da442237af2b74adb65139ba622c338d9f08c0cc1499f84c9e78272b24482287c9a38e53fd9f216b6e116f2d84a56893dd0a886ccf99a4d58d2ca443205c8a67e688948dbb8b74b4aba0a6ea45a5c3f31bc24f2777299684b6bcd00b51c6dd812df250284c45bc52db9aa980b3ea7f6359fb7fc5446a2a8bb96cab051de1d3fd54958a4803dc36406f56b2e140e49f88080c8370f048ab827dc422fb261ff78861dd0865e6f412178c8900722cb6836eb851361b7678653904d59ee96f659cd798159e2aa9e92587c9cc7009d6176112018119e655157ce5f1526746b4e99bdb3c825ddadbad2a9f833102c96c3069a0850d1b129e18190f282659c57f91141b13e716b07f2d9dc222ac741c2290c476bea1d8717d98c4a19bebce7c446a6303524f30241225fa41eb039f9b3681cee0e55765594452ca67186c1323e4ccc79ae6dc8db007a963313ef8d60ee93146041fc99819f05125254d67a8da9b626251504cedd9ffeb49a7b7ddf686ed4013a771f54342c988d1af2f42f9e2d7469d9a4f46645a809d1a5363ad8d6eb71085a7f5c4f580918c0b9b1e62f656602a631fc757bff8b70b427e76b0932469d398621370f803a5b9fd196f429586f070802978ce07df24c15907cf8b23117ad1dd8c8406ae94ec27c1353b26c8050ac50c579dded14b7cb91353e9fd51f9ea71e8c3823c09385909673dbb2f82cd252ddbeb7be76088e47432843f2817d4b2fc9f9c5b48342a9b40b17181efddbbe441d7151871c976ef0dede94fc5e27a456e3df32780377bcf9f9bc4b36ea2de01d6960786f077a2af8d4268e0d288a8008083b9daf57b02b3e05aed1fbe0e7d0fa02c4e3938cb3062194c8c873c815e8d473963ae1931b359ac49687c50f5bccc68288fafdfd1e009c0388855ae8752d538da65b9240cf84be05fac60fccd2cf9b9856c305bc70b558a0e7fde961d20ddd11f8458ce8975d1ba2cd3400973a268810783ba089bad7ba736d70770109941ecfdb2dfc5fa18d5cf752980561d06c80ccb7b1813c222f1286c14518ed734092d9afe51f64ca33d6db526308bc83e35475b97643e9a127210f4f7f2c82ade79458c26d5651b02b47e3f849f85fc782117789d84eeb002ff7d33c5515827e2827f8c912671d8788f3a9392379848e21f60aa222f2a8b95f12ef9fd480f69def768c9819a24e58f92700f37b9428a83c7062cf4bff655c5243a74f3da3aab668db0bb6e6771c3f1f784d50df2d08440d175836adc86dba4941cdf12aac108a893fc81a6c8e040f2664bec04fe7695f3b6629cbb039589bc975382ce7a33547437ed7bf7f5567d9e55e710888adf97a08b2121e2e9adf9d068d0aa29d6a8f95d99e2cc68e0266c7eb38035a7f49111376a96a760c5c5c5d97e43eb01232e0fc806abe780ee97e2e17ae9cc8d0e6bd89f952a3ca841e8029134fbd2ae87cb2ccbf819511235ec3993c46dbc880be8a8c9156cb462b280d491c6a656e251ebf262b7cfebc1372eed43fab5193456b57c7f8beefd657834b8f713ecde06180cfd59295bbb5030c582651dd2ee39530ec0f76d4d953e2574dd75b6c42c0333afe85ae825d4969902d1ddabd7c17717c1ece05168a0c48a48211e6458e0987f173ab9abce0e8b9d7d9fb7576775f61aa375b75ca472345cd88a43779ab11b308b7d7ea1dd82ae7157b5f6d9940cdf38255b04a3a33e79ffb31865af537b7bb654690b9ad1187952ab6ab621dd61c7af7cdb80ace9557a4e841b3a70ef55f9ccb6add8cbc1b50ca359de1be26be5f21a900b1cdc469a1afc41844fab6e44fab61441ef2deb0a3101f9aea661248501d347b82309cc2941d38e58d3a2f6fd849bd6adc833f5af08839ac6a99e51fc5870b997eefcd1fcc8c3bd441a3c53f49f4ae24dde13a109763487e7d8dc71fb5dbf086bb2bf6ff8df5d7a121c578c6a94ef2f4dd5aabdf0f5846f0e6c2a251f9a8c13c6aadf628f7bf824d728a40d4f68bb758217c7acbcd49ca5868ca931eca3e84acf25a51934b11d5fd31474e16c1819b926d58375f8b3a0c5dc193dfe1655962dcf323af35eead96a1da24f07c9fb9e0b9d5e9c0bd0680100d832b3fb9aada52eb82df8caf7599d60e87e6cd2189a9759ee55e353516e9c8474a44d861f551aa2e22e6738b1ac5606d8f55f9cdc24fd65f2e9408c1ce4d0ea78c6ac1a2ebc5d8335187020c778fca425d7189ad1f9c882ed2d368f67d3da81ba26734ecd0b70522231bda92c7d34b8b02cff4e5224e775f133215608223243fcf69003febd277b73fd7b98baa27cc6d73fa5601ee2c8d6fb13a8a33b363328b7b82d22dfc38e1431b62528af52b51117c63aedf903c681ecdf5b661bcac0713fff0aa6290519db7acc08610ebdf0627e9c6cd4c5981eda55a2312140b30eecb0d3623ef115ad0d0d855b8666ea13c5f4e0cc4f7a230285d703bcd001571cf479b32b32631e932bef519c90048fb59c5478511b11ee1ec85787850486eb96a6327a00cf30788da5ffff478d5cd3b6728db3c0938621850cd4114342556d7af3fa467f46d1c8965a7660c39a11c4231e9484cb2fa0b7a5067dfdc0aba3f46214c99f72b9b2c051f01c470b4752c0e7a0831b14e3307e969195a4cdcd95d70b4cfd292a154c20fd80d30b43c3c3b7dcdff3561b200d477e560f4c9ebf6e69c8a082c11fab56bf05b2c199c29121632a1e91a489acb33cb3dd386a593ba9f816afb3fd3d69bbd637693e83eeb74737a61800acb7933f7f2ed2cf584ed696679f84a2883d623a4cf53d5afd099ce6c14ac4294e0de214f86bea61efb8c41d5f4dd02339927c014c3a8cfb687dca562791c626a53cc086f5471ff248e8c907fd40c96c3ea77624b1ceff919085cc17bef27745b9337d173cafc6d7e7595fddce552696ae949aa509a65774bc963a22e23b1572667e90b9f26667fa4d23e5d62408508901a280ab82bf0b8b87f87bb98c9e7b7a25df10781b93e7d19476035933acbc30603d448f9a8db0c1c105496deed48c6a58c19252a6e7576b174474bebb5e121387398c3b20a6c621d32b921aa260681d66f0e41f1a8cb6cf7e0b9ac864f50ea60092cab960916003f4f902c0edfd13eb72eb1a854a33ef4facd150ab7d7a1e84ed9f707fa3e291dc1b788bf2aaa510adabfce7a369eaea87027df9ec6595d23e91963e25c54fdcc8cdcd7f76651c121749f92540bade4c3516ad6c2f6c704115e0a5b239e5370e98f187bc2ae511214d99705d8e7899d094a43a260669d506f06b669e233730c28b7251b076b8ea79e23c97acb44325483894812043037bc5461dec998127882c6594cc6a2c81b62cd991b0ff073d79684d329e7c1d0dc0bdfb3c9e4de05cc6989a1427061482593398589706d0c72e300880771b5c5c48ba355070184a0a324c1bee712e5598e27d6a10d3179c785db0a1f57434314dd441dec21f419b5ea07e4903e84a520a74b9c6025408032d6cd4f1930e41fb650ce1a3bad243cb57f8f3b5644325ca75e3e3bfff8cc5a8c64b6aaa34def6964cb63170dfc3098aa2e8b5d6d5bc597c211850f90710efba3d84212be0b037f7bfb0e96814ea47c92e102f27c84c02b254c18c878b3fd6eb5db89120054e72a867c65a88f1ec55da6b9eff57c9f5d594e11149992fbe45d0608d248e2ec9de7bc4175ae5f4a1ffbf4f7b4be377376f246e98679976fc627ee7b4b52a4165f183d26a454870cbf83e07d24c78059af8ee97147b6b37d626d8cd90b7a8389f4008ba66211d02d76c1c3147112403d8e2d04f04c6f440ccf466a3c903f5e963b8de5e4a80ec24b0c4a1ec727401ee07446e0758e1340653650cad853e63506f3f19e3c28396d037e1c06612a26205e80b302e660e6bb2a65811fd11dd2d673c1b4f6d057150e92010e3b7502d6880598aaa9a4d973cf723d962ade7e166c4f59a8f67e6033352a02b22123110cab53476dfc49538ae88232bda30427b8b89c3c1b19bbee554955a0b38dfaf1fc5b020bb4b9878699bace3512324b5c250a60c12d1441e468c4d852a4a72023d17d3eaac86133459582677502ea615a96461205ab8438274eeb01d004c43a7092cc27c867f91a73776865e98be2e33e18364b26558ee9c46574a0ac1e27fa7a79f2619743cbc8046cd8910d95fb170c8688c8f4fbcfb0590a2a106e89cdaaf9ac0a68d86ff5c1b0c5ce26dafe5da683370c647190465334acb138d3ad6e864d94f72930d591f536a912eedec123b3bd9cb13ef3b2d34c6be35f05be2a2f3fb9cfc9a79debc39b55caba641c656279b20ceed2d2c3157e8f673d0738daf446be0f2b9ab6496aa386cf3206c3f0d2c383c81e2bd748dee766f62316f9dd66525083010d8f6eacc3026004571d8083133c31b0a49ae517e6c2406696de488aae76d15ffcee23067d7f70f0f89acfbbf576f54e1373f28f713545a617fe9df8d49d70877af3c3abbd945d84ffd36811f9acc5b240c4ca8ca1c2ae76af1a32ccc67309100e92c70579d0bc9b9d4284da10fc563ede1ce207e2368ade6fda799fa5f31d88ca1ee987651076b89c74572e47880acda0b9f6f06d2482d9b70e2a76d2f48c0e7b7a4f332834b76bed0c7dbecdc3259d055a954330073f3ed97e452a45eeb460164986ac07242d9591831d382644f218d19a60812b73b30bd49817a21232b0226c3446e54c94873730011e394d00a7416efa471653d28c8a28b2d570cb2e92e7403e804f4b40bccf512328ef0f2a09041b500fa883e66af6699b19656e957b27b60b334f1e8a7e0a27d147994dd11f7cca145bd1d61d698af0de9a200b772c16d772d511a82d45034ba187273e7cc1c5bb9fcc3514bc433fe037e3bb0555271339d3e16aa0d1991de013db5bec61530474d6b57106b3e019e876c558df44b0f3a6ea4d1de11583f70451f93f5d0ed97579a54eff16453d4bd73046be9f374ca4452775aa76d9d8ec26e55523592f343b6be9bb8fc6d2e4fe2d7add1e3df6f14556aad92e7ea9607d9d1c8c4cce9e96e0b3370d9d5d8ff793163569b5ce3b5ee35b80060b71828135c6380105515886b955966db9e4afe6a9fee546dd3f67926368f544537b91a203e8f0af099bd56577d35c9de11c5ddfac56e9fbbc6c57a1a7b9e19c304705cd49af50ee3da7124673c065adf4ea4bc3086322f195bf3737b288db508ca5835589d0705bac4035a2b4b040728402a53c75e0f58bcf137232be70b7eb565ba95cff2565099fca2640a47dba0f036b002fff2dafe1bdc36b05340cf9ede4e2798bedccfdd797e6495beea7c6ac879c1dd4176c7e6db12569e3469b01fb134ae906bec220bed77e09d091b8373f56a8da88382a8e27d77188f826fddd9bdac70ec981d8b6653c72d8cc535736ec639fc9d55e4a59dbaafb817a5e47e151d260c64fc4d4e0dc2edff554277d599291930f64b5bde8fb31a4e9d22ead44b1638619cffb78774069437db81f717c0af860f848eaf5c86bb204d4d0f80911b55e93e54acf8bc78899c9c120369d522ff08be6935da5855d83499854565910483b7893703be50051b2e1a91a3d3cf21906cc563cc0c8ac4adbe48d608bfc5f7c49ea1a53b7ddab12f134dc2403c80b4bc58bcee45a73752b14e9fea02321e1701f0ea1d75d3b43be2f7401cb46bdd16c73652b538a1a1d94511b6ef402bd6da928b46d5a7c2015b27735d7abea0af8ad1cd0af3d4888ce26f46581370b089ba728e80b45c209603f7ed8a268e77f01eda5594477f0519242;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9e9609c478a0ddd207823f989d3e9cfa65ef2acf7006a68062eaffad927f7937b7a552ba5db3a6670ae468722581f5c36b0216d52fe1fb2a88e6c43d06cd3dd63df2d5ea15be715b877d2a2f96ffa718ae1b37b2e0d35d25a3d4982812bc32e3045ac52245183612dbb14e2aa531244d8ba6d39d4233108fd0e1fce55092c31c402c0a5a23190196d015690fafcf1a21eae0380d0c54c46c3e25cbdc0e72b55374fd590919fc7c92048d839cab52a8d1dcb197db3c164547fb646fcf0b368c04e9ee449dc8120d618550d4e16572cd6d49252f75909933c073a5e49f05669a0f4fc56d4df401132028d437f04a55efed0e8ae9dc47894bf8ba74ed31e7a241488e7619d2eb059e6d9a24efb3a2136035da3439d20933e1cf842c32c500032e2123ecb61a0597e4c131620ccb55f06e6b08cf71f9e0320d901a9b9dca93df9c5e61c2a5cc5ceb41300b63260f3543ccd081a440ee5b1dbf2e9ded1e4f3d2c0f33b738dd71756ae815ebf671762ed7b2507d9335875f675f172f9973adeb5c492386e8f2bdf368150ab2faca9119c32ce950f8b4fe822bb4ad176b34f0e147785a92418704269f3ce3ad38d04eccecd8e1ab5d9f10d1163258b9da4a67fa524f95c07df9eb97cf26b13b9442d993e876947f94dd4206abc91f7e77088a1c48c3a0d693f32283a66a864b45d55f67177f2b835cdc93b5c18954cd3705968bef65e46b024aeafde53592c11973c2d03b61a959019b58bb01b824bb9a79cd82cfd7b4c1881f777f3ff1770c1155541d2d53a02bf25e055ab97635ae9c6e4b58671afb9c3cb69258eb3b333716bc7977e47d191ad7092cee131ba6bdfbfaaa8e6901408365a3d5f5fa8a6c76c03895b1c0c295995d3b4406df11e2b9a67ff69109cc72e90e23f0c148ced348980b59aa613229b6c5f3458c982c842d69ff59fd7cef9de1d14ce32ec086faa078fd675a558fc3b30f3736d06fd1235d0e2d46424ee50fc21c5070841764c06063c3b52c0176da18a19736822685a4c0ae99abe6608db047ded95c506d83d3a22d392bc3adfbb00fa24d510bd993688b4e22149d80482f9479fd2fa89525e897173ae11213adeeadad3339c5ac5d2cf9c567ca57193f72f5681e0cdcaa5c2ed00be007d65f62e8cc7df803ea85f260d19689162a7e5fd096ba0f84b43a8496f8998e41087dcddbe8a552eb684a9c03dec066887940ba79d44ecc78c3b03e3b215af192a98d10636cba7772c732b9b3517aee2c97509cecef2ef0b03ba7ea93ca1956a2ff2caa8dc4ffea8a5c02d54228f76e94662d3e47d89c472a4d8c00c5a2326df31b1efdd5cd49f2cea58e99222c1fde45036cefd8f88921c1ee0772bed07b9fa0948af1dfeb3afd3dbb5200cabc5e0ffc9321915d80bf563fccb9319e86c0bb49a17ffb81800e287e018aeca52a562a68a3ff25170343e39de5db08632442947606f5c4fffdd837977872e704a728e7d66d4da8ca206debacaa3aaae62f2a66d58c608d9ffd6706c5c209a34626d9c953fa49c983136beb0788b60d65e7951695aeb1c2c03b544930af0d8678208b10bce46940b69bc36e411bbbea08055f9412e7c5897d0c9efad47ce55c6e5c05733dd9208cf6bc12b232c17dcee8beaf54a54f45d7a74f35c85d46851776e5e3a54aa260e3fed7aec83626b8e9f04aa3c43315eef746b8cab5ea78cfc4b3f0a4f4baeeca6dfdb6f90f53d98ad425571c55cbd6b14fbcd5d7872294a8276e955ce86407f01563cb88b5de0f28b255b6054ece125d406aced3650ac09eddb7a4f00fb378a475a1e7e8f8d32ddc908467289c05a5580932f62b015323c8c8daaad5914b78eb525ecf4aee0aa31ad03e56cb785ff2bff748a6b02b6d4ce1080448203bb185cc70632f7ec245f8578987a8eb960c3ea1b9cbd385c2bac962a6cdbadb68652f97be5b122b8e1f8e6c5c5ff82e790412cae17eb7e34b63be716391090208b0d6847d661b53a86d169968d207b617bdbcb959de50603f6e07be653438caac21ae0c764614269d9256b6e92c6fa76f6cd66dea011737706d9a17e0effaa0c54a5fa955c7e035ca22b0f2176978f4d5f6fc40f99efc765a5cedbce848183706324efe93c7cc5d591eb999af3f033ea2aab674573ce20944aa17de4cc70568ab478ed728ec6de7311353dd21b38927e564832604945a8e7458768672ef2ad571c211c94ecf542cc74d6b39fb7edf8088ec8f2d70fda490b0ac1c465f19bc3c4d03624f4a51f1b4ee699c84c7712f7d4322d3b7f893490ea91877291cca409008eb16c73de68db592c678c1bed67151367a2f55ec2f7e92eab25c4ead90b55c91059fc44b0a7f428da0e0646d15968ead36a86aac5b3a2d7b1d2b6b28097ae0610d0726bc98f38c29663a8047aced5638a35669904fcad603c28b9b9b305055245b80cc4575eb09ad07121df600e268ee9261f9a69a0968faf5e4d65c66c15f314eaf458badf2e41601a6abeee22ebab13fd8433eb8f942c67d7344c9602101e3bb8785bdfc492bc7ff40944f7619af688f9e28b3d34a804603994085eae7fbf2ffdf9337de737d24a183640ce7f0a497cf201699110ece73fe1bf8fc407464bef41061815d19e6edabc321351862dc08fb08efa74d2e83f8561bcfc4dccb5bfc0c42e7b68e373f8874688c6ab669862f71f90d71aa8ec2ad9608b825e81ea8ee48a61ad74a1100689160dbd93076dd50c7624fcbc7af35134b128bd423ed85b8fa3d56a21e99b80be6c4107b79201bda092af6c6ec2bbc1ce4c337952d535db0e20e3ea14d72e00b8f6f736eba0bdbeb131460dbff2ec5de4b1f68df172bf1be0ed9cadf6d7883c0afca8e7ade7c8c0c56d6b14cfd540ce7bcc80f0540753608e6521524aacc60adbada8b5db1fc09af1077aacfd903c398941cdfff2b9a39360ca03f6e1e490fe1b21433892962401000b588704c9e1129ba77228d2db197624c1b9415b1927d388b42f4c5f192d66cf47bff8c5cbc4d3ab273352bdf32e4ee4409759c0af399edfe78fa32d421fead5092b4b05cf15bffc76a30c9de60d649e5ed171bb75862cbb4e1e97026101081abd63a432aac48cd974d11d91ea5c0014d389521134eb47fbb4c2ac268f129e58c91b69c3f6b39145b716c4e56d1c835ec87294f1072f66fa92595bce9e2632ce14e0052e5a6441be101cc50aca356badb66f7407821d0372ba1e822e37a847de6e936a801a46746d69ec58098f3f26d693786c603902fcc7e0646ddae1cb5cf4495453f422f44ecaa6f3aff91941d0666e5b2782a6cd0be68c04c97cc70eba58fc224dccc294b47c9080a81f2d01450fcbe786b2d341eed55dc0914a52caa9e56548c08fbf47efd0bb11a08587296c8b73099724f421f9557b9c3cb961517b84a20dbd8b268b9a92e7f2a54015d3966bebcaf5d72c34590081b86fa9eec931b78acd4925ed862455565416930ba1ab42d0fbd9878eef3c89b83c651338d8cf412014d000feb8f2e2f595ebe26f6811ca73e87daef2820f196a09c89c1562cd02135dc5d879d6938c36069c0f9d2585638b81484159aa1b795a1db176299dc14b5f7088afde8d23645a139cd3838401934bdddbbb2604c5f8e36d3cf7bf48852a9fc854de29ebfe3be01278d12aa5d42fd3650c840c084c7f2e544f3c15d41d7bba79b48de0328efc414193e9666aed71759753bfa3c023d62d45e0c2061f52d6018774c459248a70e65a6281336f16a1c7a2c997b2af67d5f5a31ac69fae1386b1eb64a61d2b607015adeb08ad05c2d7678a5bbbc961b3795eef481a1879ef0aa16dc1c16eb2257e7accff100c4e4be9ef445917167b9e5487c4470351046158af7f33fee5e3fb156a2b8c9195444b84ddf28112a7cbfba449edbd16c94c0eca4bc311e7e8f70456039197966c07f7b6b004c41abcb65d5b3e13e7cfb1489e2abe15911ce7ca5a3d8f87b04da9437f5c607af2632f6664fb197d71841c05f79e39a27b52baa8e26882d453186de07217d7c1a56915ec321d33f3bd8f8864575c4ce173940d9dd46b9e9f7458c450346b736c308f7fbb9fe6ec9759ec13bffcfb0bfe43523beaba4c6a4e1681d0e89d97d28e94a4e974d28ca48cfea4b645b7ed0f785a74f79f0e1e03d3ec8dbcbe51b97e4e9b607708a0c037761850b6bae0a10591902678bb7e53fcc73d228ec41056a0a3b6d888bae8b03c11c47d35e10d53918e00facd1e838c1a475d6d1e88b302e67fbed59fcf66586c343c67d02d75fddf187c4db36d4ea4bb1d0b2b29124c25e9bd2af784eea5e18bb53342106a3d63b39b2f3c401aef6918e24e7fb00184447b7d973c34026c8991c5dbab37708877ca59757a707423e07181ca61d14d65cd97778a49721f9a48b206f22a3a3ef3a9916f90039ab79863254ebe49fda1392ad01ddf2b80670207b8ac87f51ecfd5d2192d1c5a76b3d41079d763fbaaec23eaddbeb3bab471199531ab9edcd520adba46fb5599078392b65f5723be58734d99da6181a06e6ae3d849249b8c8b2c6771a5496ed256760b2d4f0cc4c7e1ad25bab3405e1b0398011dc1a35f3cb340a6a91054964442138e59265cef9e553c062576585b692d88e1995c31e3829697dece11556af401162355d10181668f45b4e81eef5753a77dd39839821cdbde44725e135490b67bbfbf3e5621277edddfff270346a8d14a32639a7877cd8a4bc6a88b360df334b3fb57f3ee93405be731bfaa5265eca838ecf34c6cc889ac886209a6d29df2b74e8684b8ecd79d89dca5026bedbfdc9a8df146c646cb90e12c1384f41a7e0f674ed6494b3f903dffc21193a1293e97d49279dc6226521274b698db30f92d8f4046d12bf622b985a503e6c5997f83d5aa411b5387e3798cfc4492085879cca24ba133b7205ba1d9768d89f36ac45981b94ca56da2b6b0bdbbc4ed25f4d526aabeba8173829bb02f525c2ef4a9814539f3534a96e9ee314c00bfccf88924e37f25893767e6f2c12815475292f75f91083885c9bd8e0d002bded7e38b8ea5a0a19ac611562a308f36a3a3d87a19ab6df16519a9561404603c7fa5f2d55e4a4f0ed5ab19b999cc0c8f275ba81c180c0d4b3f564f6fc8f31934a68cd41da9fd2bc1c857828b7f3e4968cfa2d6ef68279e40173802ddd3feda32fcdf61a077dc276690d0cd4a86a9285f41d49f4040361484926f680e2f27948e82f55601e6326f190a4b5713074db7a566063322ed007232bd5151e6b19789f89087190272cb77075dcfd2fc1725f16eee5909a94d4ae13260d466f9c15c570abf49639c546f357fbdfafd4738da433c4b99acf59fddb0d50d93aa9e5555141f9e8cdbcfadd00a24cf65993749906752fb6ea74d0caf8927fb1e3485e9a1c2a984b85234cba27884ad47f52e7848a58c86e8a6122d8c9843b8c7e31f648d9e786abfcf1fdf58528876594acdb2d9adb9731b1eff808cd013860aed880a0e712b89b9ac997004163b3aad87265ff83e4a5f5d4dafdf8c317f3109175bb43aef744224ddca9d4e594dd84d9a8d577b7e38df2301cd775f7d96d596bd562c1b0bf33c5504181d6043cf0a8ff9d288412d375bf95835a43ef95978adb4e6242118ee95be1f0854422c216e06f90c58bc751a3666383f29ce1e144e3f81be02619f01cb2974ae2f15798f8858c2cfaca8a9aece38e38f4055310d0d57a0178000c75a4872bb8e690b71bb79fc973e38ed7a61183e974aa57b07af1b81fe2f613d964e122a7a87c09dc386c03870897fdf2a8326d7178391ce066aee2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hd1d096a1a17f37414fe3ad95c97188487fd180dbd5c4f0e82421d2e680075092c22a03e4262c6098f9b285827539d4b628757d4a90417fb3dcd66316ff4ead430fe56de294a3bf962b85f9d1e63bafb60b601940fd286772e2a654249847404df506a50f6726cb599247674de75c62f060b330dc8fea7a432dc913799fcf7772643cb84d8224fccbeb744f8a220bbd0ae97513cd44ede28a8a6063e7adf3fa14958a4bdb0c215199095bdba6936980d85f5d7e8ed00f6717adc249e3e562bfccb45795e7e9dc492c5f5d23e36d912f4ed296105a6b2ec82de17746825205f22955614226d9889c76d2db3cde637a2625aefef773d5496a1b38cc63d77e365a1f8c68810ccc53f8f833b98738ee3b36a805f85eb809db0c80639f6c7bd26b5503a53210e5ad69d3b97ecf0eab2e5f312df9739af680802c199d0262dea579826e2e139efadcb7da560640c703dc4a7719390b64885a7b49e212486fdd2bffb2931954a3e2fb34740ed132c8a6ed0c6ed33f6ec01069e23d40285d9fdc3e216a737633ec25c475b2a2974033d758f1e33d06657105c009eead1f633fc8881c7a2ed6048495458c03b2e3b5e99da749db696471aa4d7b39e42356fe16d583bae0038fdc71d685f989300ea4b90d54fa21902480bd7a56d72c38fcf5a42a8267139e88edf87d90a0c8721af950de97084b0d52239a316eb0e17e948e884dff4d82b0b39ffc67912343225999a63b15318545741ec1336cc582dc7a1987f2a4eba49aaba3e6b1b04cf7bd103683c5bfada7b94d36b3dd7c9bcffe4ea9d9c736f819127471c78fabda3c52821aee5150037fb33fac9d438bd95a8c226ad3406ce5809b9d822e5bfe7eca63c130c17ccf8f46933c976ed65fb7a4dd237d5e69534220afb67b76085117d9e51513832c37b8f43e373e3c92bae928e7b9b03fe958a3d977c33c79e0025aa5d61458f9af4f1ec1cef902228f8133a6fbfe65413b19e2823ca7f4bac9fd40bcb3b3cd969b75ee718a24641fe13004ce64e4c838c5bc52ef2eb2e2c72c7c6324b9fa88d270c1f895d4146a0e41bc81c22786338e5e9dce293fd1736029b4a8ef66b7eb35c76ba7e9b618b5b09fb6e45c66af697a76d93b87062312ae2c96c79d703cafa78be441c12948156796845b4614625a2b5b5ce525e3d1284ec6be7c898a51ecb0396447d1c02517684314b69ef4cf4243ab87074475f6c4c13a2954b74a09e5bda466481cc11665215d9fa223c52f6a0487d8c063b012712913fd385d292d6d19d0a7510eed6b575ed0f060153900753a4722aceaccad5456728f917afd1aadb60ebd72dc4b03864a9e3266474fb140d03ae7c6f43665d356519cfe0e1e8bbfdf38a910b7bd6301caf661fbf8931e3bd72adb574a42085b435c1089306be944497e42cdab5105de61d2a338dfa56fd7563546186420c9d8b6c1becefd9c037daf126cbbe9eaef0dc5225a626ede8ebc1fd912ef0db97250771b08563b5409bbb173bf14aea0efcd9210eaba35debf5f84d6c31dfbc849910a6385a819826ea03cae72de3ddd7abff62e085be38a2dff70deaea79dd4eb7c92f9250dd1d6124a0be98bdc352ea127f00b2faed9140b683dd0ca55265c53027d84f43c87d528349b161ef537c8730be996e67842e1c2d8e0a8fb12ad1caf0d14ab70751dfbd55be39cc9faccf52e94ee71342fbba76abc4c46ec5bcb1c950eb319c9d01a2daaae4e068a7749672242d3cef463a4b9b70e9a98c326807908328da243b96392e9972158f38f8df6b98a6b7ab1d86aab59eead806932ca2760912952748723bb7db5a1d884ed46f5222290d6d5c9d27f6195feaecf84510b4abd4d6173218b752462ef9116f863a55694795d370cc19dc5f523bcc35e25c083372ad8c8376b422a64124a3cae1bd7f4528a6fc8b718d61cc30a604abbb7aa2a8145f638338bdcc2b4fdcba915cb4b097fcd26165ad92a3c3aa1fdc54918df957d8ec29e049aabfbca6e2f6b1f77b24c6861d1b45f470c990917d8ddc82bdd33e409b79f2649292e6acfdbf7c43011bf1156fbc142c7c3424bcf3d27bd9c8578b07d4befdd8314ca00647d66c651055686b2d76b7acc4dc9bf57f6b051846767c8f9967075de6b74f8d729ac5dd53ffd039e2e955be186fab6709411b178117250b14aa5ecd1675500a3282c58b5dfb50d1d9e42eb3702195a6e9f558dff448d73ce10898e93b96cdf399edcaca1f4eda23dbea1ac5cb56915a0fb82f15b5146047f74adfa2a869d327e5399333f07af52e7c1e7afd2e05087388be0c249dc3b289eb296609d091af235507e050c10237e4b2ce6fa6065b08912c1f70387029d6ea69c5f0e259d00efecb0217d85b0f1edff920b30ca7c1e5c0baab9d2d5e010cf176a90689e20b10822d82bd4fac7e7b791022f85e8f53821c3836277846840ce51ab8c800ec011ed94fd8eca70aa3a3d5168ec4f308db915da1635ec8f004fec64670ec19978c8ae070f85c5b7f1ec5c5cb81f26e9ad0e08cd69b740592e82513fd2feedeb4579eba8c6efe7dd2cff251c471d79f7aa539cd70db4f11bf7bb0268aaedcda5d04a4ea2eb5fb79e34851fcab1222b0cd49ff5314a819aded21903efb9a016a67a56897cf80e839098fc930d27b754d96b7db092ea4779ab795c03d07db1eb277e9bfef941af4580e2b080e3fb376e4d12cecf7633919630425bdbfa6f541bd1a5d7d95007515bfd38d8948c9024d7cdc2b333b932aacb270b60ba35e750c90d008194d2d981d4b49d703ab6c50096d355807ef3e08f518e6fcce18aa3bfc5ebda59870b6b4e6318ebe010245f94d7e16bb7fb3e503d6c83b46ccb10e2d642ac24cd2792c9502555d799f2791c55da2daa12d1a160d2854edbdef63a5a94ffcbc858b42491de1c4dbf01c6c0b6438173ca0480a48a60249ca362b8eb9e5d6c309df84b4910f98a20fab65ea5bb6ab74fd0cde5c9457d7202b304ab77a267e7c5f0371a527b254a66a40f61aca0ff50ebf6ab2f46b876fd8f6dbfee2892fc7ff922941d38d149719c232fb1338a4f3d105ff6a5cdc670adfd60e2fc98b6d09c1631ebcecf36ebda8b908ed8be861e2634dd5d6f5f9684e865aba5d96493a73b38ec40b2d125553e2bb35d9c7d8a5d8919b92d09c4f1d90c538981a0e201ea1f33e713650ab6f08609decf360dd3ee956e91b12ebba5f13dd2e2831c16c323a3c28d8356ee2295c631f10c01fa0296c8b2e7ae4e0c3436183de50b64e03271c95d957eb74148df6e9247c085e53cfc3e5747e997376bc0ad42b40b1d2f26fe8ac26c571eca4afa6060e1abe236d49305f4f5f59b6b29173034c638be111bb8084cfba9bc7a529f48ea0b7f497bbd8c827000a013420d33dcb1e29e6b774bbb04223d5d5213ed79c3c09193389afe9703f25bf1661b6f20aab15442360d0e8940032f7a0a53aa0899034b4cf91b00501431dd6272060ff6f31616e21070b7eab89dad68603cf0635b21cda38a3cfda94aebdaffd2f6ec264beacbe1de15414e5f750fb7a004e6a3d29a642ce8a35554e3635736b0dcd3948a3f426b2834120bc5da81f8d4c79062b09e9f92628f943566f5dc05b37ff1b37e4a8983ff5afc82973d0c30bf7a04ee331d0074e45d5cb54e5c5ab2379678a6fac6e63f11daaef64967fca3370591fbb7b5d3193fb6538f0f970a2d5dbdcfcd0c164fd80733d58a4fcaa2b921c735b6a19d1ed7753fa13fe5a61788d774cc1ff26357dc5cd0e036d720b59beabb7d314479eef0ae390d0f1a4c305e00a536785fb527da3eb8a9f0153f558b06b6d72021af0cdc63618b21686d5c2a7d8ab8390fcf1e6d6cadf7e29efd9a78530fe52e307914d799b36e081cf568142ac68af35e9883203faeedb0d88777ce9fb1d77238fda19a65bcb63cfe9fcb5f87aac6fa60f1cf5d7c9eb0fff5c014ef30306a58f37c6ffa788aca8c02bb8ebc90ca8c904a3a090a4ecf587a409275e2ad860b46a2bcce5676052af730beaac461a6ba2557e1028ef6678a3e90abd98cd87772d64bc9c1005b0518d755b2f61e80982f303bc3c0f77e6b1d97caaef58796ccf00b6737a7fb4ebe027e9a0aef287eb4cdf4847bad529841f49d9f54a9c0178a70e2293606262110f9ea122fce62e392c44ccba49bbc75c3e55ca9ec94c60cb8fece9f2808c75687e2381a700954a46b79778c2373ffbbb93a7c1bd23f5e79af672c56166e8104495e2d546bdd63921a8b27b50386a1422293487887008324337d76d4e49002d51af3174b7afa10d2f6773753b72731bc3b5edf160c734df3a695af7cbaaa90f978409dc6486db9607b7bf1adbb258fdb92d3c6772287908571e7a70407774cca5a9c57d5edbe07aa9301955958f1f2fc079bf3a2b7a9bd29f34a01a1d2672173bc93cbbea629efb0cf50dced2604167a65776d66ebea05fed9dff98e9105033224fd2d93905b093848b143255fa83c83da0c8adcb26a4203917c5dc0fbb5045d93931554a160fecc3d16b511c2bac3853e9ff1f11e288a0c79352d78d5f76a6344b158c4656f34d45b0bc02f41800e58a1b340aa902b15989966d5d82c572a0d70106123ab503a46eb0cb35305610fbd42b6c86b9a0075818125486fc9c58683053e183143200cb6cd1beed64c0159fe1c234214376c4341aa26d1f784b1cfb7874b293c9f94929a5b8cd103947bd4e134dc366f8a23676581ce480b2df8f0b646358702a434ee120a25085b3e92d4b6535e164a9fe0966a6978d4f3ccda4d28ce1d1b3af11a637be6277833d2b80b118b05a787169ecd2da9ed48955eaafbd948f2fbd90e852afd569295fd360282144dc9645068f1227b635f9b7467583075e3c2d60c40a94d90204d00292130f8882ae7961aded5da9eedd8ec00fb2213d4db540906761268fff5ec8c910e5736960b926d769e91a594d4b25b411e4607d4c411bcfcbd6b7140ef7f9459c436a17d00f962cd9755b48dbac5b716f066cc9df0ab19296fd1fad973ca3cbf1260af70e55aff11750d8f7d7ff8e56069e8d4ea50ff8e1ed7526df136f79ff471944061096df393a2d5dfddf16c2fdca9aae71da55fb22c1a33ff6f0a323138442cfe9c225e36712240ef50b5dd6fde0494d41ef0a52004b1e86626a4e22c87364b35ef0352082c34fb226178a752200d74461fca19c9e6665b4ed90002c27e83fe68bea029d81b02e9064f586f7c63546ec5bef2b55de7e2381ad209481af55d64ce50ff44b4f42430c238369ccad54abe44e4873b0667e246821118482be13b49ffe9d0ddfb7f4596a10ad037dca9ac0d429a6e1d0e395954ea92dbf895873541bad1c3e06a0403d17cf2c23a52f885b286baff6d1142e19131cf283437939e1246a8d8987f52fe639acfdd629a3206e82c79c7e2e3a34d38b72a633a39fff8b8c5014d70ad93b03898b4511a5adc779a83cc628c1ee25bc19b68823c0ecc661f9da56fded39d50132d2faf98c4b5d519eb9a95c93c74a2a761d49ea5f145c24053b077821d0867e9461949e23c7d3ca495de50834203d8283018cbd0c88a374c37a420f08dad9913b470b142b5256fb1dabca7f268b13201f4220734a89bcd5a7b212fd0a5cc7bc92256746e17c1b1a442355e88826170c0347d9e0a09e27ef37cbca5a31819d60dae79832304a5429b74ee1f0f6e9a87ab8ec6901b5bc21f044cbeb2f97e39886fb59c54c0766ed875ef0cefd5a0cf7d26dbf687700f97784bd00a5d1a668b7ee0f72ac1c5b539ed50540f2dc0f164c50678c7bb653b295781;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6da64e84e1d1ba854964610d55856b624d8a70ab8b6b84045da01e64b22bb2252eb8f1295be5767bf9d491d2c8e1ddb77f280221b29862a0eccf4ee35846e8cae3bc871e44ef11089cf6afc74b8d4413746cb38c2ad799614808005b6e12ed004c229c0439cd12945643285362d048b3ae3cae2aaf5c71d53b4457f90619f245113c22ea211873682dc6664ca62253aca31565d6da18b1e78993560634588b6e959fecdebb01ac4658e9fe311aa2cd53d1acc353acd18db67dab96fa57c075ecd019adf79ce6ec85a9b465f181845a54792436451510206409f56bb42fe408047ea2491e793399d1aae609105781dcac65cfcf7241d751e3854fd30adc74351a79b5f0c48412ee6f9d581d7f36476214f5f9285eab5df74df79f3cf9b7e091ac1b347dc0d44b7662df9f378d5e5dd23aa01f55589ee89df4cd727496d4fc7f8e20d2ceebee8f61d1ad05810e4e70fba5e2558501cd7ec04f02a62e3f4caa0ca0acd5aabb989045cdc1c3e429e04f0388b13cfbeef91a417a24b4bc7c78680afc891a4b006874fba6b8d318e17ce7a8afa740c0660945e756df8d22e7f9b50f95909d7825878233c7d57c7cc0a050949632d9d9422d4b92ccc7fe63ac12e1d26fd4b01f82f37c1eae4de3e6fb6f1de7f32ee4e87cc5f9a3f44c3a78715f7d2b9ee8f9bd083c50608755e8c7c69abc795418b9229bdb7ae33fac5dab3690a5f47965839d904e5a1bf72bfcdf2ced428adf9558de2ad8bd3d6e08e8bb3d9b6daf79650ac5fde996a756470720348d9cf5fe72877c41ddcc02d68a6855d997465c5365fbc86a73d607443ed87757ab384ef81e8e26d7a809c901dfcabcea8bb90a3d8237001f526c85c917c522cec3018225cf23fb13577ed15e91d0ea81b3c7e29bee91e06c02a52b758e9e151516bb99e6a013c6529618b0b6ec85c274ffc98d0d04a7ce39daa0a979f233b1d219182b1d694df8446ee77254ef1d7bbb5a78610ec48e96a54a3a648892f5ea1334476f43e29aecfc159d67e80cc59c5bd84accd548c93b1a7873a66ed0747bda76674c5c57691309634fe9905384c37b1f11be521b1f992384dcb260dd4e4543b6e62b467716f01e959ad3530fd62ca64627cedc4948adfd19ab125b79d20e313594897e1c9c3069334ff90fb623babe571227cccb6f656b94086968e6e42d77d27877252604b43874c3b4b465c58bd3b0bfaf91d54ed8342e0e5d7a7864dc1d908dc896138db52648b3f0e845db56e2a08a86560bcb2fca58fd293637cdfd6bbc5f685ba8c3015741e3b24cc1782b7288e433dc34a7daa68b32834de9ed203e0b97e712172745f89224d37b53865651f1d48dc71753ac731950a063ae13e317908ef953e4a09d45bf9788b2056418af20de21b58d260db2e4efba35c055ba01370f33fe7b2a113440fa0cf56bdeff9f295cf160e42baa21c60dbf176ef4f59b35d3b02cc916d600bfb58082d4fc1dd643c69472a219d96cf78355b9d21a4c4dc6c354c2c0dd2bd1062894af72d553c3231affc13372f0d7ce5d476284a70caad18e06a2dd965a60c0539d8c032a37db47eefa389c4f3e29bbc3a5d41537a49bc6a9eb836449cfb1f6d114be6dff9dd63ce12150d44be9a30d41f21c20d9d2683967da9bdcac12993016809342da55e62472b295d3ccfac50ac3596466a406c16abcd369dbe2d873435a65bdf408db0fff99bcc2e05e840c96235968278884dd589696a00528f6d20eabd1920e06f5aecf6be72eae83fe4953b206f15e3a1e87911c227ae0228130cc968ab7bce36f456f863ba29e97a7247cc14b9405c848144cac3a68f3b1cff84ff32166509c7e008f88deaa25ab922f6dbf245adc59430c972b2b02aaab51cf6683eb75d8847710b9dd0131d05bdb4c7b5a663f75808cbe1554c3b85c9645f2413db374f54088b80f1c2c45ff88e9d896d98b58076c2f06a4202f62eabc284a5b459e29ab543d54a0a840780af2d56df053536f446e82fcddc38949df99cb79b604e357d8e9bdc1316f7fc0d98224b400227a3c8d7d885929cc755fb7998c67b46b00e375699c41ad59417f9ad0640a699a4ef9bd1d4a874ed5cf71af40701be7f77c12bdc8f1abc8ff5b5599f34b08203bfb64ffdc4e6d1abe2ced64386124a0f5ad96c759fbbb9b2c6d478efe0df361f0eec2a6451c7a78feda6423a0214912fea2612316225b92dd1d258ecea48df5ae30cf2e82512f3ad92d4f219801be6c0983e876eac2b9d4703c14382918516327c6e1d70c9f28d7a71cb31cc77aeec90efb3c3c7c1d2a76eb6c12e1b54ebb0f233210f131b834142512c3423993e85c679d597c5da7a7e0292285c8edcc52c9228e5ed77682f739dbe41be54d5fa92e4c102f75e888fc754d0a4ad72edbb3cbe519df20d3f4b1c68ef368a79db3f3ea0a1ddc271a771accdcdc22342114b7c868a9c4d4d4b6e374331b91bd1b11a81f4c598d87a3d4b4567d16c60220851bafa3919565f5ece2a69f67826fa33839ab4a59e9882790b7d0650149483e5d4250b010528ae3bb536b4cdbfb74a15d451ed56ecea1b57206924e3c7121f5bb00c3c5c4b1cffe87223ff3e30dcbf5311f46d29e3a91f39b3e9054490190d2a9cea2a157e321df95b326d03ef212249af553b82ec34166f0f02aa8e1ca2fad2509fd11a0b998df982ccc55d2390819aee5bd2bfa0a8997dbdf3b0369a303af202d417fdea721c98e48ade4ec909a09cbb66a00fee7642f0cf903c0e703194cf9aa16e70674a42351b0868c995847f756838cded57a6b088d6a70991c10ca84cda3b4ce7d0bd6a2034dbcd17cb58f7c059b1c280d4e0c39c1c7bc97d49d7bb3a293bf1006991a49f4ed50476db920d9a708bed94caf85b099f4d0112d51e50feeb1d7151680b012d4e4194e1ddf21e626129b2a9d707bc9c7c480f174dc8891c6fbd7459ae1136a7c4ce31258dc51d74e1fca2ab18ba63080d3aad70426d1d69c4480fd71ac30c7245ed94938aea34144d1db57c8bc0e18e65fd42aeeabf7842501fefa31118e400dd6bf4a84c9360c200f930ddbd7eb03884fd55922ad132c31131666c9a0c61139faa4f513ee4cb012fc73e59a5937586ce33166d575b1b93565fd12d3c65d0ea71ab8b8bc4000fc1881dfcd2cb1592ab2abf55a17e31bed8c3ad8295c7b7d59f9244ff63d4c7dc317855cdcd9de2d5a4b0b4f477a9d1883618fccf38fad50fc35c08a79b4009b61917c6986c8dee4c7ad7df227924eb54ad6af74b009e6f80c632686c448a4a4d51057a2420793a8ff954d81718e0c30e987e3155488546d0181db48aa01d1e1229832d798ae7b8214ff78b3a26459e4adced528678637478e7ff2ca1ab613d64ddb4c8b48c63f513ca07b43d07d8ebf2de6396c06a86383486fbe37527848681e8e9f6f3018c2d4c9ad89ebdc71e3df8c374d6dc91e23d32241231e733c15a467d966d69707ddb8b106d0cfccc881c78f4e27f2ad073944a8027b97dddc5d2f96496be1ecd0da2f5f9b609a22224b5da0b5d68e5fe1d66da719a5bc5780dfab78197c837e1b5770d7ff60d11a7aa630911d51097063775482974d5fe6f558c2d4bde477edd9b4fb75795e4e33b49d4cf50181492a64919973d9c2e346c469b119fd18255df8f9255d03e50bbbd18cd8f5ea9d2ef922bde550db1851511863ffc467b0ab2c5ea04a0e484950135afe0170b61886f5f719fb97b16c8c00433368a8fcbd81aaa39dd1c499042de47afc4d4e228023b8d833f7805e682a55d279aa7df51f9f193c0ca4b3ca01281f6c6702097471fc18981d8ffffa257ebcb022a0944a11e881967b3dee833e7c9d1d19a15dd3b9981b73d2d68fa8fbc0b129fe5a58eccb748c8a8820876193fe1aa050b381a0d365902c09e86d5da2060816c380c9cc7901111c4284e55fc072af32bcbbf90e89c46e5a981b2d8219ee505f71130fbafb887b1dd889b327f1ff658aff1d65b68dbefe2cd0bb5d63e8505ca6d768e54d591925174cb651600071e2438cc7e5d55bba40be87426a05d7ccb45dfad4b3f3d73f5bbd3c8df37b6f6fac1a60a3e345348f6d8356c773bb3f887d9271caaa8caf8023a67984392bd952851826de70a71857264a4e605fd0716d8c3f14a814070c1866e9ec2dad6febea3f21098eb66060c7b4249d55013d6a0c2758871f515da734f4f48dc9d9ec5d3aaf54923eae87c6acedbca044399868fc03a6dd29a75d1a9b67a2ec83a3f714ec2c0718f94a4ebde5308e465cc1704ac0ed427433be2e44d21701e3e600dc49b62f79ad6e68d0fe5e3744070f4b4dc51d305b5f738269d6053ffd65eab040a9bc18e427be22d57ca89339aa9a0f385d285be3b88e23cce7e977dbaab3a13469fef5998f4c85b9d10401d428f4dc44a664ddcc1815ad99f1b719f5c2b702b8501e582bb00d96fe9fa29d607fb52d92669b3e2ad5a655641b2b14f1b505f7a11c7ce2ccf9a40eef026ec7e34bcf2eece9b27202b15e4d396d04216da0c36371af495bd7eea43667bfbc3271ae627378c06885a3441a7f943e664c95656cbbbe436a19e6d0ca0337bb30f18432f8c51d5a527f1734701e28d275604240db31f0a7d920d4db5a3cb7478a685943d081ebd25062408ffd03a548e1b2c1070b7ff66ca7b8b326b4e990f17cad898f9648f08edfb83fcae53b0288bbcedfa27ab3a710aad3427ca9a12c731db761df39b66331b597b02403c7a84d37956448d8707bdfe5665ece3e22cdd8d3e3ed07c68e0634a7e252c122143984609875f2449f068b4a6bdabaea9ca46fe5540a806cf5e1e1c81d371e14178d848cf4f6f6ac1d597707316ea2edcaff2640f5702a2cafec5261e580a1b7d0d165d0f4344aac200165d483696345b1c968237957a2177827edd02f40020612407cb686c9a4eb3c6fee2c86a41d71442a0a42a8fe83d440da0daffee3445fa58561b032eb2c62926bbe672f11ddd68f31f0ebcf8c62c870aada70aea9c6b5077dff23a11db3158625858a1d42b609e99ca65ecf88bf830e7ce530c8eb13580d02dfb2db3b39227369d97b8aa8e51135f33c371f62db0c53eb85d98b2218eef518e16c6c6f026a52916d7b852ed61fb936c9f0b49121053596bd0d100d3a77627b3bbf5aef1deabf1f3e573441a4a1d93538147145466518f22f8e7ff0a9b00556018ae8f5e82f48757e4a3007c35976af218bd5f3a69f439cf16777816c3ee48c9f9536b3627d1382d2646a7cc7f0547c56c76be6e48174b264660b9b62bbb4004ebb3e3c5ddc3570e875037136d36f39ea4f87665aaa59f1f2c4012f863ad83fb0f4a806309875ac74c3e716dc53b6ce84a4aa17b5d4ead7d62ed26745d8831311557e5a87efc8305154e8ac6cf03c7819a750afe553488a936ee26899481b913da86a3c1ba3198a2f19228d0c1e5effaf03c96e0e965998f619fb09dad5ce4f48960dade353ff92168205625b0c8918a5c004c957358d0bae0f415915a3192cdf50b1ba286419e37a4819af0f779428d7162d9cc20d11a9400e0eed9c69b778e1ff70c828181ab7156b79d012d51fcbdb2bd313d1df512776a707cba172b848b3506fdc62d0016763ea1f1dd1ee786c0d8b7789875af237dde9d46696d52db4f0aa81a94499ff0b60201ed156f42c00effd0f29f9a303343200e65c45b7c0c568799edb8d6b0de61e14290c122e0d2493ea62263f0879f850e54bcff4bc4ae4b490cd6d3806ff74ab4df51dc7b93a9a1a89540f1ab62301953a19eca3dc621331692c62cfbafef9b61a1d6424;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h3b691c9fdf49470a7df1546569604787b7f45b720c7cdea0371eec83909be2400bff053dd717abc514cbf858e694816b708da3d592f0047b20636314ae048d439703497a8c945c670b275215fbc1e1cdc591833bc87071774400d0982118a265893fd21b0f152876390f4bedcda4929081e8782967fa92a448234fb6f9dd26f9494013e027668e6ee5952f29a47100c7ed57b25d52ac82114b71729aa229bb3676fb7e35aa1b07667482e9c86e4b1223cc64c66b6fda77ef359175b49895a618eb14127d966f83dbc2a60d45379872a317701c33c4d46f369d5176539d469bf02142ca9a682d31d6b6ddad815e4c2739a59ce1542ff17f19532a7c492afe7d597a12f8a458a60a9ab3696492c701de27a65d7053108f20e6af7841c9333d199c68c6d5e6ee2d4aba3970fb5839235d6b7f91c774f36a38adc8a361afa63106777b39c26625c1d7d286f84a464f8bd87f432e01c3b41ddc087303befc67f6406a3ee5997ca5c707ed298c7e685641097335ba6a7f7d7a6d95241814584f41e0cba266d39529eab28defd7323b5512755af967f116bd3a25353f5d9ceebeb4d5e96c93401d6475bdef586af5d560f4dbc0dbeb04ece4613cd30fce0312c0f324ace41dd2c2db09040236ce47829708597402c49b0fa490f6c7b60596669f45c2d40f9731a58440c7806b8922b51efdebddccd68134fed36f49190df8cec440fae779ed07d173e8919ce0769c12194cd2fc4bac575a33fea5379939649bc5f72a4bbb932154d3f2f7fec54b0dc863b6a1dca8e1cf6bc581292a4b3110a972a1657d46da8f5d2350ca2f98fe72e147bda01ec9fe6afb4dd68a1c6c0169a8e3b3b0137e8b042a2014caf56d970464386c94b106d7c948dcd5ea4f7854aed08bba03cfc7d16a0ef9e5287b7a2f87877d6dec9d3935bceca48c392f5835461294d3ded530e0c2f2d07075827130204303aae538d7178a455425bf7382ade49b419aa76165b454cd0590367411dd82ba67256616e485818164f6ad1d960bf9e47669281a7d47dd5cbd42f834b95de04b69dbf47f7565d0f34af9dafd15526d9899ac10081dbb411cc14a2b86b15790138b8e190d20f04c325575a7a52a95a2ba3ab9da9a99cc4a1125382686e8cf2d93fd7cab91a125ac3630d2856cf790777630417d6833e8a865aca7bf3f7f2f4c3f2946af78874c1249d6b46e3921999aed328e36a307a3dcd18df95b07a0e2675c2e620412434a5048b76a738131c45701e75b80eee4429f0d5fd393298e284e12caf1036e262b9bdd9a123ac6908f854d962bea7a15feaaa8cf0becad5361ae2581ad809110173b2423129b1be4a9fbce0b62a13a9fd6fb64ff862f2ec95e52a2c3440d0b0f970bcba2c0eec24ef35ae9127a60b4d2d3373b1503a3ee7d86fd2d14c5dba983ce683f04f21e686a7e696df839816d894cfd081931b1626dc22ded72707fa59ee84bcaea2f1d584d275a82c4fdee4df14330f3c4df2187c8200f5b97b226f5f286dbe46744e95b4ea59a7190ab44ae3ba31d79c6fea03b3ff31ffb0478fe56ea6548d104b2c88d0fceb7d0e6bd51fb938dd11c290175c78bab3f2076a16dab22b25493b934c90c607eaa049dd4b366f4a50344466015595ed97f39559c627f64c001fb16eb9c0d967789b8251ee34adbaa8f2f5c2c5aa3ffb9d513847b6c443a9c6abe7f30d8eeab198d493fa3fa558ec5dc0e3586bad28396d0bd36593c503761a95ec8652095e64abe4c3c4c202a93a9e735272a1edbb5ea8cb98628fd78c0213c881c1a198050797d1fb7599e15d9af4d9105a260cb9f68ae0eb909a5b558487e7bd3002cc70e9b24fdabb3d809fcf641df927963c2e195656e390e7e96461b8b17f61422862a89b43fdbbc6009480f3153d504f3b2478e22545d0b57e153c4c220c4edf0beea859191f9332b1b789ba523abd3980d570739cba5d2c8b15fc1f39d2414d673d9db44223c4824eb8b61c88f88ee3deede04cc5c1da1baf62507c8001d3eb515c28869c2037cc8e7a6b10369e5b3db437776f8a544e42cee31c1bf495fc704ae1aa966419f7880d9894615aeabdc9e7a3d78a5c48a7ab9b87361091fd6e1e178e8ed9b201ff8e381dd546aed030e8d21fcc520f526121b02f454cb314b8b5dfc8828a6ae33c0914576bacd0934c1ea8af37f00c0322da01e7c57cc42d327c2c407b3e234099a1603e0f4b933c5a4a12c9c707d0e2426fd286ff64237461a060024e8cc1ef7d4c6390c23d9594bd3891de152687e22f66dbca05b401e6b2283953a8badc8203b4183b262785a62fa03e47f1a631729bfbae754775e3a22e7c8d14ed4a63c19dd19c7a7222cfc42654b193914dbe7d48055c846bfac275469570ff39e7dd92440e5271ab0d8c4ca51a0a1830170287d3f1fbec46d6bd42a7f76921da0acc09a8bc7943079d98aa3ed83d18d0d7b7fdfde43b2a737f82cda8dbc76d049b0be324d31a7d7dd77a48bcb300bd4a4c5fbbd8e5d7c197fc5230984e2af06e17d336f7d6e3c1f7bdea966679f3debde69c52e4dc2ef02d32f455cb8ca06059e4f998f45cdbd0c93d84f3c0ad337dce916fbeda874525bd043aba0ebddb15cd32011c424806b38dc007f1142c9c2ec0da30c14967b9eaeeaa1c2aebc4a5708c485bb5caf1beb33a8c9d834bd72b00ae4a7544ef4d2d01430efc55af4330f45c3228f7efcd36a00de279d1ea0c88b35075ef5fff697fefa446e226c1406ad3d4902e83fb2107dfd0d4d3b198789b2bd849da9fc04fea16686e4927d41ab49d31252b92fcb5de6dce31b0a222615b5d678e67b0a193dea0484e76fa1f5503e1f9cc97316ebf26bf70262a726fe00d12e4c724291800888267b0264e3fa09ad66004799e3e2bc38687ab787cc07d21048efd1edf5ddae19fca17069c214f323cfd998ec9065b7e78237a891144912d32d998920a335052e478e6e9de9c5ad003c16b097f47191f6a74e3d752b2d992250b66556492acdcc48e23e1b9fc7cb625728db537d729f77d065e2b8062aae0b318339e749a136eff922e28c72749a3adab6b2eba943e46eaae28fbcf5c95497c9559505043b6d7bb8d42ae8b9a1e1a4408fd932dbc7c0720124c70532a003b26bc65a79c853148e14012767a7d4b417d9d7bbc521b8f407ce42ec3d650441763bbfc749dd6001d90b7c2fd0da68c93aee05b2eee5bdc808d973526f268c2b9eacc48f96233a7a266e23ab9df8eea3d6244b54d921d311f53d73c57b01f9e18bea39bd83b76867651031f3a3cb5ac4788ac7408ff8ad1fc15e83becb1af5aabdc3042b5d5b06dcef9f8d41e844e57931bb48498358505efea4c1818fdedce3c20f246a6872d8978c51ff79962db83d6393efab5e1e2c949a597b3b86b8b895dbaeeed37a2482f76f620a655d8c16002339b0fc7c5e944986dfa826082633c18d81c72f9e7a5e8330eb2507cc94fc52a08c980b7c855975e5da6607b0137024bdda3805e43535d44b76a429693d97c6fc342a2716c892660ad1cc99ff97fb33dac06bf8f9b301a53e838fcf20a2279c4db2b9ad8b342a1869c6a1d26be046d47b3454d3c0c6da199e898ceb5daf789f580f733c33b7deefb63f7e89860f9584b9786d5a4afe03626a7ee11de228d7954a58a26d77fd7bc9d5dbbf6883290326a7147b2a89f870a36fa3e801f8cea2159b62d8d79056ccd9205058e30a046d1a36de2b8438eaf98f599ee4e9196a6e09f6585e43daa8171a32100cd3db809a4a63a5a6a329e73e8330f59a4af76d58faed736465be003a3cfd40bad3acdad1172ef358ab8875c3a615c99f9d9f2cc4d6316b82d0a4942b0998c1bf5e39fd3402a3dea5034accc4ab71f443439285a2bbec1961b29941510aa574730e7eda9bee58ef591dc01f8c4ae325f8506dc102443ee8840c6e7ef713a7103a06dfbfa269a4feaa1d60649cea7d00333f9cd57fcdb6d1d9a8b195eb95a69320f0802e4a89fbb5a3157c82c78e411b48b3725bbbd5b49e4987bbbb0809accff06fc463d0c4eefd163681dd362ffaa82a89e9556bf6b33ebcb1b02a97f3c190ec7c144e32799f5c86582af482ecf59597b6c5863a0b57f4f9b8a04016afdd9f2ab88d2e6259928f29da98c78a0883dd8102c49464d82e62fb9662f1f86ba1fc7f66bc2bb0ce97ad4d06defec028f070303741304567bfdffc4d736b0bbc4996293ae2f86832ca3dfc6200bb31e53c96fc9979a0bbb21f89f668a86c5a00ec4fef4ba6a004d5ab96e416349529375847439eca108cdcc45b69a0c7aa4cad5d147f3d7a351b705e82962a83e472ed35386a60f11654e356ed2d565413d846ed398cfb081ac67f1f0faec83fb7e72f0f2391d046e4758d08e380ce85b77c3542d2b48d0511415cfcf9256b4677c19cf2dd56756ee5470fbceb803a9c1443004fcbb16946b4531184e0f20281a43ba407b1b30ce9b18a95c53bf53e9a323212dbc75c517f624f2592ad41fb2e4a79b194c54519952864ecaba99e2e2ea8345a4f7629d828ac4de7a1217ee3a757663d90e2ec786ce2bb8ed657d135c49310c0cea01ab0123197039e9d0e1043cad8ef103d96051919b54be641d196f672aba88d2a747db7399b21c0aef76d0ee5ddd08476ee541a70e642ec13ceb658edf792c9345c6498296b97925829695499e4256a5ef905b4ef7023bf724f6d0887335a781cb6ffc33f227f18dd09165b0ebfd7611ef714a1f7e74f1d81f0044a7e7d63d379bde9e4b1b7d93920110c1587c6b2035b2b30927a0375281175da4957aa2aa91eda1a7cf7b68f1fa7a6ffb10b9122006e3c5fce89e003ce7b71733f5fa4de242eb72fcd60b597d225c01e5ccea1ecaf2cec4087e780550c7f320116bd4822949bbc43138defcbf309d645c64d7af082a0770d0f0bf6a5e834ffcd307e5d78d2cea048660fef7686611c421b3a1afca7d981de0ef9be755f939baec97f5ca9676ba4afc04b1cf52cb873938878449852bd8eaf35abbeddccb6984c5352fe6e2bc055e813643a22890183c93a45ccc143041700f40aa4a87274f0f96c457b523675695b5c1ecbf4a869b4a154f7952fd71437ea000cc9b0a828854bb9de89168c64fb6b56ffad1cca25384ffb1798ac0b40805d11ca4bfd1493b2cae76de0a1ec3225789a7ac082f104ddbb332a8badc8b6c146745c4d80db5bb00dfbefce522dee768c3174370d8707004f43bd59cdb044ad36a2370e070f129aac39e872c3efaa898d8286cf30363c592a29b7392e87f82e7c428f2ea8f4e177d4321c79912fb8668b2189af6f31613c192733cb338e9093d120abd7a82e69de20d0acb20f327fc6af0de49aad9714f901e15fe2a3befdc34a673fd69e77d707b89a5ab1bdce4fbd010b07a88a2b1ca07f70ac6e1e6a35f326a179861a26771363c5b50a57e0d83a7ae55a5b1db886117a9d0ed4fe5874ec87447d78e7577e78ef6d1a289fc2e1acd5326d711b13b5095f5ea05d3bcf47ad89db883247dc6920d0321b88cc211136cdaa693af3a854d90a761a4c8f57dc1dd376ad8fa122f8065adb7d91b533d0691c524a941bd70c0a348fed76fc69046d965a7c268f266148448cef9903ed4147c299bcf066802fec217c949dfa8b03ee89d87813a2cb9336a73074e84ac7bce576c29f90bc207c902f9a9223f70777e93b9079e2a632d2014ab591dcbef6244787ee0016170571563d5934ae81f039c7a03988ecff5a4c19b50b9469fe19ce52180cffe670fc7a911bdeae3bb3d414c37ba55f80d2721977a891657df693;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h840d139ac5423a6e0f8cc618958b227b339e2219b1705d0c4814daff2cf30cdc7f556c029bdd56109e55efcd32ffd24d1a8f24c9de724c8e2a77e287a503ed4e97d3525cd7bf20b384f1a51fa55d40d1b789139651e49b6c19e54129754b42a87e9cb9e14095598a7334a342270ba7c26d224f9f501caf458e72209e352e06f6f3e32468b301dd7e7387b04ea326f5f982344693bb099e357c78f9daa6b8e5a4a0b9bd7cdd94bf355524cef666ba1da7c4e5e0242822ee793f18287d3afe41a4eec9a947ab3beba2665033f801bbeb594f9adaa3271e0e0e6985f1b84891d5176e6fe61768b7fb08074fd9fd00dfe1d18ed52518b5bff92619da83295af85f6d2480bba95b3cbcf099d236bfb3b97f9673c0250bdfb3a89366a9a5d8dabf91ba20bbc7fffa4c4dcf61bea244fcfec0cf4569611e767221da17310b422f94fa6110f93b9b33d9cabf410fb21e0b9a3fe6f046290bccbfd8c9e87f7d38ceb09f4b13c07c5f2641b134f76a913a7ab9cc85e8fe39e3444d1a223de6f1ab60b0f37cbe9d62be29b20b2233944f5c5fbd8e424d54ceaf9076e92109c107b3ddbafb0d0bd92131a83d3543025e0c9d833a0db2e4faf696984474648ab7a7a6004b8ad4c762a232c23dc754b62e5021033dc879de543625ad893bce737c460e48e6a0b01f45684fc10c5e849cf442b7eb313f037710325fe7a4cef412edc7dc7ed2dd1385b880c164635b97c25119d5138c9321748dd5234d9803aa2d98ee260d03a7e23d7063e16313f91eaf1736aabf786d601c20ff2cc05642399b8f7e93260313f7a70aaf044aeeab19dee78528a39c87eef3484c89feb4533e2ee0e61f0a7dc69959eb01c4828acc48c7274b3cd68b8e43ad9ea5d7415bcaa2c04217952f19809d2e2ce588bd99f40b66955a833f39dd60276c3538d0a4617d027687f3cd80d9bb228d4930afdb6f93c079f57efdf16be8123e5ea4b967c61253730cdfede2c35a1de252edcf43d26f8a7c718332faf80d26309efdaf8c8724ee4f61a4d302dfed7b2071f2c771e9f7ed7acdca90b357d6e45eee391778de5958a8a891522c541b2b5f0f6c90c1cd73366066907f5242e6340faaaa25b954fb6987ceeb7435bdcdda0ebafbc3cb12379d099d17aea2e8cf174e898908c472f0d5c23d28eb188abf5814cfa6f5b5b04f09dcb3cb984662306016cc1b1b70140ea7b972a5860813ba36a546bb75e1ebd09967422d1b74d0b56993b0cff928c9ed6b6caeb11d17d9ed18ca73865b83b97aee34e321ea8c1672be53ab8c7f8ca2038af912eaf1e860a1e1cbaf6ca0478790b761e20822f0b0db49665be98e86e9f6c779338a9ad60679ee29c1154db1fc0b9db6d9b2ac22bf2aaaf555a7ae339a2415cdef3eec4cdff65217df20a56b50e27534a2876087712ddf5eb5c2f27de1d720703e92017a0210f3892090d41231792aee910f89d7a4b5d3f967ad164cd7e1498cd249261bce1ed27462a762d2c23479e00cb82dc4c8a2bde0b5f1dde907135d96b08beb063620481c18d63a6625c39a8a801081d131aa07bb7e307c2a3a0f5edc22760eb0d143f6dd24afd34e1c16bce3e662decce090509a29a523daf2bd9807cfc5909a587b92028771b96307614d495d483a824e908c1845a97a3d148799eea1aca23a8514f4bf77f7caa5215c7dc753c4e88a2f945923d45c9017754c175993fb6cc85db49abc9eb8b100cbf6db92e452154084b4947a604bf3ef7e2711713156af2aba28138996854690688dea02d7d70a7e97fbab331662decddbe36d0335186fc2f23841237158215cef6df3d3cfb67dad5cf7a62952fd9ee6ff90bb101d891a7caa957ef97c0f6780b141f26c8d2ae429b1487346823c5005b3d3807be8a7cbe6e4e7f86ba3f61d248725e06eecaaa3db04cbe3586bee9135119cb27c9b12ed5500a82c76101ad45321f6db73d8dcacca508ed83fd14c64fbad68aab2ce5b6ee8b67e980753f44dbfa21d4f2e3bf59acce6d9ab213a90bde95786e5e33d5be220b030d837f14ac3e2224d2394e0d3d3d220951ad3f90110b2a6af7d065f1379e8075662459f73422851ef23d111eb96691989915a12ebf4637bfbd2f7020efb8db998ff72ccc5a67937e1ccfba577d70c43bb1023378f149568a7c8e07fc3a3e2a102c28ac66d9a3adf6c9b205b8d175e108c86e4a3fd5dd3396efecdeb40ac7114d69a36e5f46d91328b35335ccb5ae9597d5f9b0fa00327aba203468111d3c0048fa996a630af631d2ade532322204c03956b5c92babf50519674790450e95967f80a3895f24e017c95008ca208589111348bf292b35c1da3f5d00ea119efbcb2e28738bc485aa809f14ba16cc5db89a24532250e0763dba29dfe285834573770215b2294d38ad62edeb4aa29d1eda0b9fac8164be40f2e9ba9ae7e5721c3d5da69fd853a03b8f1da239d8a67dee045b71774d4114824ce2915feb6f653afa5726a5c3011cd55796c1ef782c6e7638670c4f408e76807b7a3891ea591d09189307ea0e5b7a412a5ab4782b76c0cec1155eb772c6d5b8281593faebf5e799f8ef3e6c33b5ede45a84e9e474ba45a1e64bedcbf20eb7886d1e3111bf3124d958be0b4237d1289c79ce042a79f26d785ebe123319b1a44c9bce159243258debf2cba097c208ee966446f59c81049d408d5d7d64963dc32dac39021a1f2dcc07c2fa9c59f5f632d6f99e5538ce3823761788a9d05342daf546fda19feb51ffded396535dd06c6006a9fc15aec7eca285e7c0fba471e0726ad2887923c3fd5b40a270595ec29a92fbede9158dcfcae80430b6f813a718d85f9165ad4baf0767a6c8ff72da1c70b28e080a1df68b5024c65b107f1780fb74391a7aecc1071a91d770721354afcd86b3d1b3addd30b4ba933f707d802f610d73656a4920eabb37b84d366dfa7613489eca7234c90a6c7d6b3a5e74bb8768abdaaa0d19e95dc4e4f774bc19b75c4908fc0bcc5b45ba2152c25f0c603ffa86b0db2aedb6e5c6fc40416a813f3d1a123ccb454c0d967be7234ea79ecf6c2df3809bc4910146f395f5da3910ef2d6fc09d489fd46b81ef86eefd93c76575129f6be0e488872db7163518d0d7976a298f34fb482cafd4c6f001ddf58db4a6deb91794dec1fe3ad22958da1e0a5b9fc448c6131036dbf9a70a51ac530d2192e463c23f059bad6c1ff0fd2eab5f1d4568f0c975695a0697b3e99101aac1a6d0b7606c1b2641411c5b2f7e25e82676a0c7a16733cfb10362835e6b9b7bedb916a927345c885cd8f5090cfb96946f3bccac509ca48143a84e0a9dead658509688af2fdbf07775b6d984b89203cfbdf8935d3d939a68b29b56a8e71b6fd38e953cb4f673a4dd255365cef483a40929937283f5b0e850c28a6b9cf6434a3708b9ede0f4b62b1e4e27ad10d49d7cb7361d816b5cd760a67585b3a792d1b59b34ef5ba463f225a358e7acfe3cd00004b74ef3ac55c54b246c7a7daaa5902f6a944127c7fa1729e581748651eef01e04a4c82f86502d415ee6ecc664cbe09581c53cca94daccf924c11651382c712d0bc70dd71d4bddb49789d403a4b155f62a0bf65e3dc517f8354d7ae40ca3411356a235ddff6a1f064991a23c8bf7e380cbcc49f664543e201c3f632a79fd98730cabb34fb7e703922d7eda9d2f98f236a9fcd076a5f64765f5ae22845eadb7bee9a3415630d341974c9da1aea0e1a36ac3dea035d4393ca89201ac0415c04d00f6eaf58de9328055bf913525b5c518b02cf43ca0a597fd608287ac8e2f2a17cb7ff80a90c77cc795a7ce14d6c3e37f057fdeb3996a52a99d66cc8b004cb97f3e75f249a8a4d39dfac7ded473e155ed2ed495da198a512cbe5a260b72c4d2e13aef9f7cc4e5d1ab757eb00eeea92db685396beb569cf923d714823ce003614df4ef144f379b334fc6f71af18dc05de298193ec721719dc64694ff0a2cd8924155430cb1c664b07aa4f96b0f41bc81ce6587684fe0e3b929fcf03264ea9837a92b8c7bea7b3184d40beb97d5c58831dc62419cd2e4a8b0472c58f89211894248028f41637e27d167f0ca5a4090accd46054d765477e10288dd2026fd6049a2803d90160cb1527278ac12cdce8a780c0792d2a8aa7c120d569e507b39c129c4b49f52272f5ee2d114d220f00e79e2862fc11beb9f5abd775b0ae7f67ea1c05d481f15836937f378cc585135a7d02cc99d0da988a8a940bc8534e0466abcb55fe6630588e9c85f1b440e5fca384f34f7a90c04609613f22c8cdcc01ad6b1edd6d0d239f424caefd9ff3a6d4dd7ee0a0d571c95a9b551c4d268f6029d8332b1f07855dd0504c74b39812603f82eb3e7ee5798cffed7ffa20e80ec2b86c8c7892713bf1fc3d72facb69e95415ab798c1ab6219b5501d341af908fe3376703da19c0ba662ed4a90f66188b74039ceae570ece67bf6b1afef1add0e5c6b4b1846ac5c00729c500f3ff17728e5166e53482be823097be5e50398d2da7c84334222f02287826d6cae08eb608dc17230612a48cbfa3aaaa386d8711979f7fa753b0e0e930e6b4ce0063ed1dceececcd57f640f34c36af566e8604415926c61b85900a244527746447b4582ec68fb521c80fc7fa1950e462589a92d1f5759d4a525c532a1a806f1957b24ba9fe7c20ba4ff1be64358e3a754f7f0d397612681322e5dd5b77e43669c93601dc138a17b916ac0cc131f38186faef5f1e549246ec60dac6c61f740138679c513c9521df59b5d4a3203aecdd37d9bb3f4c689848296a9656ad7dab728c07cc1b2e76bb73ebfba7e134d189ec17d18ae7f7cfe7bd6613489524060bf43cb757d2e78a80db4e8069631ae20392a17952037298e3c4bd9f01dfaa007aae69db484f512362c4b5ad3728204d26c2875284d3df9ce726047003a6d81f18a253f97a93797e92530e07bd158dca4f4ef6c1f05078025734d37a5f2c3bbb302c04fc1abe260c62744123c86469f2379982c36d536c0aaf85339a90a304453553d7162a9aa303a9db9435ebe0d164074fc54876b1a75cc3200bf03fc582c38eaff2009eadda9b08abb05e8fb4eb4622a79fd3e36753ab75783779c8ce25fb6805c2e1d5d13154ed7b1aa012fbfbeb8034f92afcd552a78bb542e788d30172088cba39a0d7fc16b912010617b54fd041251650f64c78d111472eb6b87ac5ca0252b713f9c1398aeb2ce23a6038677fdaa58cf2cfdd6d608e31f2e394582d9654047f5534f56c7641d29dd3eac90f553bde881625063a57a9049571fe1d57586128d642f1c3cf7a05df001cd564dc5fccf48be236a4a62f740729ea340e908081de52efb8ef0e2200d145001397cb37d79dd7d619efce03f4d612af9910f525b063cd5c674039957a3b9fb3d2857078991402a08a0d4a371c77442c3fd340c7ded0effb037efb8477d4929221abfd29ce24bc9102b80322aa2e58e28b0461546c7207fcb4814c9780d272659c5601a2f3a044b019b5abcb31a2d8a750a5d93e5f54a52575689b784fef4638ea5cd0e8eb53fef256b3dfdd231c8f7b7611f1c2a48d895b9d5671cb431a5eb65e966fc6d43c12fe738f82923d8ca77b87ac720d08034f872cd21f143a9ce4dc91099b3907cabcaf7e5aef4af193749f2a08d8adac13d286b377531f262978122c9b9aea53f12cd43cce9a088fa86a952df89981c92a2491728590b356cfa01c81b3e919a3aa7dadb7d71fe308ca21d237ff4ddb84868458b766cd30d352a16f86eb80a3e399405488d74cd024af335d35d9d592c264b002f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h7416fcc9c8b13900071d1e3075801e0ab9ee013e7d14ec93f5d35418d7962fedad77dbca91966c527db8869f4c34277d5fe036dc160ba8b77143c72e226e978ca1c5abc6edad0c6d6616b74b2ab38dc4b1fb2237481febf4e7e96c75378121ffc31e02c057c96af23a883fea262b2001ca55c3e51efe7b4d72ef654f64fd998023f29511cee7685027a7fe5cf8359d68362b8ba5687568e4fda166d51a0378dab622cf712792ab93f9ef5d66fe98886fc00af9e7cfa6d4570b4e135c236bbd827e2c8b796667cd27c52a9c4b40aef73a28d9e1509205158c462aa9225a2129ec0a5480d4de6dd2e154895324ed20d3248ee6c14d372f0b1bec343c14e565a7bb43e68e57a1b1d2fee240261b3299e7468cee64a5177e914b6e60497ec2af3aec9fd2f19759d31ff7adc7f40a56d92cf3710cf4a97a5e10efb8315c812f82b469a165232fe28a6fd16053435fc39d080b7c6a7433e2a1a3d6f7a9b57d90a30bb0ecac51a23693078bb830d2bf4fa4c18eba5dd46050c7997e3ed87c764f069331d010e47e9d1d40dbd73bb749a334abcdceb6d7c33d91ae361b64234a18a09456e88c267a8caecd863927f81fbf9c109d84baecc72586f9b591b9b917a43828cab5381ff36b11723098e27b2d7b0243beeffa3bf1995b5f8188497eaf48e6f39ba4901541b67c98a057cda6d8f1a593f04f8beeeb5f955f4c42f1909f63fb73f59bdb428470e1763cd262a1505cbece5111cf3e6dc2b984226eb1dc3d7599968f6324debe45bce23f07f43f478bc65cf2ad0873037ee0842e28ca5ff2f090f2e4e7922ca1440264e4fcf487a0468f43bfc2abe9083b8e6e551c7cd15366bdbbc0fc06977d7040b26b50ce9b760ea146a5a0b22ab416d3e8e2374569ff442aeda141335b16d7e50b9e4a894fb126d468236ad8de2e0e7d78e464ed29b9cdd5da1d136423acd1b556fea9e2aa5b2abb565d16afd2e7a811bcd2cc092cfd4dee5038be7b19a7d4fbaa4d1fda61d82bd8975bc53e2c16cf0268ca8571442f74aedf4dbd1c2cdd83e7b364358529b3913d707840afe0ef9bf5f18b921a87628b2aa83481600803c9e8f64232fbbe0ea543f406dcbd56417359edb10a2ab61c934c21055d154ebc035be3e2293edd87437e7ba6756053386f21ffc40da82a8d35ed389b2200fe83f09735083731cbda7e3e5103270f50d75d3037823798aa5b210f25680e6436ec316e858264d5c6025e85747db8e0fb34e43107d5a041789e67ebff48d1b4e258d16c437aa5d1a76ea1752ec6c352f7f1cbd068c060c15aca16c00b337c7efffe14665f520bcb69d1b8fe26ba4020cb957c65e60904cdd21c446d2026ae7e6283c868f6c36b569fc34c1de27aa3e7dce2c390e04661fe94ce1a02a3bab45671e6106bc3ecb9cb78ae4a21aae69d0a11ac8c5df22a344ebdb0e2faacc68e985f49c2e2b546604cfe64bb5da4c9c9d257bb0f5eeeed776db57cea045aca6a0a32eda49604c2c73be3f9928483619a3364e960c07144869f517aac55b7d2277b3f0962f21b6b91dec497168ee01dea7788875f112435c1b6b71d98656dd3372ef3a99154cf214f686c05d1e76f23f5d30140bd21db427d24589229ae7d363165ee0d309badf871dc9267169899616e7c2f7d678dc6c4d487981e597f22afd494084750e4150fa38420b1d5b0dd7a1c9d9d86ee884a7d5090515803bcfb036e17dd1552f7dab5cd0705be3d65ad834cbd9d68f450da4ac24ff320b0dba676271f05a53f6daa8b13bc752058e0e680249a7c9b7feada523d0a1b0147c38ea0a0ea6146e2f0e52a12676c65342cbeeb6cb7a4261b4d5a37765323c4249b63f13275b168691c18c4c7de9b7b02797a5d79ea61c740bb2f319f69acc42bffcd6b69a8d143b7761bd848e5e752bc6995092a822092647dbf3026e63e6b61e8df3932e67fcd72effdae0879e234e35d89211d4209bbb384ce4c91148a0d71c789540f8e370e066054683dd033fd97ed4992b6c5fbbcd38703d722da741366e88e5b15a0143ce919623363c12f889697f72f6494463927ac5eb48cb8c3ff2f846f3144723c6f41f5b3d2670144b18b4d2466e83d33b2eadb42b63210751a8197ebb3853694753f8c4bb4478d60fc88a4079bb1bda81814166fa9c670b42a0db6994f78f8880e4296e512caa4b82f14bfd2019c99ad4b43bf524211acad6330d8714590d7e93dbbba6a8d3c4bf71d17036e91c7535fa94c1a0737990273a96b1093ad8c690ef1df693252a430772bc8c8674763bfa17df7a53c9dc008c4a100ea43c52c5bc6419b1fb41991b5075c688b73b6351228610b3fb1eff49336b5c12ee4def2c626906fe9d8c3425d0ba26079bdede16b20f4e51f772df46f85c9f32adf388b46834f8febe2226bfb9dcdf0eddaf66931f2f03816b1c2999ac247545ad41e48a6c67f880f0e3f86448eab099e041e8965e569fc2421774b355a9ae52d0464b9dd50f4bd0ade2bbe07a6eff300885053ab7e479b12710f8a70308a01aae3437e44a37fd5e2063a40a4744464a833f7edf832225c26ee7fd8bee9b2ffb9419de984929a5853fe2f90eb9f9ea62662606dafbb5e7192f63cccdc4fa582ef0c038b1a0a12c9891ec0867746e9d89449ee02d6cbd3ea7e2cd0ea4521e35c9400046117aadefcdd06963600d6c7772ae2b34c94c0ca2035f6623c43f681bc5759bbaeea19e7bdaac0198400d73fff5ac520549f433d6c87fd77facc1064856595e56d152b62e2306a4d3305ee079811b5e97592701d85220384b81fcc1ccc8215c3f056bf1716b6708cf2c59db9823cf0221fd24d4b49b62e895da9b27cefb0d01d49810e01fd39b446c0e6f9182828d75daa422d468fce091bc053a60d8d94753b5b525a1051aae8009028a72ee17634dbade8c529730888bffcf50ad9b0122cadebbf3ff5c525cdaf37889ba43c8796546af7b14b548c89b856bee5b7e32774284c192c918e809a3217f3ab2ad853174b93ec9e58c0fdad4d2af0814726c27d7ecdb18570e34fb7a0ed2bc56d58b661a5b86a1c8481d99cf213e5f2b24fcf206891a204e150b951551d98c48dd1e52876c775881d1520a8d91d8f15fe0ae093aada04acae30f1c3a0dfaecddc94a559007a70ee1669e0a3fea8881d5b0cf4cb86a5445663a5c3b988e933c53d5bf240f6120e6e63326fd158d5b98a7b4ff9eecfa5a016f1d72f511175b7f3615c5244e02821917246bf6afcd95f6d53d2864983fbde6f2cc40307e443014d0d5aa3418ec4733e37de1c89c1b38c6c6a1ed1648f4bdd66429fd736e4ab704c99f351989b7d46ccb7b3b5a8baab1204385adc384102492702c17ac20663c8c3e0259e2c8ca12edd147bb109a7f167b3a65dfe8fbda72182b851935f8e4c5f9c992e572e042e5b7df9dbf1f26850262d532704e76872bfe107ba9571340b92ca655545326f0d53a1cd98d11a64c6f8666d16fb3cb282dc47a6beff915e28c56316e75de08e1327f7b5d0d38eddaa2f0c0aca312f22f2a84e2a9d1cefc16b9209c49b7ea753db16a3abb72f8b964c545ac2b721cf6d7c7392c9a64a89d171ee6a57cac68b83bd034e934ec00ffe4eb0a6ae80396c0856fe691771d3eb3e3db1224c1b41a336d1e77ef83589d090a1d1fd6073048281f198453b28ec58c21f707e9ffe26fd99e6f7c315f831cc99605a1d072f9857001c4c595f6ddb467b5145a247379cc2bd7cac3886aef3fa1bfe6eed52ad237ba8d186855653258a895d4b897ae6e8b1fe2c27405ac7344d7d903237fd4928b85378f310e6c323fda9cad013760f55ea0c8ecd56ecf81722ae8a5c98e1c9f91b486484822fc97d5e4789582daade1935d46cf152b51f1e6a5ad170e7b8ce87bde19e9fcb47c4d71aecc1f6e64213bbeb2142f7b1518bef36488833d6314297fedd1f3860994d5c8d0cfb8d1c825e223305c7382b8c67de026f65ee1a84766de6c3c52fb32375f3f4565e1b3ab9708f37f13d925ace1a3e1e80f6b852819809a3e1507479b8d2edbe9e63eed72176daf5f804dd3a511d806adf1758be5c8d467e65f6979f8b419c2cb211bb2ece77345a2dac4e315d6e7326af6f69fb2d9337106bfe890d8219023e407e9f176f17b18b052217656c44a33f514db6b2a1765ac5d9e9d31eeb6b41d6a47b53009f9c6de1027fb829298725f2996e6290880f4d0b748ceae78190376612425521a57c43845b97a5fe729312bf714ce75d2e5145fcf576068f8045a5ae14d973266b46f531c2cdecc359f105e30810456cb2f8590d7e64790907e4e7e861770c91f5bf4b2462e7265691a4724d50beb339ce0c49b76021614a782374f37521abbefc12cf33c90e2b22179e7f9828fa61e878045fd08b02713f972159aa05397db429ab57a1a1487486d1f2dc6517e9b47f37111d4c2e093403cbcb26b7b589ef2947a9bf3238e414c571890aaa80b6feecf00b7dd905ccd6c0e972e7269dc1cb5b55085d7c4eb65de26c5be5b2046ba840a3ec0ab51b689b5576d6c4a1055a79ad9158ee09f69fccb1db8a9287ed007272a1a350f6c81a34b0ee0633dce9ba5a33dae801c0b11ea14e0670ade7038c214b9ead9cfba58ff66b43dee3148dec6c701338d4f01e6505a2a0b1e88c67fe4838cacdc57d1912d89b27edee6065bdc16941c6ca24f0d3976dc305c45146131debf2e813a0f0973d20740d90b8a740dc468147ae621c1a42738b652064615e12fd1d7efe1ee7604ccd69bc24a5e255843cf520d7a66cf2298be4009d6cace8a607053a511f442bd00f0e6ed69d6d4f95a368474252ee7317b25bf7c52973fcf1f6f398cd78a24dbd9d93b69ab74339e27556f2dc106fb1582c4c0831f497f44b3b93de956a18bca60bd6703a802ea1e814f6567e8a79aaf2574f29637078064b677be96094deee368abf32b80d5a451ae939cfeaf3fb40f8d5ed493b1efd2ef16fa00baaf44a73eb5bb37216bd4602cb0020c7ed609c93b864c71a7ef3c1b36843523205f904efe14356be3ad66b5ffcc7c8e75472d9885f847ac9eda290a87d7992ee42eef6d4abac682ed5b33cf3f576be1ba7bd2cebf396cfd2465461992e2b0ff2bccb449d4b5c97767d67e2e81800935807cbc61089bf3febad7c8927527b35661116a1bf2eb9d1d724e8133429fc4c6376bb4b64e914409188de51319dfb0b98c1fd1e11e0f26a57db776017423f4d4d21ff494adda5b5eb4b290e9694b550c9c4d57d909ce6f01f5959cce68aca616df484fd43d0f070acb3113ec0163bcb018b7ea5da55d388e4416807302b117ef0fc92733ec20760c2cdc9518a3ca078962f1fffe78bc05d63477b0b1abbbdd50db1a5cc0a49c485fd3914d609dca0a4afbd70d67265718be9c5757639b82f9b5f4b7b5f2cc5417802f1b6639f68371019c4fc247e93a4fc31cf9630d0e63cb4b071011af9b9bf835adeb8a7cab7c820b118ed46ee8547ed4f11dc36b3670b3d2183c5e10b707523db63af8085363b0fa403c6049ab8c818e807741e8701fb92675f413a9191c3f0916e4fb263a638b2b519dc702a2d0ead55e0bbb4c38ad91d25ae003e5783dcec0bff4d7f6b08c4550973e8fe3ab253cdb6d9e050f9ac05ec31aeb686a3529d275cc160cb13d8d4c7edf8503f14d259c5afa4286d674cc8824b0c1d7f74f0502781be54b3933dc19a4fe218f7a980aebdf83ae23089135a3fc4c2d5e1e109a829efc91e330f2e7be2bd90d6c60f81f65fb0d528ea3a0c45230bc1d5455d6788a951e7c526d799c8744e99a868;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h27601e69527c1f073740f06db9141194bd5e7bc1308e9f284a672ebacc5dd69f893a05187fffc458de5279380dc1a295fca1ab7bae76854818e015e5c8f5e6b60fd5487cad8adbb51247fa4be907b8002d7d5ce98cd8ed3ed2d8088402b6b1e7bcb2d1f1dd754b42a0c8ae5db6cb2c78b88483a28645526595bf2b9508d28834185469e135e4feb55fd4348dc28f86b260e62dc226c28b3e77a6d5ba045c4034faeb46ec01b72693c7df735714d02ba5067ad31a3eed2390418768b52d893066c06fab666da3a0c70fd9157a3492f9299917adb0e42499db8671e6b3d4a655ef4d6dbdf4e3657f2f4ffa07c3c47c6cef11e98a9a94bc05f7396de452a2a8ce61c9517f4b4712b0488096fa48ef398f7b58d12a5453d4721f0a805fb103ac725c9eb3511f3e7c60f90bca64362b69d0d5c9d435faa3c260f6bdc8c076ace6e0d270e84b876340328f6b5d9125aae5143416d287e405e7a04c51da92dbe97a4421d30344f8e7261a20281193a2db353d642eaa12b8183f2d00ed37308de1ed18003fe05ffe52990c2fad0bfa9a9fe81a608b4bc91a8491a445776f43d90a1cbe80241899b809390aeb079a104532dfb00320b558a1c8b0f8eecc0ff3a17ae6890f53b7cfd1e05773401ad3e5c8e1b3d8ed8b28a67004199c5e090d0a6696c74735539547112902fe25c53c1baa51e29d9e7fa4311bdcb0f98a6c3cfd5341a4e9bbe1b75bbdfd17a6feb98ce5cbdb85eca279d0929f427d19aae4005f36a5ff2f9070192698b141e091be40ad896cdadbe5e48da9ae034f049df76d349b3348203e9baa20459e649dc6c3a666da74e63701e484286732ecf8681a204781779cce0cd46e7c98def9fc13938bb003609d19bcd7be4ce4e40e82f6d1cedc135180ac9be16730c446b4189a8869cea034d5c24d4e6561fc16400e764b160b6debd3af73223efbb7bb1dcefe084d4782fb4ca3d54796776879d236ca48637027f2820b996e99be6a66956134bf0d9f9dca340612bae8575e0d3b11e09d346a50c2862db8b412517d8177bacc813f4de2ce81396d19c385e49818e81551e0980eefeeb5f2a84906c746f5698a0556c2faf89ebf9cedeaab31d1464c4b1ca3951c8db938f98bded8aa492d68d15cf3acb3ba75415b450c0b51e729b9d7885cc94cd51ff3e8dc705fa12a283f94cdd83b822fed125d826d330e3b19dc75afafdaaf5e93c7e543159ce26d0baff7eceb85b21dd57e965c43885952371ef5d2f8476644aa5d5e98483de7f8ff59a99f33c120e459815637a52068bf7f7f14af04f60e761ad44f878cb0483888c348ea5d278f8eba53397ca2142b0ecd4d131356a00c3120fdddd7107ef705f2b7607fe45360eec3ca5ff21352603c75c7c5191681feb402f8127a4c4fbb51b508483a3b46c6b6918f0d4293d0fa02f41e3100b06ef50289ffec58cd8184654488ce5be0fa618a8aba8067ceabeb471c082d04f774384bb561defaada158499532697ed92aa44a938eef9789bdca3c71180d56cdaf40375ba852356a0e8957da9a24c83009389b0851b87cc8ef1af96cb601dd5c39c059d6a52a8f1b8fe9ca4da4818a7fbbb23ebf237dcef70a0efcb29f37c60c6b2c3b26bd837b5e1365c858ccfef886e9cd5e8bf351450ffd076a3531c1822ea1450358ee00d65ff54d4531cc055206280fadfb75591928bdc95ee1c2d88d0f1e4403d8cb4bc715e7fc658ff77d3e8c1c6dabdabd1fc0007bfac07e0b78e1f3529f52df84f08262b753bc9b12d09d3d55fce01d49e9512637ddaaa3437852b54af22c3472ef11ab437ce5917e9bd7b2a4136431caa2891152d3bc70f70090e6dafaced8dce6b92fd84510566d41678508fde034a3c106c348b811d74899f3da1ff3364674c00e6faf936c69d5fd261e056fb5429a27a1be65e5fe7216f412810bbe8035b25c019fd555d299e77e45804b9bdcfdcff9c8900740894f1248adc6c45cab1a2c8c6f2ee2e8d05d59af950bf0e93c2829581688edfd2970c13210d70a1c1a6c76296e927da57e45a57b65933d307dd7c47c9900c23a94da004c431a3d13b917f8beab87b8f231987708d71dc76754a7c7713a23ab6257ba41e72602e9db53f5a2493802e24fe191464c116ba13ca4452dff6afcca58977e21630c4f71bef7bc5d1661942adb276ed76f005bd57b58d0282d48069832bb40848080acc0fc37096438d5bba53b60b889af49477ae6fc1895634213e00b8e78bdc8810bda9593155a3cd4e435886331f50e9f2e325f99b7c639c65ba473229ec89f292f56c8aecc964d40fd88123a47fa06e4420ac14f4294e9d0ce2d9ff067be074c02bc14797857d3ad3af84b3797772b62bba1706e7d33798157bf0c2f9a40d01c6803a10098e59b4862166c941db08c6adf0a75d8943ad65f062bdd6de6af7783aee36fc0e25b8a477d99fb1fd1dbe87d2e09a2b08f0304f33df09dcfe24f4554e12e8a5436080d91a34d857afd319dbd6f70fba0ec1375717e7de1860e29d47de67f49f772058a71008ec1dbe6a290e575eaa73a88709a66ba1bfad0f5c1840f36cebe6beb12f41f2e948d79ebd11e4d6c1b2fc68c9b0e5ee33f5b7026724b467f11d3cec54ab7a4c81fd2105dd9b14b7cf665000a50b00c578279fb5dc1c389644250e3d1ad57296d96e087310e47bb0020ba15fca796632b68eb3a079e78778c532fff28ddeb153a45126af43c4128493e372ecadfed1708872c16478daf1486b94ad5fc6fef9ce17ab720d08cdc9be13fd5bbc360d6e8be6bb0fdd4d900d0d9dbe8a641a6c7b24bf985f77d91b356d495a8ba6b87bd3c4be3ecd61813eaa3e4f200c4f9075b44e1b3c15f37b8852a368d986cf8f1a65dcbe8c3020234421f457c8646e7e2bc0f992caf5982bc644f1d0b338058accb19269f743a3397db765bdf9b1fde3548903eb8058d0dc33ffe3c6f07694713a3beabea01f8bdd5ea31d0ea14a29d3585cc2547f709b6b7fba1783d85ceb2d8e9bfdb6b4b1423512215d15a8d4a7d6fa76dff8d83fc05aab6eea2061a30fb2b161088d77cd94cd6ddc615ecc272f90c3cc477c640ca03bfc99c4238f1cd97f37e06b5f40a7709ce6b2605da5bd2d9a0a22b8ad2f79ad0958cc8b9d3d8fd06deba9a1913bba2665568a0e6d2809af1cdf925cca0326196b42c8d681b5fa879b5d340ec6307a5e826f1481a93d293b3968db5dca1da4d724b257d980bf8089be846af43466f55876d550031e934ff9cb59db0fa68dfea7edbeca5d1f582d0cded7513285bf9aff3ef0f630b4ac2072e271bf8cf2912d420db419b4f8ea27a94f7c75e7fac5b6420de4766dcf552d27e6a08ef8b7b26f7cb4c65a319ac71f5389ef54d58351d927ce545245d78726086f06ee4c6724a742f5c93427732d9ff814efff1afa1ee71563384c8dd102fcbef3982294550a4c3417c1d9275c7baa1af0180a886985e89118c8d35eb0e32a1e0bf6b71a8f49749ba786300a879aa4d4790bc7f482bc7d934c8d20ce623d12b87240300bdb68fb80906ee274fd7ef4ff491d10c14a6c492230f1ab8214f289784cb63531c769c2472018532915dcf51341d40151c4f9830910627f8867f16d1e841a5c942de254f527dd0a068d96f77afb8a3757d039e6838c920638e8b752ba5a193ef9ee1f7df4c06872a4047b66386f47bf60055941e84bbf98e2b94ab788b230f6c54483cee05bf378c06d63a35ee48ebc946f1ab9a3e4e2282591a662a195b3d750bb26f636fe12bb29a05f059c19be27c76b86cb86aa105e89569d77e7944902ca3fc35173deae228e3658dddfcec2bdfe65782ec4343798bbad92b2f39f6348f901eef57503c0a677acc6007b4d038fa596dd07d19349741bed1214b89a93ae7d509760c1023d42663fbfce5012e2ca2c437439e3f7f3f4f2b552aa0a0e981d03dfcc55990b23fe8029f03bfe8e68d31258bb63c6774bfdaa244701675d5354e8792794d1000fc09d1a33a7c3fcbb3f3c7c89f263da439ab6198d2a9d99848269cf05d9ee0d6476aa120d641fb428d71373e6cf8961ddabb28ae50d458f9553ad9a7994fe6c071f23600adea99c80486822c7efc1403a91f89c655895a46331dcfcebbde40460e1bcf08108abd4b06c3c43765a818f70da6af4517a5503a4309585469ce13b7acc1389763a8470fd48812d8d0ada5e593dc87dfcc191401b3830240d16cb8d453fde2b9ee4340f921516f19c317c3f238e851f8f5fd7836db08e962e14eead0360f58a290b5766f7d70eaf2d34d7411f68d665d2f9c88949e7edb1652be93826258e7ce353222f26401fe96573bc4c02c53e3e0e1809dfac95bfd7b07256637aceeec2fef2e85b6c445d0b8cd0ad6dd767816fa1faf793b96dab329aa7e27e6b24a31a5729de1850e4e1ca902bd83f15acfd07a590e4aee1b3f826a7a24ef0d7dee084f5d4be15dd5bb9249101dd1bea7d7fa9c8dee2733208f1eb02abef9db30d19dc9d6144645f9b3d2f76b726d7a61d7533a9d8aa3520ae31ef13c89e3c326c9fd995425039b741aa873bf30c9f5a7af47ddd3c866e70be8ef85c06f47f7b70c4872b32c5c65365de55c46193030ae0eab5c96c359e8228cd8e4f955451de267f913feab92330823c5f93e3ca63bd624ebad835faf50b74c501c18695967c6f73644db5f1b3714a2c3e2d1d31bfa5b60d699aa3d0379e6890798d9fc7b7d1eda9f019c2bc56549680b36bebd04929e4d9a0eb7965ba244ce96712169d64f59d6e4559e363ebba2d7141e24167e98ee33a5b974ef78b9c5f8ac372e4b4ce5f808785b781d364753e36fb6c11b50088270c6c5d9bf8538fee72ffbd9ae889797a52493ff33990a7e657aa95fdab83fd10195e2a938a4382b2c8976d192df4aad335dcd1bfe670a1759113e1035980e9402bebd6c47c1b772e558e15e90a9a448499f2b2cb388939d5f3f19fd94bf7776baa830ee81a52c2bb2ef98cb3ff8e5315a57f495aa597386702e75c15714fc8d2171a5733cea9e83f8a4ce0ff27e1a422434ffa6b2ed9ad79527a34570aa2a95ee110aa5fbc4f88bd45edb4f28586827f86f661d33eb49e153b862a8242911b4dc4d76154f50ad3b2e199852b0e67f75db7098575d94531a6ab6351aaa5483d08c59ceeb3393e53a2cbff6178707e4a432cabbcf2969cc2dee9674bb5e830556c1f31641527daecfaac19ae607ed64ec6ce5a8b7f2df50f56ae7c385a4b3298f78b0a372a2762ae4951b5300100a6bca51b0f7de422bdc9c750e3e662399a6cf59b85f97f5d13fb23f1f7a97d1c8ca9ae0b9487c792b09754f3127d6a42f9d2725ed256ef406d9087082438363c3ad4f88df314d34d0a42167cff37335418eb5c063ecc6113139b565f12bbd0cd9d0ffc95401bf78899339633899060c663692524cc63bd8dc10bd43565370e86edfddc9f11fa8d4f1a16bb11e45deed8715bc7f763ad18b3e0eea0e139c4a24a007376e86c25d5f9410ca075012a102dd2599c0db3dcfbcd1eded1a446887e5bc43dfa697f093a287bebf71420c5c8468e2c9bcc5ddb7eb9bc720697a3202c1d96d40c5d9d53ca611355e1e3f15e075a4e7edaab7a5264242db4125f371a4b81b51e18beebe133eceb578fd1910b18a4e41877111c5a4380364218666ac51e80e7fffba1691699e790a23a3fe5dec04281d4b098ddfdf7f419b69126a960c6c032f5b0725c9f96b7f638c9dfbe8b65133dbf8f70c67376df4848cddd5ecdc13af003ac9612e42ab561c1c7d4fdf2d2b6c763fe2e25b213ced1380;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hc03579ca7738cab5d717d3465dfd5623ac47279dd4b7a1538a0a7c5f7b01705180ea20c6dd072469cf92fa480674188a89a94d810748db403d897489a71d2ec2d673435a0371ee9d76f6fe117be47850a64ed96b16c2af9fa36534a028d0813ecb7b5ec73b250cd554512694b9505fb5852977a586ea239170ec8e48e051bbe1ed19f0d39953b5a13fcaf828c706c55f996d328a489595a4282919bcc02f5025aeace359f34c24d89bfd53b8528c786086b508f66585e69666983a3709c0441b32b6c81ecdde1e13bb6136d15cd7438e762d774d0e4637b4ffb9e8d25d728be1bab6eaff4cf8cf36cb29acf9eaf4af85d226aa3ed64462c7d757e0394cde00ff8330cf4b46d0fa67e938b9f1a0f45bc1da9cc322c315267196a6f8d77f9c5629524f3657d1b3e00af51e488d45fb2c1ce05c9dc072d3bec0df147e66bb7ef470625ed949ef7a6c1dde590849bac4207f603b63fb6734e03ea64ca8bcc771d2307a3c3ccf97a012ddef9c76f924cae7d5f9ad6b993dbf2c11d5da7c1bf61ab4a7be62e6a548842171cf49e80cd88fa956790e5bdbb00ca36a9a16c202a99970a40c443a3133fbdb7fd25f8bf15267c8c0af5d73a5d8163223608fd25273460fbae9ec00fa40fe984c8618bab4a93defcc4201746fed438b0021d845793f4c87a48737d135e29703d7bf661a3c49261479e321e3d70c6c15c4f5406391b99bc9d4da153ecb88bc53f2fb1aecc42f8d547b4e9cfd4ff338fa9a9aeb73a960ee997a93d90169c91f36b49879f42f63837cf4d0adcbaf984f2ca5cd4122450a4d692b63389b8c15c089bcbfda71ca086e9502f1d7e19d7fb85495731f4a54b763ba9f238535af46edf8877fd298b4f9d4a0ff4de01178767aae9a025b797ef4cfd02d6687225c138119243fc54e7764bdbe49a8f9c8cefc39cf0474c3be723ff9f4be4733ee5304e075ad61f60b0020e4dd8076e33a98044375d36ac15e5cb9b2d10b22f67696484cda0413bb23d995897a1da12d3cbadee015a2ecb44d99bc72332816e19a41f81ee3a3193cd741fac33d39e3c5a2270a7532ef5b1403cbd4a43f113aadf4edb44f5e05a8dd696aea7c4e2ad4e25d894e9d8b269f4b7d48af15841ebac536ea20fb09eccd1d656f2eb09cc4534dd71a21671ce0e2df3b35483eaa6758b3bf26c9facf52c4882cda9b6d6ad4ec44478ed61f5d121ac910e84e07806a22a4ca0a2b63179b5d36544eb61924b7a83b75bb5024712db661250b44df98b3936a0a3d61c3d585a00efeb266e9b73d05d29c6336df482d5fe915f2b037a7663c2696b0dbf390130354ee1b94b564cf67c431db9485d06255b07bfb0d7d18143b7735f26602f3ef92a07d5fc45c051509b7faa6a6c644be8382fbbfe084709c68c1e6a6303fac8940bff3f793ce5078fc146a72874549ed8bbcc7a28dbe07b23fee83d72d309b7fa328e4622d9dda8a31206aaa41534486d7c9c88d34563e6d586e146ef504cc3b7250df458c3de7848b8f26bdd498f94fbe35d64bce0eed1f7d8b028c69d8212a2dd3b1ad501f65d1521f0594d1b849a0118012ec895bf4840c38248b2e0d62a7758c18d300e108097b9ff3f413e911a7bc715516643b278b88210fef2abf299109c65114e992800e5b5b0feae1acaa206dbf034e806e551cf35c363239fe558c372798a39df096d943dfcaca91a09b1b17774c31490b210ce61835f971f5763b08092cc41f25a68c8d3eb2ffc799c896e6da3b74a6c68003a5dcedb90fc5583b37fe42436b62033c30929563626a2879a15c5097aafc1a39f79a44912da5207ac964a30c7e06291c89309c39f5087ff8f91caa009210bfc2706f6d71e00d19e02421e16a5ff926f0f37e341740994f7420bd5316694a5ab95edd60d141e95aabceebfd73ac4aa9aaa8da7ce513577c2ff735aad5226f7a139ee15e05d6f49c1f29e2fc7be692920b4b714588a10461e897eb566fb3e8e15edba4d1ad44f490654924dc572073817ade13fcfd816c5edcf88e034eeb05947a17fd9711bbf08e24b69b90a675f77f52d052c49b6aa12a9f66a8f9028198c8ca79a9714cfc1805526085501f3babba6b593120540fbd5913614410cd6529c14107e7933c0ea937981bbc8b2fea2a9ed8b6489cf96cd8758a96cc2e1ed55b378310214723108280a2a296550f49f873bb42af68c3eb91e47e88c0cc8ab86a392b61b1bb7138b04a17b775b5e4502a5f1e0de20f67c7e9287582315ca823629427245440ba9c7a8a07188a5697ccb25c17eff0f34d158fef86a39e35f295dcb6faf815774f4f4a18feaa47cf33f4afb5cfe24ba684f8e0c5568d4436b7b6a885fe22a73045899cea4bc98fd519eaec543585f5ffee5944772f1fbfce4df970bb13f989990dbe64b8b27fa9e40d94102cb974112b82b8c4a77a0ad88f6f3249baaa0218bebbdfcfea895d0ae67a66554e9eef2c215e7ed1bf0ca64a81a996e88de5a0b4d4cbf18f29811aaed71bd4e0056b28e80821006298feacb8ebe2e43806ef0ea5e2eb97ecab7052b176b939f4f4b85a53a486eda02fc3d6bb67137eac426f6848e221540f05cb2ff589ddac2b5d2b97a4c06d2181621c36be97ec1bdf7968d903d65aa5bdc07b2859180a065b9f427fa0ef4fe2cb281ebe8b05616f07103bb7ce301ae79edaeb37c79c23223267ec4da3a8ae00f805c468a048aa28063f9aa2ae7926de81c9eff9ba3ae1f5f4a3e9d3fb8f07375abd34640e1b988302714790d26290258c80d4002a697861607296b1b6d67e2b6dcade85dfeeffe6e8e999abf9dbb1b4d3fecf58aa633bea47c58f8c4533fb6d61a0dd26aacafd5d5e16af2a38eeaf7b83c722b5433c86aaca08be88d4abd70f22389bc3f800f3666b915e62fda97b9b9899f522edfe259fbccd36078b1d3a82ab2a6780a32b24fe64d925b98d9547e8bd525b8566e5cbfaf5535fd6ebc691a18215129bed550822f5f205c37c6644dd0c2c5e5392c7418ecccfe4953374eb34ec23b0d296cf8e26a98441b7c076a963de6f3a2786453edb18056be13b1216545a724d6b7279c88738592aeb9686838546b180070f8c052f59e36d687481a69e823e80f99d2f2e515a26f8fa71fb3aa37031258bbbb5a904cc3c4cd6bf6b6e64a9dded260b10ecad06d619fecef901688bbaf8cafce7d15ea14180b274411f5e3ed7a6605f7f00b624ad1b699c528cf6461210896cb52df085db0281aa42980340cf8c22457333a21e49d64da89adfa0980c13e9f94c737fe2131465ef636fcddf199cd1aff3035e88c6706d8adcbbb42fccfb526fedb03eab3db46e70d052a08a505449fc517228bcc3db216f110f0b8825b29a6f6c41ac92ffce49152e565d8446c772975a145bd2498970f721d6e60492d83ebed778eb3f02b163dbf9f350d3f1ed3fd0e935db4dfe3d72caa116f9cf0f8346cf97dd9fc527482fb5f23eb3547a7f7a52b20f0b570d37d9b76cf5587371782f4593216c350a356203b8c97cb904c274e08a33699d94e7cb3fad8589da9e578a68f4b3332760077d1324589781e784be25f4370e47f8be43b464e92ed4196bd3fc5b7eff6b1508d764ac314e17b00c398b2295615e5d5ee2969f3085f71f3ba31cc2b97965af52c529c6aa3b5f0c29bafc2d9ae38ff8d45ee852ed7c6410e03926ec028dab969c99dfb9791ff8437e497a55653904423088515b3a544f5b82024e72515339110e4a048afbdf90596fcaa66d448a5da0f72eb581140e4238df0050c88c81818c6fd6e1680ba00c5018be5164711ea78ce2c124bba77f04974f5c8b435f6ec9739ad2bcb3efb1a62bcb897199c79c8e3f7792d7be111c281844a57dc53bc8194062852ae52800005cb720fca065e5ccfba9010eed8e4dcfa309bf2aa1707400fd17b7b1a75dd429311066d463ee6248bc434d52d4e243e1bc0b5085142ec78066c1ef3dec58f6621bd3995727065aefaf1fabb8369a92bce163b8343e15d37953d17328dfb04e64a4c1689c7115f29ceb6ee90314a48b54a02ffc4cd34e8721f8336f6145d97637c0e3645b3a6c50ed4b7b4b4aca0a4bd3403cc524152d25d00ddbd6714a9aff94b63ee9b69c3e8fd37abbf274281cab1ab93c4fb17dad95556ef5b6f68bbc8c8d826381ea5a2df9f1f78fa04d3553ef1457c70f79defb3fada3b7c13ea907421693cc3f8fe09911c8615d7aeae47728fcbaa7a8d9836f391818303e7ff7a97916db648042dbc9dac11ce05c3fc247f44965180fe6b792a15718e09d9034107a7add9afd1e8644a8ff764c8744d2bb6434bc93cb1f83bf9d9542a7075f39e485f5d56d1ea2c2252927455d4474d7a68d3d895d66c127ba2e2a634ca246427f5f3b909fcb8b67ff20f44116397f0e63609e504da5e7a037b8f67e1636ee2577137ef7995fa3860145f29d8d648319ea3016492e11112cef1293ae26e8920f0af9e86a1a5da4281a969947b0ed6a40cf066ce6fe6ce032903dad23545bf16737e0c79adb8db0cd5aca2f63b88a8de2fc4d3f5aeb689797e2605c0d7dccdab5969733256e7e097e2f3804b9ba70a8294e416f4788b1738810541f911034fa86021ae0fdefbe96d4b379cbff63657620442380ef27b5d6a74814f847d115529009cb6cfb2b3f309fb483f8e1b39307797a9d921930fea758597c0be6f3ad289d510669446a80cf8180276974d84315e636e1870260577bed37a91d43c71791de83b0c09340619c47d138f91bde384e68a3a2de9def928fced83bd1fdce97054f8cccb4440e863de7ade27bb2da4221ef559ee4da1ff79fff12516fc6fd8e8771f36b6b9c49f2bd862acb9416c6f4873365234ad0a5f397aa2641f28e16c5d4c246667a760aa1cae9dcd5446635c7bfafeda6086034cc8d2c339726113971721f9039daad5158ae2c67ede5ee954378665e845eac401824c31b62af52e156913454188f51b5e56a2bfe64cfe7509bb8bb7ab7ce9f6701d2b70ab4a0a2631be73306b1f20dec7b41c35679e2f40e67a8e6b95d7ac0f656a1e3bd874770aa6a4321cfffd7b11d2d423659695e4ca40bbf8411892878f2f08b58a12e0c41d44a3829c2504dc00e52659a91e73c3b5c8d7643c246ba0f68b95e66aebc1eb7284436222cae0b383144c47995893196b18ba9dcb46d61631beaf659e39bec3ae876bca4f0dae4071338b17c06d9e47b773db0e5cf2c77432d88ce970d480331986d9520342766dd3b1f3ace0bddc5df21d9cb43a31616cc9ea738f79305e4e24ea14fc50177051fccc2de707eaa8844f60a9e730264fa2b715ee7714a4e0090d53bca75ebac2209396c9321a4688bf1ba5acfdfe3cdeab1836612862cbf5f6de03dab19d37d24dd267e65e50906656ba0d252e8512543128855d42534ecd54015ad489b008bdfb631fbe914f0a53142c3038c9d45e219a6559426a6c56339754c2e26fa2a97ec2eda14ca57dd0f83a4dcae4a8ea008baab115c733e872f7ae655df45af689de2283801cf5ea0a85636d77dbcc2e48003986b40b286b11fe8192d6a04512e069ba19c88c01d10b4cd9c52a422eda5a635d161523474c9222281fff46e8c5c9a4951e3997a7320f71b82dfa62b8517875e8ae7ae19ffe6eac16ae89f627a778c6125927a22c730fc5f51e0a9d45008dfd51dd420369e2bc30da15b86799fae290dc4eaaab318da702d6abd0f2d4b7a8f1316d748f8b191c28a5537c9fc5b684539d873af3c165e471eb71fb70197a5b95978fc1c1f24396c610526bf8e00fbf6173c0e3df12bc367a5d1b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h39af4e819a661a996089f6a3a2b20d09a912a99e991f9d9b79b6f1fb35ac59e19c97ea0927a48b3e528278af5153834c4b9ea3b8272a7e35bdab7800fce119ad7668ed7959665d0c9d3571f37fba38d39148b79c46e9e31c56341ca86cabfefc0b066706b42c43e9fb7cdfb7580f2fa2980dd60b08f15b5dd517321668ef6126c9a23af691c9d733152f2fa7de6d7dd9a7c51fec395ee6fb13a5f25c4379321eb4479064fafd4638f34597fafdafd9beb48253e4b131fddc85f1d99455e459fa262ddc809509764350786b96a8bd464f2209410412f9a430d05358169f1c12ff2493e24d7cf5b03c375fca2a98ec2753ef2cf3373a36f69261b44945709b614281e8e07a8ba3a12d3c1b166c59ec2d8f63a7dd7d8226d593208ded4e397aeeb5fdc19f169ab59598f1f2c3fec83b2f3e6860534c5ab9a64797a008a0bc5c60387d094ae2caaff4165d2ab5de36630c5428e643fe9367dcb0d9c85cb23098f67eb0b8c02b1f0537cb2a784a866624a84d20b08b561006e296140a28012b7c8b8c7e7dd1486e04e2e342c38230fe6387b1fd009605dd02b7e59da8bf4f7356a6a9de39bfe5ca1b2d66dbd0aab4265264d0469e6a17893839842b62bd4966bb3110134c65f7c96d72061724fef04790c3cabd40585c4e5111f9bbb1ca6726fb8c12c34d55e9cb7e4d0cfcbdb78ee2cec6e9494f8784180718f43567c6d12b7f0949df51bc09f2e753dc52be609475c05a80dee3ca40035afe8897555a6155bfb4a0bec8b2d6fa83dd75dd52c33d177108ffcd459caa1a4c3073e559af2538314ed1615145359b57115ff3785aca2a26da7450bd2cc494d3ee0bf958d4665ae6b923db72d12139cd8aa61ea5ceb1bf0417577ac571b10979457bbb309f8dbde3a4ad5191bc6b9b28e59469e357aa56c8e78c79b74d65a107964b7d38813bf70cfb42353190b7802eeb307d6b454db530fac531eda5e3df119bfc08e281b12265729452d7d109abdb40ccc016d5802c05ea461e4075a6c148d08e78433f7d8710da14714d8b49d55b225cadabd8bdcd4f108eb2a0b9242c59b39a172551e9ecc8adc1ff2ee76fe4773542195cc6e8d714faf90b5c6db328d0d133c19a14bd1949cb2853f8648aff2c23dce4edbfcbbf1f60f3caf337bc1dfc61c15c719db44f60a7dae4490b4bd1c1391b33ae47acd6af303b83ad9152c5eddbd58256a14db0c45809406b45ba1b0783a83e1c6b983de2869e6085b992c6be0974b744c31eca5f6775061eca70bb19001b074bf86d73b0abfae81ae9c21ead5dfe94dc3b3294158402e738cc9853e21a4b61d203962d199a8ded84f0f14752138c854d91fb3625fc4d71050905f46509cc5cf110e85361e3835276cb31e82854753941e2097d27982a67a515c1f52a62e3314fd65521356859ba6987dc6ac7614053fae52f42851cda261d6123d46a47cec32a5bc01818121dd3c0585846aad508dbf7a8d828825ebe1362cd8ec6d98f89dd0cac86a80cad87914a9fdf7941041bade630c6dc7a07ed7411f7fdf20e98e06451d296df19eb2c6a5978c4c62b6de8776a8c15c2e3a8c444503864e4aaf75018fdd91acaebac274fab6afa249f32cf0c84e37988a0f52b4ffdd4c2690318d403e9d89f764fc2327639b2a16a714b75b94f9e79154bb9ca8bba9b460b5e57cfaea62e47f05507c8fd67832cacbe6dd931235182ce24648ace3faa05a2d7205ca2ff251d4d9a03fe03f875b942fd3a64745a9017cefd9831c58532d2a6ab365aec4ba7ccf776d5bb6212570a0b193712d52ae8b0783f4284034ee54e7cfd8f251aa9ea3b45d841b04357bcb15380515fb1811899f68588edf6807f6f4c05d67fea840bedb114fbcea5a8bef54e085231d89d312e481118238f2283699b4c3ed9127a74c4a7c6a490a007b42fb6330fac75079f49e8a14a233f4e5deb3e337831c57807dff7f0192ae31ba6cc33f07a120beda4c461e479254ebd7891f6f7be093803090979ec1dd61be394d90b83da385c29b74903eb8c5c7b36daa8a1309740a606a61bae67ec7354f41893fa3c0b7af8020c9f531982943bd05b9d6727a5412242533a8723f30da50d938ec91e4ae419dabed73a0113f2c27b1ef8c05c04de042639b97cdb91700186585a19aae1e9a7073712cedbe56d3bde750c777a84dc9fa4954e335cbc5f4b283ab7eb0e948461eccc3b6e3dda3beadae129e48f769723927d83fb27cbbe2bddc8bfaf799ca50a231bd5cfb01adc36bc78c377f07bf50a9b5f4ddcaa878fae8dbfecfe64b3b6e725989338ab4546d6a909b35932a0e665c819079ba59629410c64911fe9e9a5701fee8a1871c4d869d722daa4a3ecc524ad04f2004d77fe368abf32d5be9b042e1597fd00670d73c88133fce6ac2b4c49f6449d83a65eef25922cf81596a1438d7cac812a5880c328c8c89f4de1b8a0d48b96e4231ee2ce33d708986c240f1315bc37db9ad869b5808b6dbc69396e86e8f58aaa43e5de91f653c0ea566373c75193312bdb10dd459d4b80e9598aac8ce586d57eb0212aba6d65ce89e2d5b3e39f491f358b0c25bf7c2d9123e80c5053447479f2631c7a9971e3846a40745d20490bc0d54cbd8933b133ad48cd6897fe251e27b3a2d7e3c3eedfbd4edb0b920882cafffd1474a6fdb2d4a60bb4a33c7a22773e4106f4d62de42f82ac667c4d54633ca3ed12be4776d88f36571197fe7d9baef5d961ec80a4051e3bc083a25526cd9e654ff09e57c43d3842aa256b0c3ac8065c90d1cc572cf491e56d5d25cb1add1b3c65cf175ba026d1e92da3ecc56684a6d3627bf8ed0e15231cfa8795eea483f548a88979bbb988847f3382a5fc6c981a1ed9ac3040f382e44ddf2b6799766b367fe9a77fb62001f2c7d8a1cec1bb8c8f9be8195d04f255020706186a4db707d01e2b8d74f4bdba9d701a59db7568fca9e5b28267b606c2e5eaba37fc736d3884cd70b77c31b36a8251eb43c0581f361b4a1f5c778b68d6857f039e55af7b5cc139e77eaa8b1500d6db1ca1ecdc0743f0c1de253842a332dd2adbab93525cbc7304b273cf672d8234d01a77d65ac629afc2b89d8af6aa39ba977b945df4061dca13ef5a5abfa39b43bb877291c6eff035c1b78d38fa48b5d78f63a334dfd59ded6047ce3d662278063a72d80feead70ed6a46b2b296ff6b3d6634499a6ad71197de3ed55bbbf077f36a15feb7a11cf00977acf97b13ced295e908a0ae37cfde5819dc965e0f5883ab18888ceae80ac1e55fa2c2ced5634a10792e9c7b63033166e2972eeea5854589f027f966b4be6f7405939f399aaa560ef53827b56ea8d5c6d6c8941dd07b1a08c8868204737d7e1e30bfe64922f5b8c09cec1cc916c65b3ffed596426889a956d28d0f367b9ff11405fb2d110a278798758491e87912ed3055fdeebf5c5d1e4f5806423cd405883068cddb474c6fb25c38716f9d352ae4c81c9e8dc0e61c9a87ea05355d0fe58be061a9d365b73e8ce1a621b0ec7a029e664f40c14727a9069d1e2f288ad0189ebcf0effd15406d9ca353ae38ae0e720ae4f4697a8ac46cdbd267fbe6a1559464ef8548fb4fc77708579ff19e62dbe6a267c88929bdde8d2c4e38f2fbca0e7020f7fef56506199abb143aca1083422b6bacb5ca56b04d0ad9787a84165c4ab6befbcf5e6a1072f0e1df796f3efb8422a91899e99ff01ff6b9cb78a005619745f81416591a8ba33699069f3443e60bed45ac817225d16e85d161b8cd82ce4160165ef6d1b67602f3d41bc946f793ece1ac58c78672f86efd0752b0f34688bc7625b2baa09a9b7f52c30dd9be489f2ed74ad83c9f2694124db2de7207d9755ff60a1693f67e653874ddf06bb9e47226640441ca93de6d4aca96f9f5f821a1f97dafae85c5dd43aedad8c97ec4265798fec3ea186202e70c4e631725d7a8e928d2133e7fba15b989d34afea3f867ed10aabccaa3a94a3ea07ee636c76a7731c6520beb52e18f9b2ef5d2bb191a4745a823d3771843480af9c481ed3ce1b35d6cdd6f26f934202ca5faa7de2562aa17c9b7238c11e6ac78e5ae62e0b0b4f8aa4847f991f745e6928837d6bcb86871771e793db5290d85a91db9bba9c595be27e76fb68553a9030b937e738b813461003fe41ec25678270673d905034aa611e32fcbd38bd53c615495da9fee565198b051531efbc8e42e266051df80cec0cec6673c85611300e3addafd3479ce9ba3cbe399812232f74c7b737f629ac13d928d1e6579c281848b99f94903c1ac148b6078bba221c6b059502948be4508e628667232238ecf9b8ef31a7c47d4dfe7a5b56488c864f7f708f1bdf53123d5c64fed7e86ed94b35c518046d34de90049e2d1fcc7ae2c4ccce95bb1b2067a3151aca46d1f51a299e27b9336d3bfd3ef5b77668ede56fc155bdf1805c8cda3462ea22bfea043d5459b5f498aaa12e9bd8304ffe3bd544f905efee70533b164cdbf8aeaf3f09b336be511f7ad2de84bd8ba1c414c919e3de9d1c10243f3da193bedb97d3418fe6b45b3fbb8165a9ab0bdb4d0355883d1b681b514ea908e6f9204d5929c97366ae1e899465d94956c8fb8e4db815cfb226277dfb3d8d877174133cffdb032c4ebe5bfe334ffa0b1568a98075204407871d6d2d3890d2f35a6c251a6aad4bd1926996272ae3487b50568b9ee29f75b8e4682fea995ffc55e478962fdc3cc574937424319e0361ceb065e1ce469ebe0dbb2b98ef057a6896a2bad0ad65d493040dfbc242fdf38912b2c1836d583482911caa85bc2adbb70e47ce20331f580b1b2d680385198253779b57e1fb621b35254ed8f40b334012b9155c719b276c6eb0f428fad08397e2547678f475b2f022b59b973a0bd90f3aa58a7fe06b48c6c1c34a4810a9ab87c9e06b90da6404e9801228d5f7ba8955849b42686a82fa9481d5ab0a6cbd7dbe69bd4f087a9b98d067dd367680dda770d0635637a5bf95704e849649e2e4183d186f058d025ab255e9d4f105198196556a7d54fa6ad05ea5427b9eaf9007149b75d3c62533f308763ef9c7f4241324a4ea900fd1876f7ea1e7080249438c978a1d8421a5e74f6c994a2f037a60c3dd1e9d9f66256253fa03e3b1bd247fae374f4d8715b44c55ab633cd3e61c16c72c50922f3aae7ba8fec0bd492e731c3304c34a993212b25f1fd8eca99f9f0f2fdd15cd939570af3e7042fece0ec682190dfdbeec4aeb009573ef5e76524d7d193075a7128033a4fd9795d5c4e54ebc136309937577e750ef85b901d1e6bd1243e6993b34ad277bc372c87a1edf9b0126ebe8e1782d43a1f9bd52549db19de15d4c33c8965e250a18a6f7b834cd94906f7778ec641ec3c014d61e0148e48c5124fe3ad467959ccb0223b82b1da6b210827799ecb91208f60313644f2cc60d2ba80a662eefd6106a022b8a937efd60fc26516f4a8ad9358c6c523b8081d27b05f275fa5232b518a33d0a9fbfa269ffbc954778856faaf095dc964132b0946c40f3e7e5a8b59d1e1fec5c017c53e5c144d51ba17ae29a8f8408583bed52684848fe239091e53fd4dd0af053ee8633fa494cef5f11e5958c990d031594e8342966be3978fd06d368a410a7908d0fea1216564311c507d011ffbb1085bf0f0f142bd49b0c790a980c1a97567536977a9c2fb8d6bca2ce11f0e067d970c2b62338d2e568055800de209c3cbf4796f4b33da652c4bc23ac14147d505f93561a9e6dc3e6e4285bbc35af6c97501257fe6b63edf418f71383d726b3efd8d762501122d886b12f533a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9fa95ca8bc5f89698dff6f7df5dbc16492f672c3c43688b0a6d2536889f954b9d7120826f348c803de65a10434cce9dbba7f48b2a15b551054aa2b04b1b6ae934d098e313e026152d034f16de4c0198921032e681c3eed352d6dd1e4ab89049f6978fdbde26075ec38f8b31bf2e9d533b587592fda4b3d0f745afccac8d9698ef0da0be42c2e0017d31a94b074ac8cdcd82cd7b01254b7e6d466f486cc42b1c9f576e679805d71e31187c9b14c7de1e8d5a924eb5b0b0c1a23576a961c1d11888cb84839bf28d8fd26df1cc1a45bb7d7f35e615f801ef7535b24eeab1342fc77f0678423ace1bdadb1d83d3484589eb65ed08c8b885a63d26bdec51eb63d020f3bec95d3e89d1673f7f0c59bed99e2122f25cc7313d20e5cc60638c890ccd4dcb0d3b924ed76edde2d8418107d8e3ed957da031ae4c54c3d5fe8fc3f4148456f77b24773cd1afd5a10d3b30c608c80221ffb2ad0bbefe607ab9eacec5d2cf71bba93455afe1886b9048172e85190cfd20ae55078cd698571bac2e0c28acb1993e6abc15e8c3aaa71f1262230c78c979514de842408b165d6dc8b4268ecfd20fb08762a65c64a84e40977f35d1ce65ed97f7da6e552ad270fc2513eb2f000908af46392062ac0bff4747d0188e90cea0e39e2fe05542cb757fee80fd3476aaa5845b471499902fe3d25bc5323ab02b66292af3ef93e49659a779a2cf115701aa0812caa7a343ed834dcb81614b3d69831b879ba5d815372d28f51e4de651e1a58bc04e830f9eda7993609707d511edddb4cd745b61c9e17736e92f94597b085b7fc172f0225d389af78c47dfb001b6cf14a3a7d899e8294bf7f6daa8248ba33b92cb84a47dc59e6e9766a7321aa509a6f5062f3d779c59e3c3915ce879b2d73d9344f5408866e8f2915541ac41cc6e73bb85f18a667c0642e04f95b8a96c7e7f5406758a25878bb6809dddedc8cd2ccfbbf58021c70b12d5f24e3fed552315c73da52936d03497c32e60c67b4b753eb6ad8859a779d44d3fb825dfbe45a66f1040966f7ae2e1a881a979c3343b18f67bf60fea6460992d4454655241e5ca66db6fd13f58528da16d6f2e849cb2dd92ecfe86c3aae69ca62e2e7eb599bded492e7aeaa429e4a5cec3ac4efa786b723ca41ba0a215c164a137d8c27f2b423dee4cbbd1d0913ad97f0e125167e5ebd86501d04edd91e68a3dadda2e905c4a81f5763b58f580963eca020c2b6621ea33b0122a90b0ab4671e415a1e58b4059a10d0adf0eb4572c74bb16ae06a9bd1d8523c9133a9b7f6e1f55bbbbdae0fe814ee3090766a89610e53d4980ff693e34e05723bdd7d763a634d00f9e2637e15ae9f6970f3d896c956aae2feffd44ac765e7c5267343dfa3381945b3faa79c4ba604d60a0193d76899f8d5a74814e67ecc9c786ae85c70599b323876077a9dfdf0ce623db47435305f9cd5b7ca4d20293b91ddedb1d61fd5f541cc213df82323c572ca781e81a69bfbdf6ebe83e981cb3e74333bc9a704deb4f61248ef13a2a836de51ab5d2e669dd527382ff91221a01ede88c7b33f90db7a96a9bf5b0633363d8eeebee92b9d0370f7608bc1de83de4d4f9ea2eeb3ddc498c2f02954dd834e83712a8804a5cc395ccb8f2e5ad22dfbdd98b7bf9df51629c54a13a4f68cc4ba24c8cfdc5596aea644b39d3ad3a4fc26da4faa7b13efd74b12929b1f99115538b0a8d34f7a1b6640af756fcdb9c9c6969e70c4eaa591768d87092a1f5688262b1cfa9370880f172f0985290f2c654ca9bd3c9318be766a2cf3a55ee56bdf4e01d33001cc005b27649443d2edd17b9422ce8eeca80fb24f062457d0d6d197ee08a2ca11f40b012bc4435f43712515f511d064d48288c2dcc6f7a20182c1bf07256c33e5c4d7d3f6e4bb50c9e3893f255238a50c98e53468aa8bc60975be80d0e65e7188c39c7738b817a0d94692da2e069add8dab28d049abc891af39259f59b5f5a56f210b1bb91482fc561742275c1033bda18d73b4554b25d326b1eb47b6210067a452bb32cd8979003d8f9457bbf0fb054654549f4b0422a7cbdc547ca5f1cf56a6cfdd84bfef748eba55cddddd2735fe5665807cb890150b17e0089b61ac279c98c744666f095fe96246726a64fb50afab82e26ff07db152b1d8912aa3fdb07448c4f0d73a04ac54c8aac5e88d09edc20511c4daa8e480787ebabc69bc39eae964695ac566e081cdd8a941ee8baf3167d2ac57d1745dcc310ac69650ca204b27731ed78c74b3ea323d35730e9f1f731dd002bb39bebb2c2020bfdb3c8054e0526246d896afdd1a4963954b2cd124b878716133a9c61bb13f170082a022cbba8a2de775cdb239595b0eb571c11f1a9744875edece39c5f8562fc8fbf0560f6073ea88db6b114c61447ec2e9ac3ee8d19d9a20db31aac3ff4b43942cd46a59c6619ffe8520bc514cb7e1282ac59963a2f5e2b76ab2743cec4400b70e8e5a396ff19c39c6f3071a950c68964db3d70323fdb9327f081de7038d6e4f1d4800d2ffb6a082ab53c142c8017cf14d440cd362ae76bb257dcee463cfa711641354111a94029b5202debd3699e4072cdcc9ea03d530bfc58bbc4f807a3e0217a54e3a7be1640291b26541f5249bfb1a741cc3c0bc574c72a58bca206a02447875f903cc475fe2adb127dc367688426fb2c7f3892aec412afcb25bf9bc8162b12423fadbea7106d55ab95bd340c295a96d5aa98f6eb71b806bd8f14736bf83adbc80a66500c5eb43c04e4774d095f6618fda7a49de8936df017afc7237f3341db57db819cbf8cd292087b9e066ecfec2313e8d9ee07cbb719c3d39d82979c05e2e350e8793144f6efe0a4e70040384c707612ef48f0add8d5b0a62cfb873ff2ddd3a6d50e764077abcbdff5f35e158129923a820c0a75f99a51ac84f966addc35a0a164699dfb645219c0d89ed4f053660cba40ec90cf6b99d49db4178f95dcf7ef0095dafed7e48b42743457b1119a98541bfd6fd3e9df9498eed6092486acc6aff696491bb4d7e93fce4d957742dc1b7d9ea6a56c3c3ff98ebe9ee67875ce36a4f531c967154985edea9e09eb7f78b8224a105effd5c60453fff8f8b2f70852addcbff3c8515d2b09270f67f3043ae1d984cdbcf244c48cb687551f82bca24e82f0466a962b15c164f67e70f3945b8b403dce24b4e36fa1d0d90105fd04e28b1b95996e37294ce22f03b829f734f0e253797130eb6c81159b27b8deebb2d839ea64b2261f1743a49d1e176bf571b9cf5438ffdef9a891f53e823bc46872c58266e520782b20114dd4d5b974ba4852d07e1afc5e9f80b096ac884ce5a6c651aa2d0efa3c1854bc3a1719477e9559203a6e6ee4456569e3aace3e7911d4281b39a808c4eb7de895c7d745813a87dfb8eb5c2cc9edd6383d0831e73a337e6d376726d79f40b5364aab30462f4d69c33b712b56a356bb268aca48103792a9e46119f5c6c6ff1b6675c8989f043d837ca901f7feec6fb7f9314bd54ddb462fee6896fce009f44875f0e0d38543e97f33e8bd8e9462c67fe21e79e21eab437a6ad23f79ccea166c8682b5fd13e55c73b1f6a48dc4be0fa8bca547821ff010fe8b76e5a5f9c55c0bfa93f77751edb9f7a4d50a6a80dbc8dbfe423db2389e1ef6ba4ff9eea79aa14bacabb8579076cdc249b990c6717054576c28989d6119bf0e9e4242a998fbc7dbd284f6bb930169347b9c934808b23622667acb6473c27c69b4edc2a985bfd7372d9f2b55238f3b49bb46562d5ef4d81f249acc394be28f316650880fbf6cb8c7a3ed81b60533118430cce2e14f46315b16f8f7139f59ea3fe000cc1fc3f43fa30e9341895fc33483a77a8a6201ac92a980e78abd70369aee481c554534a54685379d4736c0ffba59acb5331de05926d15a17927979f6946a8fc180735d39d24ccb995e49c1f3d67dc4cb7db29696aeea33b7ef6cea8ea9f348cecfb198c4f9e6aa7626029613301148b26d2b5b79363361891026cf3a18393aa0100cc939087a27359b765f01aff86245d2c2a59960eab01621e80a76bfc6260430a9cea74474a7d2f72f2e5caa9075f528c77959ec98699cadd36d9d9d0932d51422863b7f7dfbadbb742fe75e1ed2d569862f2cb2d2cbdde8d664a97b366cef02a1bb632801fed3a5fe4508767bf6deeb2ee3bc950ce100df8629f7f80e67db2037c6533cfa202bcf7fa789f8f78411c3fefefe15ab26291bb5d5beda1ec05d1d910af0f23fd7d993a6567765c7be80e0243e8ce505b05c6d672a1cda0d8f1b46e8f7d5967c9117031d20fda27c19d1df68799a6dfb785df8cbf441149ff6f5c00009776e97193d0e93700ee15d246d7c8d2890aeb5df4d603241fc57eb207084520ee21ac56792c47c3b15593408bc6cc17aa4d2f076738da19ddc399ec0f76cc4d621770b1a93bbb633dc62f617316f24aee24f9d8e9fa274d84a507079dd9b576dfd3fc3170b37e8d72673d320d742d85ee092603f2183f26dbac64f82328bd3fe8d945bf3ad655fd3ecadb3aa50789233ae4dbd53ea482a184a0ba4754a1b21209a841f700f6aa46706bfc2aa8eec0934f2e814959a20031d734743fcdc36eb231f627c406198dd2dd5914779c8048f086679f5ca5fb44825ce308c7a7c4f6400db8a953cc66a87e6f76a7b3deb23b40449bfbdd0fc960b4a7c95ccd27c4fb47f138eb8c86996f5c73362cad708d368c81ae2c74ca05173e624364fa0ebae7d72e2fd4c229e2a7b7d4743b9d235b794194b4834b93c6d2bfb118959ee12f57f3831365117a214d6646d425c7483b71726ec0fa0f694d113bb2943d954b63b4e793666c02ea4197663414e878ac77bca0bc746112b41d3c36c042716b63fcede4bb44d1d38c260b19ffadf3deb74f73c7ccbcca9321c1c43f7b5a0ae17975bba9554507c35cacd404ce4c42f7fcb87a5d63a46a80ffa7133f2b2556bf99f4c9fbd9d85a25dfaff70698cd24d933d57a045f40b026298335bd4111ab56d5b8e186d03c8001559928eda0a9a43f79adb337182a62f11aed3abdd41630959a16e55b9085cb46cbc4a932c852789e4325a2409140605b7583dc65b34bc17707cd3163280c9b11c98e4e0a97c2e16fc8546864df41180d7832442f827dbc36b70efa038bac8377cd86255172cfed27066b69f7e8acbd952606716dfa8ea28bf4cc52e0b082494a1d3963730c43949b7db428a97638971f7c9e4a40aa61dd26120e911153a5fc2e361124a504e4d9e2626277a484fe6544187fd9d7cc205e9a7409c5d37160d9ba43b728519a58e511d3df1419eb15f0a2fc09b58509a226df57e3d49f77db4e32eb3f8f3cc5f06cecd47a76d3087ddea004b7932b4857558b3698633a8310c52bd5157f548eaccb4c73c57afe075d4f7508f300fcd01f58a04ef6c32243b945f5393fcf87b308c1e4b85ceed721416456cfc82b51e53aa29e6642eee4ab7099ed7a2100de464bccb62cff55b7a641d19792ec19b6c93bf53ba3abcabd875dec0b3bc936b861bd50250f060871e3136850c66e139e44796945865ef3c864d896524d2c922b941a19962b839eccd110c17b81a4c1a422b7be3df049eb0e53fdd643ed935a8a235424f5b718bd984e25abeaae8cfbc2e780e80e0ca955684522b13f76a9f99db356e6e1d54c54a61fc25a9e048d466447474c6db1fd9c579a729beda08597c05c0ed9e3dade67f2df8dfe82ed9946b7ae0599f258d81165e28844266826cd73e34a46a8c521d9a4395d0e551ec853ccbc27e7e7b4cbfae62344ff116e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'ha3ec2ba239ba8cfa6923338f06172e22a9655142f9355a21d4d015084078026f886a429feb6fb3eeba06361f4b20851a50f6b32a63de82017687089b6f04c91048a960653fa941f4b9aec15a0a9a1ef2d8bc2896eb92242b36c087367744149046fef6c87d8c8c08149d5bb44f0ec7dc7046ec95ae263ff2f62b3a95fab0102020fed41dfd60e36140aa3b014db75237d0358d40edba4a13e06c22a4115e3f48be86070ed6201c3c68f99b723b9e51b38b52204ae0106c0eed3e82464a8fd8f4176f446425117616a210ba35b9dedde2985572ab8deb7a40beaf01b0092058f5fdf10ed29ee491e38fcf532cc6d6f5eb617729188c942c607669cd1d1b512812c5d22230aa62fa297440f5456ab9b4d5c4f66d602f30f4bc7d484d1d6edcbcaf8b1587bb191f75068ec818af3e392c1b86df7ba3f147cf13062bb8db344ad7ee392324ff4648efcca5448f5e1ba1484dced3470ae84f347b2f42319a1ba51276bb3a9e5220c57ab47921212b0bc33c39f6a94316ab23f3af0b37ca07bb09ee367c3104bb612b023d77c335bb99c886e818e69206350599837f3f996975662dacf1b058bea09aca1eda297edb3f3007a5b3b11605da99e04312e74a6b18ea4e078ebfdb48c2f24b0c2e1bb9780ca1b3796c01d110a1e0199284ffdc3d0a52f541afb2c9cd6839454585e6e5504deb8f36a35159d51354e472566270b9448a7eddf81976dd8efb651fa3e65ace6e2fe6900debb48ca01580b605786e31d00007608a486e4347abb30752b49f0d551e7510822530e659bdbde7ede1772ac5e373e88d1cbc96bc837591b230fa6d70a808afbc2145d052cd05d8ac85982c4298c068a15e0f7307e695d3925d9a7ef56e7776d78d4add4928d0be23a193d743edab4eb9c5189873a5b0e4e40b2746d677cd5aa354709d3b3b924c66fb4b0c66be888314852c0567a50cbc5591a93279a3de670da00a5b84b538345ef46f6f3f9de214869c13f34d168b568670f018ab0d42b1b17127677c4adcb78e7692489a76a4d394a3569cac7206806a14f02ec6d249cfb2657d073ac7aae495e01bfad94fee145894ee756287d00fd9fc81d63373d4e50daa82771f29e227a520a9bc64b7e54089872e5c1cda0a4a48df380104427adda7da6cc086c5e6a2521ca5507dd44f683e6544b3652bb39dbf850472786f6f21f088e440888db4983522db75c158ad3cf4dc978b2a4dfd4a9a900367f121628aa0a3853bb2ee53ef499f5ed2f21abbbb6147417e007354d06509b4ba88acbc1101f7b914bb777dc15da81fcb408593219bc62b4b84c68c3eb77793faa5f9ef6e93d7e7e0cbb56cf66fb37e5ba74191d8795c042571ea1330d5f3d96218c9c3c63cbe3ab79e7721daad4b81b0fb13f15ecf81000e0643af4697160e43ed410360b377ec4e3c9eda0726cfb41eecce98f1f888829793f31424e80e3b4c0749fdf577a761d5df8a12964059665ab1bcfb3411120577e1d1eb0b8168edc69d26b01ca25589a8c88c699a5214af80764ac803e437b8170218d435ac08b6d470b43422b7bd0c4909ffd4505273913d99216e27e6a2b14a5ca78d9305a6e7873961751ac76c5ce4eac11094f9276a976e78deec56d0e79714012d5669dcea45d0b509ac3051af16bc718afe0e7abd465b02a7aa4476fb4581cee6e33267f03579b11c33292761e6579375552daa70c99a8d85c1856ca4af8730db725a889b2d5388f9a7e51ff8ce1f5bb22d78194f695112f5862a0f073dc6900eceacf3df95169bf040d9279b0071e4bf7155885a19c7449b9f2675c85bba0e17fbc466eacc640ef335cf906de0ef0c703dcaf7b79859fe0f86353177dfd23a1bbabe6179a2d4d14eebffeb3f76f56b2ae23604326879bb336919a149e5a56afb0a0a3840ce3bde9c2b777abe10c9f17e2d00d30f34eba17f237ee4e5768f67cd1ff84c60abbfa95e68be67e2ffc5363114fad0d4522b6b5627f2dfee9adb6befe034e62ae95d435fca0fa5e038b67ff27de49081589963e4a67c99f88efbeaaa7e0448410cf9219564c7817f44a11467b6091a0839758cb7acb9cbcaa1bf8ad39568fea5bbf2d8ead04c03fac571a0ad61e2e5928501215375f39deee20ff855cbe1e1c63a42b48a864e303e4c0f44dc09c3b20bf3022d4270ce95dba06dfe9382104beba99cf2eb19c138b31cbfb1b9000ab19f0267a4d53d8a5feff2a5bfb3469510445910ef5350bf2a85e6c6b680782975b4bad68087beec5fe29bad3fbef0f8ef3f2bfc4c923fa46cb3a39e1bdf45cf821f9aeb5e700b021ea553aa0c7104f89ee601e8226100ae3f432d7fcf5afb2202ee13fb85cb1121c8167b9b387f395db72ad0bf835b7a7a35802f5fea50062b8793a82a62f0c2cbf6231e761fcb3c46c10922065727ccd3bed86c3527d3eba12cd2f5960b5a30517872861c52d66a7aee3c8bd22b9779b52bf40be85d55f24eea22b0354bf55df2354bd80bc6e886a51cec4b38ac50e66aa783f5b457b09a67e52271a2a04b815c3554bf25caab05f270e306fc0f581991a9e89a5feea94736c3965a35bc8666be83b59e4e89b76d89a5fc89236277754ebfee24c7663bf0c3ca0da85bc951160ebbe61d6edf462a68764ed45d4be39afe0bcfc5b3ddb5a4bafd9cea798314c74270911a7e5a04b185c82b8933a95af11721c94fafe7978de8409086418553a5a4cd3df81e3b36f0f4e8c0c5c1da2252e7a9355e3ed0090eb72604df9df7e352e26e3ff68e4fb22cdccc7f440ac76a4d421df5382b9b5f93d1aefc5655341fcd66f788b1f1e622148f7855b4688de51e8812611d4c2d725b45dee83e004556b8eb6aea80885e8777aa28303fc26536c63fa3bcfb93c326737be44285e20186e2db966f870bf1e4a1d5544cc425a1bee4c1da5909e1cb341824a4591d6a3c32ddc63589b4f930054c0fb882b5e645a4671aa5309b587dfe472978d7a9c6a3d2bfadd20de206058e597139b1fe12c795329c97f4e8462257364175723579e09b4c2a2b9d0dfb70f593e4e60748db49e49b71a5eb5976b1c16d1f9e975229b2a53b9644994db7e36ee24bb1d4d070653c0119eaec3eb15b20ec8573d1f3308ff6387f7bd60bd8f0941f614d920a09af231a2b9cbfdb7dc4376a90b982f666f504158b81c96295602c472eda93974f08fafd32ac2c5613ef0645023646a1cba6cf47c8143acc29e8ff468cd89e19c1ace8a39e531c57355b6e29f2697e989c2fa000dc3ff89cb6f5754b58b173f3807ee7de9b09c94c9a194f7e4672eead5227e6c4a8b057e494b237ed5790870c7b157cb986083a74ed1a20f1bc16712c0df2a624ef225644fcdf2bdf5dc95a07939412c62a05267e9aaa3a76394bb538fddc45605d367d7efddf58a2f32f98d695cf06209429f1baa901cc14c30d18ce9e3bbf68472f4e36ab66fe4922b23b1ee3c2f1b62810183d192b4d70be1eb45c4e2371b55c65f52e3a5fcc36b50993fb46c3b5cfa4154dbcb07eba244d917bd609b0b8b9e991570c1506abf739ef2164866f4aadab6348e6495cd8226c8e721df06403a1ff97e8b6e855d58d98c723fbb7b488d3d505b4c8157d222d4fe346f4b39c1b037cab09356366dba71f72bba3bb2a4c1e07c2fab2ea2222a9495614db07a97c64c6ba6e5e5422527dbfb04e8828e58d276c338011daa179b48e8a3f24aa8eeba9583fd784d9daf1c806ea7d96c564ff756a2eb096427b439f9d6caacf1a6b836ecbc049f1f37bf83491a13d4b29ab2f741f4bbd739f812506fada90b42a310afffdbb119531237ce66ad9a54c189b0d972f8f70d27e423440e01cf0b2e58b2728c7760504d3359928aeb38aac62f943518fbfbb23d86196ba94a80b50819d5ffe8e84f7c71c53cce85b041487fee835c740841271467000314c2614e009ededb89d899f2cefea2423133486200dd78318b07073700ab8ee702e1256e39da6399ede181ba923c9bc883a7afb0a04cb53cac57587635b475f03639fea0a71ff8f982d6a1f50c3e680bd46b440c9bf9d74030a8b71f3b8b61cdb2d1e9c05878fc3e195073db4b699b85ea294585acd27eac56a2a743b189ea491b2e4aaa6150ab258f593488d42fba5fee65cd616cd4ef60e9a2d7c5b9deaff6deb9fb40e267c66e9f6b894417898ab6b4e01bca3887c053bf4890a68cfd7b7ef8e36fb44b0124b515061994209b5fa8db6ab096c56fbd55513cf88f4cc1eb3a309f15a310ad3a0a48e2e7af9ae2042b0d9b85fa0b39fad6578821b16c82ccdce1119fba9e57b8fa4eeed2aa8a6977203bad3b1f79223f1c809c12454d79097bd495ff87fd41a95e9f9c64b8ac5ff75bc97840280ee474a4849affeb76134892e233dbec4b22fdd95e083a1f45935063c709accc39f137e5d2eda2fd5484b9404b8a1ef27b1a472e287c0a4cf7169a58b77643e0bdba987d25ffdb422af47a1e7b30a1e32f7d969facaf7b5ce84c83934fbd42b25c8fdede45915866f28d85aff03a4d9bd435e3534797a3008f6d3cf29e606b9109a7ba5433aab50da47d79751fb2b8188367ee4e72290b85985515d9395f9f02f30fb2e632d84444bdf1408ae626c4afd0475d2082b8bcde9527a462795e8d79a92d572283d85edfc7af479a24957a0ab11c030b89b80fd8c21c57159a7e8bb0f3c82faa901226bcd98c7ad70d6c878e8f231b43e5995005a24a6f3c5c2bde35d689dd0ee94a86fe5ccf20129d96d8705e2a2425927d7b66d46044a8b0a45e19728bacfc8299091a8109d1b221516970b6474d47737e90503e8ce5c3a192dbe79f1415b83081cd1508ace73fd46044a41ac1d3fbbe5057bdb5a09749ed0aeeb2dbea957c95871c94c99411f179d8bbf6120b20c4bc28c242b38e42d2278dcd0f4f880fb5e979b6be535d32ffe9e234ccbfab484c64ac3648081b5fd08780199cd0477d4b3b09ea7e2f82f74ad4a2374605ee63809fcdc2fef81285e2115ec7d0a8bb4a2599764f86ab92cf1bee61e4c4d9fb3dc61391bc0d5c08c0be207efb4b963d8159f5380d399ef6a7a98d18b0894ccd26c7ae5b8dfa890da3c29d960b5c7b41a489982aedd4191fa247d1cab1b0c4807367bec4322d0c1c4723921871f0e95075afbd47bf200d8a8333fcfaf292dee8ff8eee86a11c9a1e0eb5aed61b221b5cb6b53c54251e6267ab9bc5133a63d96ab0364eca578ec8c30fae47c8b08723755a4a53e44205e234278b4b4998110d5378d31f74bff27df951006ec94ef6c3c36bf77ca2b6d61bb833a21f8d8d1c279acb1964482b806b2b814ff56bc0c88e7742760b114c36c29b5903d198cac06edb84140d1d5aa8cb4e16867737630efb0329ca0ee61944f08784e932080ec73826e755f41512c44defe6afd7de04565a2783257c808936519ae9906b65206cb4565eebcb9c6813857a06e95a93210bf61acc4abee822a116dfcb495bb745c873d32c8c35ced3c31802f7b17cbb0d56daa1c57dcd4fe03b80d2b77eb58864665964ae64a7257a26f56b6a1fda42e0ecf49efca5011560993ee5e34fe8da49145411dcbeff634327aec78a54cd7cb5ef8f32c7020d335e8a1fbeb7346bcb15a58a1481ea1fc431681e095261490a995a0b75abbe0626394ec98edd4e970deb16475d7ad58b6844ab8a42568b71ba6233798616ed55bb0d4b5d203e01f16822eb336fbefaa7bcdeb7b10c22f2192c271cddc2e7d477a52aca312a15224daa63b731ae1ad9f57d61bc6fffbf3338af3679c5fa84f99cf97b39f8b66d37b0d4bb8d127f8b518;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h5fde5ec29b0b1a5cc85e9da22874174ac8a16ee46561c77d3abcaa10bf1890d5dcb2a85ea458dbda550823bd692ec60cf2c3ab2697d66c0d73320aa349b85d3d608d93db6c249e5417643f7f47cae670c8fd8a3191bd9586fc93c9b2d9b14d635c0e7777c806faae72f0a01af8bb4733bac7600dade051360fabf439e11f4564848a6cfe1319c512a7d8a3df6c05b5e290f386cc0eb5f0327750cf5aca164118b183399e432ac32664e922776257db3aab092ac3818292b301ff8f60eb0af5972f9099febee34035ef6c520c773e15a778efeb9071fd3b438a28531420b349e5940e153dc7c2d69b16c45c5108aa21e630a17352e18ae993ebf14face32f7f2fd9a2a049a760cd075c60ec7e537a11ec18c6309deaee3532ec3538a3944e83f5e468b82ffd4d412a29bfb80baa69eef22b9330536d32d46f73bcd96c3b0f7ca36467232ea920595031425cdfcab73d5a22c6ab5d45bb24712f34a5c70d7c989061efc29f086f441c45b14528349a80d17fe60ddf1c37d31673a179273f32171bd33d118bb367242db87d632b09439dd338036d61232349e8fd5abe727accbf3c3bd4a68584012118a2050e176892a907490971e38eeb5a6ae857fa5e59f9cbed04fd7736af0433472f71524a07982e88233b8a314a9fe292333abaa55512c74dcf00e3615d6f5fc35606ae49c1431407f539ddd66755be8ff292967683dc7c7d4234b2f777d895c49f7dc89f8568a1b6f267a2585d0e94aecfcfa93ea3b05f34372a7735530e60e67d1e3ccd47ae371e83f1ba79d40cb191704bb33c82f3047775a99b678989fd970b20bd23d92a3f1ae0b667aee06da94a10177d42d31f8320edd3a4a3f8f2eedb78dacf1d631e7c6b54c40ce68eb868dafb2b9a26d189c70f33f7c1847e94cce2811a69779818c5d43270e1acb7fc37c59396aa15e0d97f3f3248bf8c30bb59085f3978203e8978fe3518c20b72fb2d8d94e8df38c3e707a1e4e6120227402e54d30e5bb63d26f1f04409d009fcce28dc2af2ebc1acc99108f3bf7d117e2864f9d6f98041aa88ba1506027160fb0fe996918851e3b31ebe6239ba404b3e11e8fd724d56a23e6e2535eeaa151c5495791887922c01f72d5cbf14f9b846c3051b38292bab1dc5bc17c7d4651149d6fe5cd534ea7efa21784548f6a1cc009d410446312567fb3e6d9b71d0572934f06089eedf9d8631bc0b53c4063fe252bc6991d003433b61e6df227446ef95c42ccfbcf79742c115583c0d871899a70229f9cea2c94fa798776293a6b5eb50ad404f8f2b2529234a8e4f3e4e07bc9b1b3567c73d321fd24724ca4deae15359cc501cdc03a5ec82d7be4b7487000354aa2e0facf94956c0ae92ce5bcfc05d99f89249b26e80eaadd353cb47c4447daf813755de45980d45697c30a3eb335014424d34233282f007cb683cc3d5ab0ec8973da7f430486ee3df592aa7f7939e5b13c53ca26cccbdfbc75bf252108c1d24ea5550028eb7bcb2df6e9d02e8c93a5a44a397b4cf15ff80f9400448e2ce1703fe3ca9e8ee36ba5ff9972275c95256660eb49f45fdc19cf7d50dc78e3dda72d39d5ead18e8b220cdd6f3ded0a43e2452c085cd6628b046b345d0bd3f48822f189966da979fdb4abfe0d5bb513b29ecf8b5c1d0c0ef13bdf0910a0abc1432b2bab2914bbb48cf1fbf9a4a729a76179fa07b0b81fe9c5d217f10e94b4c60ce8c8a49d2589c89a18be16110bd49caaf87e4ba28dc8032890f24941d785ee69f33ff400beaf92f475b071991418b71a750fc9f18ca405a7da1220a467926abdb9ac8ffaa9228823881de720501f5d4d143950dd81e9ae99ed2804345d805ae4e517e3e720a8a5d32e8c4e98d200dc40086c0cbbeaa42267aa63ea1ea83a75320514c6395d8c3d3759cf0fa0831f42f745bb1a5ee00052baf13b4743d6a2211659c0587d3fd7e03c918761043df2f6058b3845a675a8e2afb45381ecc2565778d9d79410a7a38279b280eef9a938a38bb41a0f4ab5c46756120d69c3d029fbfae429c706355060e27b2760370c698efd9a7164dcf74763e3e948d226303def830b347ea80193b390d0b04cee7260b51319768ea6a21e2f763376057b3066293c65a0a4ba5ab9d587ca6629c1f5c4d788abc88f6a4e9ddbb4eae9ef86dcb95d52293477e061a4da30bfbfd8e5ef98e5f5cc06c607dbe82df73c32167378e24d8436516abf969b13dd7894e9567609c7d74b27bee0673577e2bc40598f3d41e023760d5e9b0ddb01f94a6d6f2463330a8be1222ba3a87104038b8845d4a5a5ee4b93d7c1ee12306066f276fbb2ca587f9951f6501939f2522b7587abb32b6d5da41d638991e889764bd683a7940ecb637f325eea55a9ba225d601c074bdde51df17ba9bbb8943cade8d98be8832049273b5124a46f586fb26d77c54892bd2aed7f3cbb85e7bf3d1cc5637caa71b0b029e7ec82917f5fb3f0d8685421b3e57baf19db61725f13f5f0a2b3548a5985867c8a98612abf40cd9df3036a3594ba01e4b66dfb7bd6763f4c8552f892694cc497d727d085df94a815464df989e692578772c01c9f737d14865349d909115bbb335c269bf06badd317332968bbd1455ba7cb1253a76f5572ed1cab955bf21c1b4c5b08d932cf64f00251f574dc258dc88275c8197cdac094d5562f0b7298b63ab36316e9cf9f88851afeb2cce4708532faec3ee3cbb02652e9bef87860c9610552bfdd484aaff572a1679c9e6e62e3ae411f2048b115e97ceaf87f64c3bff6bc29baf0cdc8083bed59999daad9c18309397205f0a015490ce03d225163e45c1c92098e2c17f68527e2eab71a2a5880de36f2cfa9a008df4c8531de810944d1d0447a4cd938e7c7e991278d85aa30e7c4a11506adec187c6754caa72f0480d9770cbe3318605cef336d35b7d4a774be0afbd2d3d5991acc252aa7d4e3b0e84e35f1053e4c2f3a92aebc177f920fa48e41a12fb9e21d944b22cd2d02928500e63bd3dc54b78cb6c37a8426afbfa852fd83cc283e358afaa9cc62de643f29aea0e773bcfb36697e47186d8fa9245b33fd0932500f1a3a59d167f94ed0dfd5bd41187f1a9f0e82ef7201a24cc95300e87a179e28bff111106862e5322817c7bd70740348a20d48c041f78a40774ed1b722de8b31380a7281193e46e11de21b64933e7f63ab3133008250bf052ef3115dfd2fb4c0d8584df925c969732c6e23eea159a203e5c9e4baa75d16707bc1a9e371ac69e1aec386820b346a1473e100283a89cb36e1ea2989ed99d2ccbc65c106ed8b3d9b415d65acde913748d7b48d1514d5c4a588ec72cf943735c839ca24dec0b38dc0efb538b87f8a505d915c9e19936eb3c15b50e258f6cd4b9873e6cfa6c47c55b21ef53ae0d5abebfae5b0928c98e16379d99a415e9e12d2a24fb216f49a32b002cba970e82efff1bf2ef6788c47490b0c906f107e6af14ff0ee6f59b69d8c4d6a82070a7134f8869aa9ba689eca14c95a1d99a0237bd283296b6e8ec16542391951c6ed5a96921d2e40c84ade1bb48dec2898b13394c8864b4ecbd1c05ff1c2bb9f03bc7bbd3a88320d9ef72b4c7b7379d0b2c74cf3ca3f65132e40f1de36ef134c4e6d420d66913711960839c51c9e5e416d4ebb2ea643771f8cdb4d15cfde3aac65051d5e616d8686baf5cb716021ab464643e8d02b0d5dc254dc7c7b5282f3a7b525ff4d60521088a45b5179cb24d9e90ded244b2a8975d0a840bb64f666369f4ec2349acdc37879804352cef3bec78d0d07751029ef68e771b99984c5a3669cb514df66ab601a8f80c18fdf2adb29ac31b4b12f2a0878d85714fb1797d8460af4eee3a9808d08b06a0e2be805e9a4fe9a33ce71c5526b03a00b1a9e4dd0369dca75535bc63953e04c60a24d723c0831b40e8284ee0e998fb2bdaf31d17ebc165e6124e3497bdc2e55858ab64b2d359d4b2e78317006fccfba679b2821185dfb98ce96ad4463329975bb7e74d9d7bba5085a15466e526374b17d2f70ff4dbcb235c50014d6f180397704eb76f97ee8728774fbb69eb1b8aa7b2a372ce0c8144f56b6f2aa9131eb0422cf8680eccf0bd8efc77a5cd1e967883768b094694ba6dea0b8d31f7e3dbf340d214f82390ac4a7529c01dc3c33ec6e45ba514d72fe0e9fc80064bbd0607a92991f67960922373a39442d169de74e9dfcd489b7ea9a0720020cec0dc58de3a60d3a807b8ed3163e99a838aa88aee0cb5a26053bf88b113741a708851c7d0e4889dd33e274a673a978c2d5ac46f0f6731d9305f7d4a9de4c610338cdb6576d9030ca45f8bf48be29c959dba51d7b65c52929a10fb7c9561a4770f09461df828142310bd573e652d43d6c9ab1a223ff371fa78f8f08f5e9f550b3bd0abb66d549fbd58cd1b6d27901c875b7538e64efa8bdc8b8404103185bc81d36f7ad04e2223758364271a9e5c6a678a738b6f5ef9da3c8a3baa581df1c5d82b8c5f3a9d539d369e6e1419e207a2b27e6c10fd508e45a997af64a4e77ddaf00220327b24545636815b6ff5a8e3bc091243751d3a25d5dde51b2fb616a79eee8d1db75598dafb630ae83c19b3e2ac9d4b57107fd8535cfa4918417fc3667b8126aacb6557e2d5dc0131e6b6c419238a195ffe553a2fb60b4b29d4c7e06ee4f9ce1ec9ba00c6ca444e11fdf799aaaa50356b079321796461b3a3313324dd734ca8ab5cb8d469a5a44832f19db73c00ddee4e87a5875db1a323d23df3898cdb2f369747720bbdd23649db83ff58c989a8ede57518653104011998f1d66980479a2de911454c2dbc47c189f317bd4946e24e0bf3af4c3e2be45c061310c902e3105bbb32cf56424e34007899d2c4beb92859365b55c6f5c0457824dc219be3639aa0bb7c5a56697ff81b2be81e04ed54867715f96802de668e4d00181e678483f657eb8c40acc7b64abac72e73934aa9b246c04db06b4d770b2047142ca1e0a43ba42cd5403bae4a10c00697caf26561002dd756f4111bd11d323ed152ec72e2a799c7d1c4eafb0f3a89b656a4a41189001a915ab895b3628870f6f4257948b37339e768bc0067abd11a2ef27c41c14c40097c0fbd28f8aaca7df3983a76a7fbb80251bd6a5b776f8ed651811d7ce84ba193e38dc631430d8024716c3323d8f6b7fdc65c933e87874a896735ee49966ba0109d0cbf1957076bd64016d1fb04a9e019062c48270b7d8382ba5146fa465d959263601115fe0fe0c1e7f39f71ce05728d0904be5895f7a440d8012d5fc2fae509003c6e27ae92dfd3dfc84e89ce89c47fa35c9253e7f1a390f6f957183393b687656f82af0af22af5725e6d4f2c7298e7c78e070d8c83f7dfd077153218605b0bda39a705ae106882e322d37673aa86dd32cf9f5311a7cafd3f20b4edf4a682335a39948a442e307ce88e73aa83dc0c967aa0d5f20bd6cffc3d4b27d69cbbc4853b5d86a45bfe32e5e8a783a3461387c435b3da34ca17fadb43ebeb349874bcd11649b405ae57d4e070764871878b84ae397d102145276c32c3c8b7e5855b77ac1f4e63747764f82a4750f4b418142a3f87f744a944170e7fae3696f8ddafadd4f4d0494d26e78192df7a6a22d67d8562f8b135f05698c37d2ff65c645a5498d29aba3c5bf3756e160f3035dea29087a70a7cb4d01187588ef308c8329da1b4b882e795cd4aea4a81279e451ad518ab93eca9bfe3003fff9a08b2dadfe4104f291d42af191d5f5dfe6a91d12944c6f896b1223b9d03fc713700ce433e358a4782808e48e1fb79d9ed08b0313d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h758d8dbe6eeffad4b66ba297cefd33521ecb980b29a9d79b2b7b954443910af1133273d7d7144831296872953a21650bafba85fae461a8c2180af525a61c6a1abb0ebe0368e5194194500ca526a6e8fae77f8e971f7c4f6b0f85cdb6d70710980236c00360feb0c645e3628c748aaba13c515b2c68fde5596d805e9ccb15b20f0e7f4caf8022beb13f81c52aea95dc2b8a7be9b0c6743c59535d0ddcf9f270cdf29184b8e0bb495b850e6a3b463b6df9966243ce2ef25133260f382d0b23d702f025489d27577bd7f5b9bd5fad0acd740d1df0d9a4db0ab4ab4711d370933693f40485b76eb283d33d39b04ddf749038b242eacbdd2522f856e81f943e0aab0f046ab42d668580610f8fa36906ba3a4606303b46e401228d4b601667d214ae5296c0c3f4b87494bfd15d2a744547ebec41a905fc94f1b30d8b4ef0257b6c43ebd6a6f71b322cdc5756587aaba8540db3cc60759ff3c06e039987c9884b1dc5bb0f4e4a458e1e1375cf730972ea6ff0e2bdd20986ccfee743323f7375a0b18fda0cab279904fd1802ed4e11a801658596d51edde3ae4133b9c4ea00f94cb60e9bdacb58ca2b78b6f21ed7586dd861b33c203ba774c07ee1ea8a646117173271294955028b42fef6d6e2e4a3db03fe78e20085850787a059efcfadf88beab969ac6b6a7a7b1cc73a034d5b070eb2263322fc802f5052ada1d2ade392b55816597d1e648c488ce199650f41146c9efb377711f887bf8fd8e22007e45ed78597f8a1b0765f9c8f5f3b8fd8df07a1fc91147ee1401369932e14357c6175f72197c3159455099f7760e762347965a7b4a3506b6e1a8e31bb056ed07078464743636022102dba681e9478fe9d3c2c5d65404d0b0d70ddc53f82ba46f8c34d8550b36a239d3451ccabb106900c1a9c8b4bffad2c5138ab3e48a25efe77bdce55a40b65db22e00b57fdc9f1538fd03cc3b66af641336f9f2c95033555d2c69e641e47e0391d552afcacbb085463dbaf7074e850619ebd96e1c78ef7a6e837adf5c3bfec721850aadc450db7cc7f55c7cfcaac9602907882ef09a0f28593ecf1d9a5650464814eb1a165dbd576abe09a8cf63bf0c35bbbb84d4e1623317c58eebeef92736fa96fcdd349aef90cfce7c179eaa63b97334d65a1745161d6ce9a57460eccb79cda77c3c2dcb2b80db41fe290bf3015a9a1d034dffcc199461fe202239a8de056d64e4a3055d68ff4d0e739e12f6a9414cc8f06cc2ccc700b0f83d92e78f184b092cad7744fcffd4e8c0191f7f80816f384f2c17537c8f84a967f191afc1dc210cd638907be0de23da1d7b13442f434898f4319db30fb502e9b262c6fdc0d5f1ebaa1b28097969779bd36e5152b3bb7cbdfcad2fb67160479cc66259f8f718c67662faa4730fbfba2aeca3de41e3b978b2049045c612de60de01ae1a527457f117ce8caafaf8ff5c92a0892d434c05a90947281f3d2309bbee0aaaf235d55aa7b3795a8b4ca97d830d2dfe136396679794a528cdb0ddf8c6dbe404223e36abd94bd9da7f95d403d1d6c2c0d198c81d5af86a664d91655eaeb87a9c5d8fed7e0fb71a4ea38daa566e1a5cedc5e61dccde0fe25536b91b090d61942e3aef6993b9affe123766d88691a7ea693e982747084d9aabc1a7aa6da9ade6c0081e54998aa57e820e18b4f6a438f8b0664da4b8629b5ed91e4a01e27c0ca1fcd8eb9c0c8117cc43e259c9d0cb34d7884ade0ed57ffed4fdad3a792ed75c2accef20ec7886057e6fbe8dbe4dc848f5a83407aab5f81cd83b2c33f49997d54d10d4e87ae5e522fe3612653ad24a4a15725b01fc1bdb4f533905888d5aa0f12e01656bf655ee9c970b9c4279a9289ef4b328cc4648f99cd6ac83363395c8ecd8a2214bf45ad8d58aa5ab9b3f010a1ab48005258fdee10c2b9c0a3430d8e25c1bdd91c3ef1a0045b8a8f00c08e32f868e6275821366659ff76b1fd87962d8a230ae80b9b31b9c2a4c063dc61e03556e96fa70bfaea935c793c1b950cf30c8cc286baaf8c258467be17c5790dd3a1a86e5b90e56b94ba2c6f8e4fbeb89c9987bf3bb87671069fdb3adda6d153ca52f5a76f6c1be92b9a07fd17004662e8a930176ca275d9c4878f4d0738f55a18cdc5bbe187063ec909529ef6e0de691bcf2e73f4c11d4da659df88b7f5cea3392d5f372dd2fe1b7edc8ed2a73e6bfd74be19d7644215d5d707e481ac43b7d08097b5ad9b10779cb0161343525c8fa5f16dc36c1bb65b738eb31817bffbada09f18fad77c714f5ae3e7bde87ef84548e3a8cd4b1d37f73c0742835b95745c50efcb94197b2a1618cd56627ed04323e2fa6363e16d1bc4bd34a2efb9fc4cef072e15410393160360f12a8153e26c24b83c69a18ee6de1097f0338cfad1e637ea9c2fe6f7b3fda6b3f1874799a3ffa880d4151c0b1196eba9bfe457d76720582ac1671b0a0a7a53bb0cfda6c2fd4c860ee45cd2647b6b2248eef5154ec9bf95d92d4c5de3e6f0f94a9d1def5f5195056135724fdc8d500c1db572267b8472d8a8a8ce5d20e10f6c26c2bf147c4c5565b5aaa0a7781d9d399f6b694298337d04ef803a8e408f0349783dfdb5cc62253a4054adf1239d12ea1f255dfb07aeac8c4b415fcd19f509f5043a426916387d1144ad99113c9f67a50230e86a0704baea385caa686aade1e98fbf235aa35755af11a10d36ee10d6b956087fff74c19e64b8b332cffc40cfcb71563ef37880b7d1cf545d064f8ab7558d80fbf7cfd1b2346a36197f54d7a1f8463f5adfa14b50a9f9b2c54029a11fff6c22d8c5c9b79232037a2362f49c492e6870db26627961927841c184c7bdd6261421eece4d2298d71e74d54b7b46cc12479cbc09e9ee7549972b5f4120447ddfd9440a4ce2303799fcad60cabc12c948666a8905e66c37b5fa40d20b8892188385e82d2d595d3be2614161b64f4c0380f113b2ec2b04f1bdd01e2c4490f1d8e6390a65dc66c6162621e06992408e164cc226aba5de1c65b9118459df692eb72c5126a63f071d3a7f48dd88541cfdc3efad5cdb58e49b95ebda0e6bdabeaa84e4c531933deccf51edfd584cda6b3f285e170203197ac2673609476c1f7f5a21c5ad7e2db95dab6d0a803c72f9af3377798f1351dbeac558ff9c634dfcde8d97ca7b67a961590a46f490361238230f63b7d392efaa7c044088380bf9968481f621d3a983382c6d22704889b4179e27aa91e5d5902cd32a5f687cb14550fdd8221c84da90f01005c42322e3c62263f055f9dfa31bdb34ab4d132d6ee866d09b25d922053a58042b410c3527ec105b123a1edc7d86c2d56b3162ffb36ee6b13c021da05145b12994dbff8282deaf55cc3ad9fba26e49b6e51ac0c9c621134d9d909fedb6e53eaacf08166584882c46d2a3f3ca9a67739c391f6ce8355d9beea1ccc4ae556eb220d07694285eee557d6ddf9c9e0e4e1d058a4480c1bba44904b6407e7d79b6395b56f41f6dae3e46127292c0d4631aaeed4f046d1b1a5dff4dd3d8e3a4160069d75fdf883da6c217016f1891aa7c3eedd97591024e8817edecc1ed935bdbe9921d06b8a9609bb0b4932b4e98ba5f9bb14067fbf378e6d47d7699c63377e0867c9940eb8fccf8aa0c557d5bcbc1cac8b35cc419cfaf30184a3299e2b83a9e27b7e8860b54bb0ab4978678a6ff9fc31212a8f8f6f705a85fe971cc447f89f8c35dbd90b2e097ce5602098bd0530a1e269c09454374142fc31aa97cac34d4ba2a726cf4fd42b1c70caf663772104f29f4d2e5e63c6bed045dbd8be14c78fc729218cfce650a41924ee058302b200b56cb70f47306b78cfe048c763e3ab46d9a6933119604626c830561db155bceefd713229de90d0d57f284634797087c8b58c084e886146191bb9d0db57c7d952f92cd8b08100f2fb0375c5a4438f7b24dcdb7b4105bb877f855ccee782a1c4aa97bf5a93308828da4bf82cb72d4f01ebcc4fcf7f1cc8ed4f47dca5d1a544d624e4a9938dce46ef9ac4c703157592337fa18e6ced045ff9ad778e5ce497bb6550cc0c08583d6bdbb63b54eaaad8d6f44fa37b362d8894f5d7ef3922c191ab1216f36f8eb4ef97df4614c6d12a9681aba0dc023a53f23495a915d8b61cbecfb6575a21e0f12c356668aef4d1a7a9b026417c3dd36b1ec20b10c23793ff1a2f6bfed58075d2eb6a074a6a08ac88de56693f22a68c0d01f731720caf966f2356a510100eeae2e28d59fa8e76be6a9a79f18bd45620fd103326e316fbc5d2d32f6da7858775d18c40141f3f88e3266033dd81ff09044ba998795dae8cad93bceae1d9f14afa62c27223ce2cdf85de115d523814040f4163107cae4423b731e006376f5c8c4c812dc42cf56ff7eb15d3bd477fd020e4d529525f2195f3b8e2abc98f7ecfdca5ebd2e63d0f8e0c34ae865f15a0f63f35012b5c0e16657641e267501ac3703073b57148bc8695c5a128cd1fd8e2c1947873868cbc672ceabb8456674430dbd824a593f52ffd8c8f30bba5990eb2dc0da2132dc17daf06127c639c5f6a8d7f84c7292da5d5f4ff65b45b736ad505dbd765e2cfd6705bada6124e6dd36ef739b925d63e67d2d78227d413f5d915f543c138f1bca0678de35403ab968d6bc72157d2af3add49e765bc565f68eec2817681c8b34f8087cbe0d994739217c70a5e46fe89524f7cb52ccff13b16f45b26a9f66ccb7d5dbd2122ca45c9dd4a7d367b326fda06255982b52f55e6a343f7f3734352e7d4a37ed196899f399168ea182d041fe2d91ad7c34f2484426d2132070058febabb7125d0a3784f4de97d90f238534751e2513ca73164f189243c06f8e52784f0a5ee5b73ed697c83ab4cad9b1912d3fc7c123101e6038f11c082100cd3d0dc76252cc98d7529903ceced8b010688ee49faa72dbc9aa9ea863558920f80d60f6f0f481e530e8cb1c3147ff1b71ef280eada9f86b7650d7123d009b7a33155abd8694161bf74fa9f23ddf7143d7b48c3262267d7b90a44cf7a6ea5a786f2e7eec1fabba058f0727aa3a25fbe3fd6ec4528fd8f5620e7d9780129a571232008efe8303bf606563b379053debd8d6d969e69a7e767b7a2e227a75dabf52469716c998f3e8d7f957702bbc7c3fb07e5bb75373a98ba58cedb626ef7c432c16673c8535ba14f2850378f6ab6ecfb7c09765489f49cdf0e5f814976bdea88ea5126e23db44802a63945254386f8ffffcccd92f58c9f7abba66426a5caf6610c4a1f54d3ade2ccac4c21c96c0259540ce4e954f117512083b89fe91794ef97e89360e6f3e25cbcbf2173e20941ae0ff0aee9d069a6f6668ebb35d0df238f7f613895ce2fc6615bd91810322520a3d19224c16551a800334f9b3265134261607aa4f9993f1e79f01b18e2a374b4b763401de81c9ba89ff56ed7bfdc6878d629908b9f5918722b66aaf8489d65cd4e97e309a22bc963673a4ac1204b56a7c06f799638e1b965b3e55d89691254ec4bc77e6f4ae65de2c6f03499016d8728738a1517bb0de2493c30f3c2d9bd86aa3f28282374e83db5151a267015f6782cac7de31f89a3fb6d1807f7cb553df9cd5e208db6b4408564d50dbfaa3acf051f5f40ad174c5dc5730cf3ac2c20cc5e482865d457bb2c260689645f134b18518f44877285316d7bc22094c058035b00716eade4833a7b61c2d61b8c6baeaf9f2c569678a631f4028390bde1b5db1cbd5ad7a435d5e380d2ac505ac43361d1c25bb71dcd9f386adef3462805410c47e926af9cdb990a53bf3b20127ea28a3e45eeb49da49d5c72;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1e90bf0426cfac970874ab3453f073d95bf171de5198f84831df65aefc3d7fc5c0cc6626cb2ca4a07ea1f5a8e421fc39162711c204d04d9d1a8b8bb9a47caf017127d0ba13d40ee954f2e6b29c5ef8170a67aa745069ebbb5b235433693e7109c8396c46539301efe1eaf46baed57829be841eab42de4606bc9b3515f37910bcea97fdbe5c9bf1104e6698640ba7900c3efef39344b967467a87537f055dfa80d009fd6c6f2f3e9b3472fd36948bac00e4951a341185da4978144dd8083f8a0bfd2ebd216705fade086b74e9780bda37697d5fcaa0d04bbf5d4eeda74f252b46c4bc6eb23a83a1253fc74b5d1b1190b432d9523b6e3e5262ef45fdd218c1f631a240d717092553ace78009ffc9ef677380bcf384fa288738859ba676fa8ae52d8d22ad79c0f297f0c1dae4568b6f676bff694eae31a55d9fdc71b11885f56b3d84c1b43a627e57eee44cd95b5c70e7ec9047ed9d789faf018c50d29884d8c6c84369418311df2c43284bab1d167a991ea13ef87f5b938ceed46cff14d10a8a1c16e63df98ba9603e7827f4c0d0423694fea8568982340019bd415b98d55fd30bf70f4c5d996afb845bf0b1d18cd8519cce2e6bfad0d7485f7d90df8ddf54dbc6a8523d501d3a04a26c8c7cea6c940a7b95be335b520aca128eddb479fd08ac6bc6db2b8ebd2757a8f2826578b40b6d0cb1ca8479103186e55a88de07f4ed67a89dd5cf53e323f64de1528bd3a964442b2f43381db7e92d336a4d91e957744b25b13a66bb868d69ac4951986256051fdc57fcddffa578a8f4ba171a93a4a29428dc468921c724f77545cc41e8c9d4482923eb6d06f779e88201215eb014795c42e000ecdd5b80ed86574ef5eb545358e4b25563e25b63b8e2c310ef8f3caacc2f2448bc5c6ad714184fd6014d9b54426e927d00f2f0bdf115a104271f39fd9b100881d32761cd8b808a6aab7d11a8c976f9ea933040053fcd443028b2a9f4f86f0fbaec70dfb8854f75c942d94041db1ccfa766e9c38c24b3edb846da4d241510d2c7e3a8b67f5d2843809877d87a3bca4ee896dadf558fb4e22853d2fe51ea887e983a495547efd22df8d79856faee5ca4ce6fa029ff91d82e0e529cecdca32eb8f154e0bad954644e0b63febeacc20eb13861f1d5efa5b009cfd946f62bf47b20812e706a822d8595bb701f40a15e4e73587ac2ed45f6677ec78ed32b3a03c93ae796d9d9da958a06f813d016305e07b4bcc2f1febd7fbb8d2ff11c90936e785fe6d31b1f7c511318bc477fe63df7e609325be71e2ea4645869935b8c59e70feeeda6e70d5408dbad11f1e392e67fa0977e882e1345599956f52ecf4d59537355b10f34fbadf8651f0b206a614daa3e2a4df46dd7fa038658538cff5b89161515c29a8d6c5143c8a94681d1eaae4ab564b188bd286deeca55d52ec9d7b4a750876fc5d06b35a677c5c9beb8fec9c100d745850835dfd1e06de2b91a8d2f0d940abbd45b61265fcae1aafcff8d2c08e423a1854c7fbbc771a12669c8ed7009a8cded35044ce466d93509f2fa61b822d13bf42a36adb103d432f218664a152bee334ea056e034cb4b568a36b332504ac5e1cbf563a4dc5c1cb189079f37b6b2b25a52efbdcdaf123f459a95605511df296ca44c20f25bfaf365fb25b71e61c2cacfca7c2e86439c45bff8e6b9ef02e1f006958db43b982187f3ee34933aab76ebbebdbc917a3180691f8c11d48794dbd01a7dc2765109925e75642ae67c08f7105a2eea4fbb1a508c473e5ae995b21450d6e5907aa46e4dff5dcc9e9d1fa8b884f8d7ff9473d6419f53e5cb4f0d41cde5879b18b42ea129c74ada3721f5db3501b089ad2f40a87a661eaf7337217d5178e55241636c06068ec7effca3aaed68d397f6e8d3de407553ad0b53b54be55fbc8f1892d8425a1642666c2d31f216fa6582bccd370acef9f810eb461f33105599456e85a338e1e998c54cb74b121e3ce44ada63387a7cb9224bea6611d9ccb943763b93a045f3fb28fa8ef3ce336532af2a0a32cf96059c06806663d1ec4f3346ecbd6307e272c269795bd6635fcf7b6e8a39260db3bf05e9dd851d289906153c48f02ba7375d6a981ee335a7d03bce622f43b9e90b89440f8eab719a66fe7608780475f7b21b857e7919936e67210874c44ea9e91f7382c039fdb8697f5e3c1aec672be84b5480a71144ce20f0df8fe22b4b9a798c7b2e021806811eacc81694c884372df15d5a11b9d4e28c21f9133ca68d6bf756bc92ac6cecd41a9637280713beab47da5e3c24edcccc16d68f078bae9e1cd443856701d2a9e92292ed4eeb7844ef30edffc82f0cd21733a776b4445847433c203e546a93d7923d887b62c8bd5973bfb132727b3677fd6f1d111b006feef87c786d14cd83a917341a2c78ceab90bc32914f94ab7365437fbbb8c69ba158dbde7c2d27ff38233b8a7269722b081c158971211e154f95210cf71f1aef1fe46d201e6cf6016d39ecfd396b22a16e0d31a1c1f290e4ef4c74374f6fea1948b42a5db8d95d5f5a028b13914ad625fec126687da83bb3faf263340c0c634c58abec8d0b2f828c32cbc44363437d1563024d7ea5766ebb5a5cbf907adf708381a26f58852deab396384d7ed39b3c6374924b22447dd2e98ac747bff36ca1ed75084105ef2bf65e89cfded9e4aad48274d0f63b0ca4901fb23f229199ae39de8dc9ff194594379bbcfefa6655e53355d0a2c45b7d380954f520c1aa5814401cfb606b5348c66e0f767ad1ca671ccb43ec873f0cd53b504396356f7feb586c939a17c15b4daa90b49071522aec32d6df66710d797fdac1c277c07262058e370e30e011deb6da4fc8ba5ae2aa6900c4b313d0b1da674a3ac5fb0168890ed74080a613b7f8bf85eec54b06c444038231d96e33ec54113135b7a1bf10b7636e5d6d1b05134b810960dc028cee0559592a9cd23df11b9c81dd0baff07b50b301e914e6f30696acb41c8d57d75983901b1966852b19e5a1dc9ce574c678a9fc454d9ca8eb47eb7a1a689b18f4b2922a2399d183a9703dd1093ade075a19bdab0baecb3440e9f4ebe9a8ab39ad5f36f87cc41aee558bd7532373d98551a7aa55de914f21cf1664f4f6e47b602cd90d7aa93fedc03b8d8245f47fb5ccf086466af9c6860f85efcc8f75d6d4629fa3166f42cf121f9e8210102c87583212a735861189a01b46fc9c3121b80437fe87538548d0c584944ca6653d620bda5a977870f58ebd491a1749be9d82ce43e4db3d59431ca82ae586cde0802b6fe9b947797d62715edb140593985dc5e36ee0a96cf77647413749ebb2ba4d00f1311f1648d99e68404f8a18adb9e5674b48c8867d81be05c8e22b95b2b1e9b1420db457cac2111c4600f70025c8aa2f338a3dba22e117d9a3688b615bcd7be91a386e3d0080192afe83cd542c2460c12f3a66e583e96adb4a09b2eb754a1650797431de5e69629066b741e5cf24f77ed91b1fcb9ccaf2df3e237932c990ba3723bdb97f886645de1067b688e06b51aeca3c53ab5dc448aff6687fe9e8b1f43bd35a22a8c0880c309a67daf4c267e13fe93c0f30040941a39f11b1bb1cc03bd537102a96757f091b6c2b05018467b003920cc0e367a0e3620c8a2abab3b336bb83c3f373f1cd083d6fad1fb873706e8d1af230cc4d5b340131734dc32629b54efe0ffa8f3c98f71ffd08c1a77cc5df96b0fa385c80ff61e9bf3cf95785d88efb1873882066bd4cc8c2716dbd323a850dd8eb8988a406ed20e3e7435aff8318d5bca6047e78a37a6b67f00000bbbc6e588d273dc39039fa0d030490f6aab701efb7e1f7f6d31794fefcdcb0620484232215eb9948fc6e4a69a4b45eef8ca684571cca40591f947fc759085ae74f91ddb202fa6fcf8b0ac5355072ff9a6393e77360fa1fb085b4d40437af95464c20d25ca59eed0718e7149a2ef48a13207ae72d68e08310ddec105e7a95fcc95ccf19cc7db7440b5c14f0dc0003931a332383d56c4f42f173e45618df8bb34a0234c1ede608d1217adc56b3287df1e0393d16a31d600550c2a80cd57bcfb125726c1f284b7cd6c2139fc6b5596a7023bda671f70665569fc62a4862e0d0d916659e2893ddc419bc6334fdc31e3fd44eefc4587cd0b31c861c36195b16f5d0c983b95075efd533ed3615417479b5f7207e85d2f97e406cd9910256675f152b4478abef2e8a447eec207bb556bc4d651616e3379deeffc1781300f3bf0383fe8aa975d0fdd2ce7bee21192145ac4401831be09b474ebad74747550d53910d15e318cce491bf5a06994293381766bf1b8c152de3424b05d7e6e74c49c009e45f64d814a1d993ecec683c9952ea67d89019eec927f07011b87a373c3470ca31aeded9a15d18c43099551711c591f4e33e95cee6f33d80f6ff270b2b4c474719cf0159c8ac9aac714b8b47171d92b7afdfe247d4ec733ed8f6625cc577c91fe2ee0d56ddcbc9b1d66857d1831f44d7a39f08c49fb1639677f6949b368cba196a94a936e82688b82045fa519228c2da1b318018df6a73f3aedbcd95544ac5935435842146fbc623b6652eade30713a1aa4db88a5884c1da976c32732c891bc2d5e070bf91f213cdc81a3426637cfef09ba5953b95ada86bf41d2189c832223e2750b2cffa2e5c904b21f54ffc7bbe0b057b674aebc2df614b007ab48950d296e87533d9f93cb896a582db7ea5d2930cc7f915a1a23a117e797353b5b8043f24ad1681eaf5d0c90a87d581386ebe2f9759d5e52f647402720fe9e7e5014b1f6b42c9fd08c437908d84e804ebd8fbc6e59eb1be2fa97d41c1336cfd8aa346a371e6e8b5dae31bc3c5a05bd6ab7274b904ba82725056cf7e26117204779c985b9cc17399cdb960dff7a4936463db3e395f004a6f6cb57a782176c25f191070313729f13eda3eb6ccc1ac46d711737b2017b266e76c1e231c9ebe9040edec971c6bf4e6ed2a84e3c2989c75102fd79738e43c63052072f69b167a55d083363d97ff7bfb50b122e8b099ff3947e62ec4be60990bfa523430312012144f80a87436d7ba9a6dacd66d9d90dc9f57efa701cd9fa0d8188ad0c31a6b3c2936258b59d7a8c967b59a68921828895979f4547d29d6c56d34f5be02c021940e2cb71d06e4f319312354925855fe55bdc105865a3f69cd849cac36b54510704dd8e8bfa3b856d8eb642a7d8e11bbc75edf7de35f89cf4018fb11c27be49ca55ef2b87ed07a9a754f1bc75cb61074708a696b74a272f37d9ee26ff9ae1fae5197f70ce1059de9749e599c488340c66a729b3234a2843d061d01065ed41bcbaced44dcfc26e841b42fdfdab02f7e45770925c634e11dec24f4094c660ad2b2607f7b7cb7884465fa235189015107ef98e32782fd1a9f4bb7820fb76d63d96886098bb10b34d994ad4ef628233f5f061c3c59f48e5c2b6220368bad627e98c12f7fb8545422a6164c4a9510994cb510cf909210c06e44ebc9febfb398f5e24d1a07c2cf195082392c8e15309447294a34ae29f717cfeda3a52afa5de0b91f0fd34d8f9794df9286590eca8db22c5d5e81193d60282bee078acf7bc7c618d39b76da5d01ba2e4cc32c3339708e8adfd2c8f944186c5ae8a406b21c0282e47c3492eca0b88981bdcd90c7ac0aa1e14890698f6828fce39437b8dc54ebda8f440fc80a065d219172a3ca666b129f4a4794b261f627b22231848ba67fb276d3779e20ba7f321c2d37cb05aee4fcaec872852f9691e4765f918d5f6d32cc9d5fd60bc618a7831e686d68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h1fed8c34ffe540507d71c52c25a3ffda3c1ee7a1a4b341661e2801ca01dd64ff9f0e02b1a50d66f4cfb88e26a904e9571dd320b14a41374950f54148f68d0c61e2363b204a7b2db4d8f23ed149c4fc5f28be6e3277843c10b107114d62391508b3c35d55a8e9a927f1eaef990b05943ff80f8076c7a1731c1bdd02b9945c3f0f6b8fa305fa49b3fc9cdd4f3bb5f2216fdc8b6b171b6652dacf9cbae9d8fccc5abb091aab531e5476ee9b8a7d4cbd6bdecea2743b56ce0a5b906b9b7530048f84221971813534c8852d7df5f5500c42a78c200e7941ae355b478b1d345e4a521a2ab11302009020f668f30ea8df20d747dfae9d19ec75a9d4ef4ac577e36787aadb32c325658f3364444a487d3919adc85ae002ee3a03a9514b6b35aadec12beaf9979519c827a3e6ff865ae628881aa12289ccadeacb6f5d5c7b012e70de820d6603fd9fba728193507ffa0097f9c169bf83e904f2c6553c1b8aa2aad97baa9b2b25a4a36956dd7b03ccc89bcf541cc60098195fc58a3a84e68785ef7eedc7ed5b82a89aba43b7d529ddb28d9f7cff7b4bb876c0d462b9f8fb4f3ad45a2654e4088516c2178f466257aa2d8c316f3c9d559117e0ab71e671df693641ee6f35119c3e01742fc25bc43c5f48aff4c367ad685b2dad651091dcc41acb505577f8750fb21a69ec5554e8c347b0bc7fa8e2cbb12ffa7d724054bc3e0991f46d32a82e6ed54c513edfc69d7bdfe7d01b8991a8cadc1accc116e1d830fcd4d1492ad9080e33429d51a896235290d4fbc56cdeabc728d11df50b8d3cba718084553f219fbcfcd2197888b909b250f19183b0b28fab6b4a314a3f3f9fc1b68f553758d05647472f9e9fd36f502fd80c524eba62aa139db1d92b7aef155868875c7ea1763e6c20b2e69e6d7068f7726fed9d21a0b70f70562783da23eade21c8da9a44f64f1a5d1014c7033d4042e681b013fee6ecc20217e9e80517026929d0803f2edcebf3f7bc095a4865f9897a3c8ffa1cb19df364724839b4e505e99abae594ed8b72812f5f055be8c5295cab87da20eb953f5bddce8a401f680695e5ea759f7f9212025faec2c8d39540a41b5209031fb29d487190374345aa4aff04d0c1caded6eabbaa8d8f4e9102abdb2b85cecd2abf9d26ef27730346cdf533b15df80dadf8bf73a88c4e27a0f75569415fab705a6f6cdba746f50bdf63e48ec330448f53284d17b1a56e4d9e2da5ab57df84c0d56b1c9bc14660f3739d482b6654c9f835849c84cdb60907e4a1fb15cd314617b94e491aee12fd10d217e0bffccd86c2e630ad5ec61e132fdf589d0bd9428a2ed4e09941d521d3a0ec29ed555e6881c9e99edbee3abbfb204939fe9e220f4c695f6d99bdc676a22ceee3827fdf08847899d8c4eb356b0e93d0bbd1323a97d37314583ef5e97a0f435ec4d5d84ba0ed13a638ac64476588e32601bb2d6ba0d3306351e6466f8240adf3fd13fcd9a3726284bce6c7d21382ebb2a91df991253a357849562d6a59c954ea885c4071862300f4d18a95c4dcb82e807105e7a770b2582ebd63aed90376afdec65f18e28f2dbeaf3e8d99aee5ffb31b8ef477293f8d2d520fc86d4ac9bfa7f1005cc147ba03e7ce57dd80c134f30be1b4b65c45706da5b5509f7221f70ba0a52ec737f9e4acf47ab01af14141e1ce9f7862f74884c42f6370a01f78bfb747819a1eb1588c3d71a6035b864e7e41d2a50322531bbc09180e4317487029d1b4ad64a415de34b10bf9708d10d25eab5933228ac1e490678dfaa378ed6655df6b66de6f1224bdc22145c5e2c3d2d190596c82ad232ac658d5351df0c4f8382791a02d3de901d535b116fa94857498c9949a96bd045998afcf001706b0bdd2c6527936394344ef0ceb5ed265efe9105ef71cf7e26e2b4ff999bc0be5a4c5a4b9a97441c295e1476f9b9edec4ce85bcafb06b886046a8833cb0a200c02d8b78408da71153367c95bb9dfc4d2f8a1d7efabc9c0af69d9c92b630da86602ee7314636183e08072fe78abd931facc9f96870e125e6839215a5b0874cbc9921a9c073f0c49ea5fdb6a54f97c4db1482aeb287e05bb3104f385682c362706aaa4f7998b2dfac46b6e79ef858c9e0d8af4b8ff0bbac1199a0b4a6be255083252c27eac0e73064cb653f6b020185093061b2b75fd304b98bd5b1ff731b5ba098325cfeb67f6bdb9446f607e2c4d6fa33625a1e6167e5e0f29e6479bacd699dadd9d40fc85681ee7f15d06b412ed1439c5545bb076b8f625d2890d525985031f5d6903f76baf97a91d363efb5871a23517c2bb25ac32cfccfb2ff869fa6d6541807574768f67f022dac6f9535671e23651d6d05d4d5f463bd1dd6a9157ff5adbb818db0ec62698e1f83ce12daf7edd3be6dfa37fa8d5310671599238b7043bbc574a42e245b3eb830ac15c1c7e26b24d91518ccb278945e1b407249ee570118b46fed3b0a5efff57ef2c133418bab45ac7983cd749f60c46a46a91b1f930890289739dc67fd21432144e89928ebe68acfa68bf75b62e259be6b1bf1f058cfca6b5a559ab42b9b5cdb829fa01a3db95c8f641927ac1e08a2d1a06072471e6cc2ec49a37b92c40b9901567e026b56a00dcf7439142c19a79c84b3b98f86c23f50b37d48f3a6b52ed6102b8a152514646ba42fa954e3f7d65d654eda4108c478cb7a629bc6881766f8cfeb5ab76d673549178292d69cde3040fd9cbbcf517fa7045a04aa9d8022f3c10c271dc6d08fe7498783ab76e6112092c8ee6870da7376eb18773f1c46f42fe964aec32d02c13fb21428caa54798c1102a47812b1d87a5e95a8ed88b51c9378d88cd11f44b69a9a8c7ae1d777607b5cab4cf7e1eba9bab4d760b34fd17efa732ed1a3ea4cb3702ece96b7f1277c3f0faefe1bdf8204828dd204239e4d94e1d61c5717d52b69f0d3b5f7ff3523b072257cd17e53e3457f8eac4a7e3094f2eb3083cf846d085dcfb9507ef153d310224829835c26aa85df933e4c51cf7ed38a2100522cb91a18be44ba51afbee143a6f7700b813b864ea4910a06dbc09a5fc2878486da31e4d5234cef9ddcf4b0978c32c83dbed1ca80dbb8c17145f2b71281cb76a00800127c45f072e35a0889ac3545d8a4d47878f57bc399a876b4a806f7907b663ff993e1db99579c19b4d8254325f3b3a6d943e31533a0febb4b15ca758f3508d214eb9bad0b42ec9eda9351e8ceedb6575ca6bea075450d10f3e0d543b4eb1dac4569389293e2e52b96b6561799c6d4e5899ebedfc9249bf6d3bf4b8e63a6200110a68c083837ffdf5d454b3d0d3f8e8894fe0a3fd5d3ff0f8f30ae0242efde5480a74f4afb6ce533f617307ed7250ec21b670b73b1831510b9bdedb9f29eb1295281aa4031c788ba57ff1ec5b9e219a0ecab03450e8592ecdd331d31f06e9f209163e453155b60f5f3fcfc0dac12f4081df434c4b6e9a61c0bfc0d41771824852f6175d08e4ca6f15bc98c25fdbe26fd1805d6e74a592450beee8eaf0d364ee6af93514b5edfd6ea8a77436073e4888d323b1ba342e7b99860db17703fe87f08be6d9ec589e38354460f26d83795c0436df9e2c657d50219feb3f4d90c3566bbb4970649371f1ead28e464e4983bbb32c64e304a13fd68100f22480f4ae7c987a33bb15c435cdb8fead7d61bc76adc2bbd23ef61309651dd3f1bd648e5bdaed9f49c41916b56640c81c58331cf09362d5eb1b44daf040cd3b4db753353920067578ebe5523817cb0d571579bd1d8752e3032400f90cf7e4e154fb3d7a2d58eb19757aa0a167f61414b406bf040b448b59ac35171fcd7a58c218ea85a2ffb358dbf1bbbb7745aa225b5769aa706075bd32a377386e3c317e847a276d2f820f0bdb39e89f95a45249ba72f4da4a88115b9c5b5fea775a3908d5d6742beb810252dc753cb3a98ce26c3ba9905bf7b28ec38db9335d747b343071c275ba525663d82e2a60b2428695b713c6400976be6ed93c2efefbf427c0791a6a62df7d9c42abc4084746714657eefaa37c3c5eccaba05e3f353ff16c68e3240cde18faefcf6c3d9594030e0d5e668c0208e4f21271510e2ae1c0a32ed63caf76510883f59965ef7e52d0baf5e572fa6dfc3466799b802a46aef70ab83ceb3e1eceb852607b9014e8f7af632e29cda053034c478bcd3d6af4cf26930e94b3dbd2c9fd0dc8085d333123067fe1d7b2764e23ce6384367d5c54dc47366893ad2ed2e9378959acc47d6c6aee49327732d1ba1eb0439042e4453314f6bb5cdbb1aa4bdeaa51654efeec58d44865712eed42ff71e916b4d3a035723b1a796be9c9df47413d3e5ff2cbd52a5f2dfe8344b85c8544f2ad14d1462b12dd35d1a0f763bb380b5d8c3e65d8bd609b72b22dc327b2d1a4041297421021a889517ce413f33b32ac26275a03f46a109a29e2b5b99005bd244af9c5c148bf91ee857206346aca7a64bde799598ec947c996ee46c1eab18a4440ec1716a55b131a9e023883b041fb3b33da7b8c65f8a0bd006cdca38feb8a9b01af0c050e38586061ea82f72426bdf85cfa8db1844ba35245d7142127c22abedc9f2b22d4e6d86f593988f0efda44eadf2fcc5332de12edacd2809387e1561dc39f61724161e33fdee5e6f709b5b553367906797b2848b95c61cdeaf8187883b8e06ece8d7d1d663cf661aa601fa2b4aa5422c13d2a0a1536a0859a8164b75362a00f4e912bb5ce1fe5105e3b1be9493b65ac55b3e806a2106a444bf3d559a28c466a72f65243f196aa4574dfff43b702e94f043b8e8ead3df1982a5fd4ec32f2d0f0a4295386e1e8dff56ae74b7a3d4415d642be8250b7a581e14bb62fabb8da0b1dfd85da63548f4a31d1605d9a6d591963b152cf213297104fc48f0b8173eb60e5f5eef1013c60c97f7c51fbcb1ea213c75157780675fc294b4420580181874226463acddcb230956b682c4116f6466e3b94a886dbc79eaac3fea371bbedf7cc40003a9621648716901d9573c61bb6459b0ad0c80a2ffe78c46a0ea03ccafb5e72a6dfcf6b94adb7427c8315b4f0db81d7aa8432de0a161b7e61d9f3d079a61b5eba482f4ad6f82de3507a9cc6063905a1ca9f049c47afd01076a1f1183ed849c006aae1bf0846e0b6b1bf70654d4afe53bc49b4cc3da6b894eed36c2968bd1d5c28783aebb98db356d3f46002cb1d01aaee52605319ef5a56d35bcab216cf95c4e95943d5883af1090fda9445a249214faf71b607b92ea5d6ab7e935c6705b2ed3a2f4d305cb10ffbf312aa847292090e2baed4138064dad16c442655115756e0ffa875835b0724f93e3098d62cbc34a36f95250a895b2a53716d07fe618b82be9fc1f3ba9a10cd3960c7c70b3e50f53ae8ba6c210497b20cbc1a63f61a5c222eb9b549e4dd13d5441a7012618271d79da1fa94490a2a4929fe51b764d79f334b264f130ba0a07c14baf274efadf6a2a3e41a81a29960ab8094ca5a3dedeaeb01691d71375ac432ad01360f84725e6bdfa76352129dbf790ec9d73bcfa021cbc1e7ebc900071e3ed7dc051993081822fd13812ea0de376298c57f13a52b75b773efc671054444b70d47de08d2c171fca57e4066eea2ed3a447a83bab35b9a5ed21760a12aa0538948964c6dc1c92a3e54633e1263b7d40f3f4f4ba72d09f2af7c50ad1f235c1ddbfe1094607c26ce7c06a5274fb7b7c1dacd9204a6aeddcba2d4cbc59e7c7cd0c37df0670e4c64b529fd1e6067f1544096fa476b5836947e746878e3d9dbd4490f599991d62b773ee64c41626fc1d2bbd7d334;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h40b5f63d5cc50d2b69f00cf022a59a564ffc6e515472095b5227b360afa4b732da9e44c457ef96d2d952e91181524e566051dfcc0f0fae23af1a1a8da5445d100f9c7eac8112dd318c2e2e206f6a36ed7b5969db162f514fdd3db2cf4390abc6dd3dcabe2cffba69b583e7676432e125663b7caa6c138a9a40b2223553d74b4138f1dd4510f99c2d599ae5ebb573eb5e29ff6fb13db43fb7a98fa1281b3e73f3cd64ef9a7e4288a754d7768e6c4f504f1737af93bdc1734c742abc9661eaf0584de5cdd63db1afcebc2f26f064f72cdd05f151074b278fd8718b52e428fba47c2767db89ed3481a3434dadce1b5a9342219109f4e276fa4d5713227f4e82be8629fc14608ea742278da8124f7879737d9460deaa54dfd2f8f8f1a8e5e6f1495e9b1f864c499b29adadfd935523e53437493ae334e1cdbe6027b60e5478699bb7d892e23450c2bedd0b651eba65bf78791de4a68d3804ff7e49a274e114cacd96fb2c27c7d6373d100f75d191080bbc897bc1005926f765a82f3012d518313edda93f614ae5a3ccaa777aced17dcbe9d41352f4e8950d19751d079e20326f61ea3c546f35687c346a2bda25b699defa4bf8016da12283f9e96382f900abd0c6f10dd1b2986d83cf69ff03a7dccd1b8f97e74375f22a3ef5f57b345145b41d5d089a098f5f8c52b5def362554444f32e2762b17cf3c5ebf480e7eef8291a73df480b407f9f55a1ab88da929c8f9b5dc0581d2a78981bbc24aab59ac8c7bbd137b636cc8291bce6ce576eef9a87e1729b24fa573e565806b468a537476a38a13d06551d7e4142a41b74a853227d273b7afa6f8b61f01327ae458400cd390257826b95ceee0e6e2bef80a25271b08664fcdb8ef63cb0cce348ffe6f85eba2ec015a886f20bbe957af78833f5e96d4b21abe3390d36f21707972e6d40ea935df359de9e9354c1d91ba4bb885cf168c6f7ffb8d7b7f8246d4caf5181613d434b7301a823a89966df8786270aa9630c512fc3cae1d7a4b06a725a3b84ea9ab272b85ab98217630c759d4fc2f7f0db3466e0d305d3db6b440da77bf3c91f3f243c9bf32e42e215b0370da0d3b979732e3910ad405ef4341ea1beb41c918e0efb10198db95ceee7ecbda1771d8f45f6a9a7c132b00398a950ba81d816c4bfddfc30b40a3de3a73270859b95a4fa805d9e75dfc7cb86e3ecb16961e10982e507b9e3d41108c5cea0619ebc65d4dc2470302d06311f4df12f5f97c4f9a3351d4eada15e65f51608958088b0ecf1c3b75181a2d035bd5d204f93684896e38c81797cb26b9e78346eac20ccaf6d245b4a12b45bd37a483f5eb48d01e081af4388c01c347fbcd38f964f9082a74eca2568a57d5a239285361e3d649d2360898fbca3d9184d28901704dadfba4b240972937c26f27f29c7fcdf36b003ad7cf221cbd5530bb111d9b9aa95c342f97890e904480e2d2ec2f0da9feb2e04b2c52e4cbf9abe37f5ebf20d8427d08e82cd7541e2e4ca8d95a0393a72a7882f08c721a8f0a1a4003f70313f399a4f35423698eece6bbe9f7d14e3ed7ef68269c086a1fdbbe46bad0500c404f2571cec27c001a76ea74d269dc2d38074bba7b3d40b538077faf23bb9611531ea4c7c45186b9bcfe6b3ad80425857413127d5718050d3684341879a65619bc75c341388a0e972468e336b6deacc3b9f1ae2fdb1dd24b432d351a89951dca393ebb36e911062538f18fcc09c6682ad70b63f272de06d7247a093d7dd38f67d05a13effc94349627089fd2f21779cd0f53267ee06c1941175211d0e2ad6fa580bf68357037e2a2552b0f4fbc93f58a63d114cb3ee3e466315c414bf2d474bb6d26fbbf4f0576513cf2b189ff9eb6cfa700c6bae864e7a4d384bfe6feecfc9dd59b5062ce7900461cc81fa8b7c2e38f700f40c836359d53eef7d66d6529c96281f95b9982495afba2a9959e40fe681cc12e37c5d9511e6a8654c63949fe42bf897f3d46b0175363fed14fe010050d361b2350347aa9b3d289c31317d8a9e2c6b9b790253adf077c030c473f14291cc5d1000c0aed444c3f27b26118b483f58e59d6adf40b266d38f62ff221f3f7b2acf0a8d69aa5a37b846bc19bf7d818f32cf747bbdbb1981ae48b824b6f72dbd866f115ebf9b6e24384446be862ab718398c5330abca43027cef88b63b6089c1dbfb659467a8914d594694d13958fe28bb28aa56c6b745f5a77f1955daf007940afaa15707297e8f5aff87494b24367340597f056a0834622c60ca28583c7d4bed3bbc68c47c80ecbc9a0a98434f89fc271bb912aa7f110ec1932c161e9ab7ee4c19fa2fdb9a6c59124e84a529f36fd0af14739685fa9adcf35be78cba80d6e4db5f380f98c366467b82022fdb11fd9781eb02d2e587c48d128070637c9fc8b53e33742480c7e9a02da7e499d628aa0d67f6e68b4967550fd8ef076a91df4727845253579aebd9bfc3abc4add4f7132b5beda5b290d87f6488e08d7e670642b251d23a9b302060383e5d4e2600f4cc04064d412954d3075294f76378021beef04884d91c23cfadf4e26349d12dc75daf5e4a2b5a5ebdbaf695762b2595fcb881d07f9a3e5554388363a32d3c7228e58610dca2ba58497e4fcc1c22f15c68b1f6e3ae5349627a96ee91665f85d693523c9c3d69841270af778a14478d97800a0032cd01a26597c33e3e4208d3c1fb791c7e4c103be470a6bc2f6305e989ac0e68020f9f1f64402853e074faeb292a5c8fccaa7fda0c43ad807a720f7917f42e74340502443d1fac7842b868e8a42c42d85538016a8e5a07863a7050fc3a9fe6a294e84c186a937c59e1c99ef0ff7daf06061e693864e44cac1e267993d07fe1c8801b3cd7bf5c35e2f9d05e0b5216637f4afd9c19223e0da7fee22f22915fb12a3334d70d7c09076bb62b7ebc2ca816d01e29794673348510d9b7ce4ff2d5a7ac1b7ece5f5d86994bab5cfeb6943a78fef8d4adcb42e535287611e7995659c84cabb7f59b5d37d9aa9790f94b4b48f66f087f4411d0d04eb81aed184a6056d3c5e1aaadeebd4b0e87f48de2b7d79fc9457f9469343dfcc90937ead5a1bf2e7569df79798baf999537446227ec1dbb8ac6ca09900f255ffe5d2bc76faf86a632a9a3733a635d5d04596f58a4709f0d22e15c5e1b87f4e62731718b48f833c72d2147dfff0a16a00a855d45a41e09e67d4036b1bd3cb39439c2497ebf4050321b25cdd58b95565225bcd114aa27b34a1f028f01600d0988f80dcaef9d4e1fe750e464c618ffb0748043436d431df038c063fa36a3b4594ecb7394cdbb9b8c3a06cbe14acaa328554224d940063cf1f6edf296516c13871163ba3157bd68b0050f00cb68b5c2c52ffb3402b1c72b5e72fd385f7baf03aadacce804e60ab222df2a1e2804b6bb982413c832d87cf67efaabd07ed7044f704b85bf4f3ea28b7a3ed26061e1e884a10a225da3b172d98b35f2bca638e4db825680a3a8d8fbee85a1d8752e476342df9db63b0161af235a7297c029d12cfdacaeff1a91aed72ce49e7277ca84d0e655d2e263295453f67f94b2f729100f67e32cc4c57d06f1cdb90a96cfba09a004d9b94895e766bb4bfc1e335dbc5ba7f8434040a30c6e8349fbd09d661ec4ec19f6330780e7c53d1718055879ee4c9e5664a5f93748f08a9a6037ab573465cf37b7b0d004336ff1eb7f9ff9ecc97ef3962d50a31d2f4b50e9fb0f9ed5613799fae5a82a87388e5840fc1f9d9fe04a7771a10874c71b814c7f5216b241f8d10b6da8209e6620a36f40a31caa7081a9617439a3158505b4983d9ac5282164e75c8c53524e8491ae785a8f3fbd035e9ad8f024947f5a7232fec05ac7db5d6293687bcd332ab79172abbe020bdd54a3e5405d4cab276660f57ab7e0d747c8bb816f7e775bdec3eca5dee0b96d9b7760db728072d280bd28fd455e007207fd7cf6519e34e80af548f2727c8248553f359549cc012f14b6187ea1642499265a8b9930e41a7bb5182db1e76a430931d475e518c419cebf47aa18ceed07a009bcfdf4d61eb66b476e151d431123c8209bc0edc1d1ed9f3198513275c0d832623241a8569ec98733c40c2c54ccb97bf6a99bf964ac729b2ea51b862839f09fa0232017d851fc857e0625d9862fa345d4fb091ec22db2e54a072afba80652a2ca2786528384216e7b163c79d113d8cde215e4c773896b3de1707f2e0e7650a458949c995c6ff5533e4350713dcaa6d33b1b68b252771c4857f74f36f9a7259512f19f124e75b59f4479faa5fa5c7112fc34c3bb97b8aeefe75bee7b1f3406aa885c1f45d1fd100bd723a62b55f28c6037fd61c2fb722ff509efedbed50c5bceb7764620ae6496cbf06146a843b6246cb3c93a9ab4bc70a300b7ff6d0476d7129a4ef31d3433c58e847a9cc9a028f72105ebafe98227e3bf7bb12e67fea0d5b47c4a97a6c7ede6f374aed328d628f197082088fc406d6a981f61889e2c8b31c4cf725856a6ba822b94b0beead4c404b53466abd3349e18e66cca01aea8776e4c67970b26463e63253947c9f243503fc4a9abe62e65e6a5837a7751bd2a496d5c5e6593bcd793f7ee1359bec866636f5de9330711e2d3fc866e3fe5dba65042a891a8d4235ef8a53e467fdbfa6c6e92f91de8d47abd36fca9c9aee716b5cb8f6ff52ad4df7b93e102e229e2e61b79bbf45c572b90dd03d9ab3875d9e95c9009e430cf02ee92c1a3e82048b27311707f14b20287cad9f6b68757b1de2b21159a10e924c3163d0575d771e09b78518a59ac50dfe8c2737e18e7d2f51659166cfaefd700ec34d97b1debc2aa8397332a04e5a22d95d14a16992d6ad5cbedf3444ce604d424e8de32867ebc4ed8702192b9c69fb3c2a0bab53728bea5874ecc6121741c42c5a12a1a45264b8f498fd146e6037bbf13c87201c1da2b073e4de078e5a2e45d019df40c85debf23f19323c43f24595e39bdb970500ef0c6c47c7f0108960c640f98e7e0c604d0ad862d0fa946a09b7cb90c64b407094f71397578674d1f3c982f807f56f9132af6803d7d9c385b24c639b39a387bb5cf09bc6628a7a4d32d83c964eaa8664fdf80f062c6a00387acdd3e246d606c1bbcd1825b3339f10e095b09e791f4fb411994282c1af8e7f495d8e307fa98cb092eee4570554ba0c1a251138ff4feac125bd7303d22a627329bb3fadc43459147571aeb59f73975f0814fd4e01c5c953e45a7fd75cdc951e2944a097249301c41dbfb5094bef247f3dff8f0a399c9b3cebe8a22c841b4ce1144126f8f63caa36402c88df0986eea650438cc41c82c25b99b4ac70ecee78e7d5045f9102c2bbc08a0135275c21ee4540f019e5e2bf1208fbd38bef3788b0ff70e19937895ea737df7994f423274b7ac6924975ebc88460211eb2e0e5a0ac1bf98892e1c08a2486751649055780fea2ab4c2bc8e400801e5f71be9db8bf65234798415a36ceaf4795d60dbb81767a3a7aa0489da15eb42b4d609825515e05d122933601d59d9bf241d07f2b250439a17a889016bdd11318cbce52ff9c37f787ef3b14506ad22664b179e83e66ad9a02456b1a6b93a7b4a6136755878dddcce0e5fb6c4897bd0f966fadeeb8e5c6cab494ec15edbc83b5fbfe1f23721a2337521102e41d503c5fa2715ad88420e219906dcf78362cd06876bd16317f049972e5bc50f1e3cc9cebf688739ae9978afa9a9277b9b6a8fa95e81f8ad8f137343f8b2ff6faf2bb32766444b04dbc7e2298fd300829f9a2ebee4a7321a7ca9b9eb875ad262c02b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h4d133ad84cfd6b50fb3601bd092dfa1217ecf22794f2c4e39f085bb098ee41ba0ffc863a0d1fe8df0df9bb4c69706dcb24d9b9d86d6767372c2813d2df90785d885b6bacbb2a13af15b2779a7c89993ea61365618c71ca5e0466b7c98a1b082f544660ad937d4f2db224c8e295a7eccf2a72247ad17bfd8635f32ae576a4aa33db2fe37573140e23bc3e2f75f8ae7a20a0f2a65dd56d59e946d438137fee79292b8067548f32a419fb1a021b59825362850212d29df562b3655e24727f38767f41ac06e230dad5f28336be71e8ee8b119b0149b3a4794cef0d65d08fc46ff05465562a9b613102cb29979e81b6f2fcd14669cf296d3ca4359a789c96f7e8792cda050d73dccb46bf84fafd34b150e93b994cda88b5ffee8ef5a60346f26e215c9c8cda528ec8b1e6b56d62a3de1a0724eff7e0893ccfe7446a135412345ef50ea91c7cc8ad83afbce98dfbcbea990f5e73190f11e6970e1320aea4b6cab56f26560c8c6b36332a9b2db3b5ff977ffe2aaceb2cea01de56c077d03347e39743d978488c51785c0f360730f3277da34833e8a1560cae218322113a8a088ced0fce6ef3f40e2d5b1223a08f3d79967a1f86d99aa157c5efaca306cba65e2a742ddaaff016328952d099481a5ef61f701995922629ce54db641ec7004d6b2dcccd8cbcb9da3e940357ef982ff5dc895811c9a42f336bd5069d3d10201e8a2811069e07533869f8424b05b5f03c75dad9d030308f2aa8e7257b9eb767ee96528a9dd676eed3b98d532028fb0fdc12592cf81399387db95d7280760824bd131f4364a4034862e70434d3a7abf44ed37d9e744847b10dd8a22aa40977057f61f8ae5c82f5b1badd3bcb4cf8a1dd7b2bcfdf30c4ef1ceb6de7cb9dbcb942dc11ab19d31fd18c576a4fe99c2b8796845ef114808d8993795a5f9c34fa78c8f27609f6c993948a0c4a8a20a156724bd70d50437ecb95bfed0b5f7c812bf5087115134ec87285e8e83bc8364560bd784d5fd4864cebf9dcb82914bb64173c11521cb64b9d0f263d352575d61c0323694f895fe3c20432221fd223069a967cbfa02a61e66096a20a320d387434ea559e086c2bec9249c5ebadaac7a7a205516582fc012260390011dbfba1e4cc8c4144ee3dda0d0904f7b813ceb170a13134df525f1e15ac6e730d7a902f13266ac08b326ec88658814a6e2da3f8ec834815023a6eda56abbb8cea6b01d857f2e9975ce4aea8e4e0fa509218f6e7b5c318a95e3735cb9280e06bd80a4109d9805129f2d112af8e063ca379b6ed0f83052d258b921d08da02dafc309e50fa3acca342efd481ceb9af5085e4eae62262a09b967d55c370f2cf918a475ff49e416deae0a0bc0ea2fecaaf7ff8c6dcbb5ca83cced71b52d18d267da35905b96e27fb9e13b7b5a382c899b68626f5dd412470a95b82240d74a474d4fd01d1fe35daca64dadf6f3e4418427120e6c09fa15a46a12ca4841128314c8571cb345be3c4127a1d53dba1b738ee286ae2791c92410b01dc660691d66c7138406d754539be92a2032a55947ca5eff4ffdac75eff359e77ed2aa60390f3d982583d60c04f68a2ee149fb5be75bd2bafe1de355ca74929abdc96d1042025b21807505555826cb0bb9821cd7e7f7c3bb3f0fc1231255ea6bd48d3b89229efa2ebd427525d7fe8ec51b48659328153bb0dea2b19f49303a65e8467c55170de16179dd930cd1c9680e25ff049ded65c3bf0cace6b865f9279451057bf701a583314f28fbab6ccac5ff7aa1d894d8acf1e21ccdc6e2958f2f251639e36f7d89ba7e74448990884bf047a5d4ef74bb2546bee9ac9b7f6100f5df26f254d907e0e07f79f87095d3b4de4ea28c4055ffb01b22e3466dc51ed19d38a55d5a7451ef84a21ddfa10fc199d6892bde3d4b30a723ef551104f0c5d2ac0c6c0c00072cc8358e80cf435880a367316a5c4b29178dd162a28901dac9e5460fba0a79aa8690747352a9dad80fb7a368c1a86346507235d164c3e02e64f93360792ba6cc551fb8c56a7570a15670b578fc7f87c7b949a92f34cbc4846cbb2e288c4167901745c8d2608ccdc4797d743e58a5b62cf483b9225932818caee9e3cdf1fed911a2b48dd76bc2b66534c1ba19eb9a9d29414ecd6c4e4031c90b5c7f7c36783c4f02cd02ed45610b1170bd08f42fea420fba53bb45ace4086fcf55ca98985a07ed5c5b6f72bdc22bcd1d9b5bf1d55f1b90960f7b7770d1f196e2d9c0a2c2b4d41877328038bb54e29e144ae80a33d1367904b79c5a15672f53d7f7aa86f58c89eb448d3f597256dd3393696f2ca55549df616e69425fcd6ac701e33bec2a7419f502cf4974951c0614267c08c78d98b0d5ee4db7cd006e5849e2d95ebf0996f4c73ef403b527178a119b47a472d832b143a164331b0360651eb42f1b7d9807a39e518827d064b01627ce2729c6d65af4ef123b4e5493b6bd9fb660f7b75185615ebe26b1d00fc6ec9e83ca28eacfbed9b3fef3a1d11e6927001943eb2a15f56ef59a6a64f48e28776197a4322b800a27a5815fb457e419facc793a72f17cf9f2f483245c6273a9b40e136f3d061e821b86c03d4980059ff233c1166aed78814f3ee2bb3aa1b68390934c6f5420e42037c3d3bd13e3b263d61c00d8da2ab47a0776c236ef43349563fcf06bb6419bddf956107f4a1b1b3353d8ea6f459df9a37975f351a1ec1fe33d4861586bdb46e1a7a20f40ec71dd8f26e4dbc26cf7e22c0697d767c372115d335d18fa170eb118700a254b5ce2492ba1c558baeb2c8993be546b331188441dc6b0a96e54c5790f48674b7a62fef72d8a4a0124a2988cbe4e6d205f04ecab1a0c4bd18d7194e6e754aa8a7385188c9403760cff5afea07b0c8b9e6597f08045577ed919705fae1460beca04f2ea6dfed3959d36f54c7b3dab451e03fffc8010011ac83483a09afc4efea84dfb30405b11d3903849fc30db1daf173e71b77a5fbb636b33ea278f527c7d829ac6a913326e3e3d8b11303ffbfc83a488f5d204fd5a03c61d1944fa9da1faf7d8292f58009f3f954d46256143908ed818cbbab0999cce9c3b765edf92cb517be04e8c982880bc30690ac82259f193562487bc1a3da7b5cbe576af4390fc8ce4afa07e9aaa4ac0393f48c2b9b27e1e23cd5815659cef76f27700f3e092fbdae34063d7af6ee75f8e3fa06f7dd590756075fdae3eac5d8c32d6ecf55097895a262cdaf9f5dc7a3b18056650cb254c6041ab86875e881b9bc432845447704315cf144cbd9f8097270ca42628573981ae6169508398f128dc89a18c13f4173c370f86bfa9756bb1239339aa5646bab40150bea779632f7fe3eed1801de375f3c3cab43da006c254a2fcc76b85913e55e3d0956b45e9a85281e9acf1207b5c35fa3f89891d925118ca0b55c82a29fe7eba6f2691f1120059a0a5856d529da667c28ac75e0b5ef44afdb042ec5e2a23b22729f658d1c43b5fa8df72208d3f7332ab542f477006eb6f29489a41f795e50fde289ace9edf971aa65f06115717e9998f982ee9d49f8b1dfb82fffcc41964a3a7678e3f45d7904dd4f2e01f970d2c07026c04356040fce8a641637615bf348d37e3575f0884aa47ab583823248e5f07c99fe419af43c892ef94ca39eb520db5c79ef151ab5fc7681426f9b19f0e60267057a360bbbfb257116225aa11216514ab2b3500bd413529347929793aced307d39f43c274d4e968193a8fc8565bd2e9b161c0709a58b051ba2610d154956a2763d7adf22c67310cd6571adb73a65de0ba9513788e5968b6ce84c706f91e899e2f30f296f50ed7144b2c06817dedad20799033b6340de21d3c3838273c962f03ea5a9ee41be5f80d8849ae3397a105098471e1fc1a8404fcf87bddf4b25d649c092b17b2c5a6145709ad67e4d0569477a6b3496e9f4dbe97eae659be12be25618d30d53f1fc18e252b3866c012ab210b8e1882b1848d743e7832787de72f505397b313691e79993662232d54d37bf127155394a5db5ae72568e948c6a5ef880d7783ac2d0003ba59a328edcd67b6ab30ce42a96fb47884ca04b2c41472420a96b3d389dd515465b0fba3af35ed04a4b2db7a93fd7655b405cb9e0fc328124433140717c6010a0050634f46136ab74804f2bc28610ef9e9216bdb68a0049d03d800a911781483d96995fbacf67c0479a30d85a3165173990272bbf2f3f387ff107c010549abc3b4ba8f68ce4d61875443bede116118306c030c9a44bc9d53d6f3b00d34f6a95a116f86b03787bc902969bd55f5ab778f0b97e96fc3d08f710fa731491db717b80958b0b29f9b2eb60dcf76d347eb0b14da4072e03f69451327a5e90b4b32a8dd6ee071c48718a6cd83ebab25cf0f5215c0d2124ed2bc296017f1f983af3aea9408d2b0b58829ace8526844c3097699e16492afb1d6484120fc934998bf4039f4f4d825b65dee39e3403baa4ce4a7ec5945a066a544833a951553fd99a4c4a4bc5775750d2c7d40f330fb529032806b660669c13d6512e75ae06e20acd05eaa81ab4c808f9fd891074e734d7c7763a23e134ccb9060d64b9f9388037b6007acfa39e64bfbde5107056efa20e707a4bcc0017afa50e8a018d17697a6fcb0158644714679338fe068135c6a57383e8c7d6b27b46a0fee604ab11c630084f62bb55e10792621e508a3409910b8625560e29975fdb48a2d13052168ead1f22affc7d4f0404c12e3bdcda97bfdda903335e96bef48f9db702d3ef3c3dc303a59a4e81d06af693a8a3412ebad6ad4ee623c8f52bcd176f29bb3b4ed3f5450e364bc60aa5c951f447e63ebd02fb8d2f6774438fcb66b59748667ff0e6de329d7782a330c1ec9c1a0a9e6ef878d7701522915ae394bfb356947084c02ee99292dce1d53e0842c6603a3ba7bcfc6e049981dd99b08a4590b8c97cfb14db5b9669c9188d723686936696f26a5e5405bd25efedd1a8a520971c939dad9a1679b9f9af49f7e27fb3925b1c26676cd68598a7fe3a9add764b2ae0e51b11f996afad644afe5567507255c48bf393a24eec577cc659c4b4b9663c6ebce09fb004b4bac16d2f6ff677a464b6cfb9050b5ea745bf779209f61e656f91d3bee7f37d48926bac29eef2d87bb90f5019217acd6ceb91733e8826c5e2ed6fbf34308b2af738aa8e3bb91cf37c21416c3ce1e6a00b990758a07cf5b07e6af008a5654b51d4517cdfac8e0b9811ac3a400cbefdb0b49f5c9fb96b7fd99c8e3c73c9007a0f02213696d43b583bd7dca4fe760b21ae2d932eff1aa847615aa68a4c1b93d5634c8b317b1022fa6cf4acf9ff85bad270455338f58ef1c7ad6a07329c01e4ee7eb97bef0bb175c2af24e47f90f83a4e916c833b920438578dd38ac09cbeb34cea7b8f07650b6f86a8598a24b38af4d41991989045c72411b6d0d2595e923db241dee1a583243ba3b943dcbf4f65b341bc6484e3ff4846f3e76968edd74a92b2fe6f720299e2075f8b0a3ab4a3b56df38faaa9388d6ca9050755ca078578b57d352862f6c2259af12f8d77bcd633b8a98f00b549d2665091a499038123d420e8d0aea76c4658cc9c7ecf5a6ea6705425e69ec300866adcd2ec650466657075752633d75275d4e1f1c643020dc852c4ad55a1ac86c1415f1cc26c2663e564144f6be5e6aa671e8ef10fefc89aeca22f70852f4dfab6872b45b364a7a1c87cdd7a5659d2c79935538d3ba84917029114fb3bc5170e172ede10a5ba207de5dc992ffaa1efc391f9aca13d8d578770f461472fca42ddd1c66563;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb166a579d0e6fd9a0bd4d4d38a812a24a341566471b884ac5ee3d5776d4f9fd3e819487184ce251460941ecba9ab6c45ff26e48d0459d208f030b255f230db3e4d9e3040526976713456272ff0ce8a40df7825d3902051d5e706dfbdbed8c3c7c9644fca56b294da306daa63428a87cb751030c3917796a3f4b6b6fb15854d8d3af30ef5083c7f7bab1c3b5dacd00d20d4f8683c04d61df898fd95234956ea60d968e7c87d390736da85e558fadcb6f2458db3880e305cf073a8e34c7ffeece0508b76c04c6d5e401712090b47072a452a00697e5fd2cbc4cb8a2d47a47b0d61a811f5afc3e1b034bf73b412e96c405d650ba22e3c2f3fce993b51305fcacdcac56a6f03242bd2ff93ae61f67af7ebb7ee2d89a8538ee7cee8cb8c4156a7305b1ee08a73f21294fdce062f73e8fde7799075cd11d607090d6fbec354b234d1e667447dd912025ddd819e386ad7df0c1ab4e0c876a2050d47b800c61640c5e77ff01cead1c66fcdf9246247d85e10b30d0cbf98d01df47ab55fdc80a3f4188958e1033372ba194a5f3adf535a89c90bc2053d2f938725ecc3b9f69709f921d6c10f3da42d75a114ee166e6eae2c030ee26d9e1b6443eed996b423da6a840d53be15d9c66784bae9f7bac6090794f8c37cb40a163fb37afee2b02290d361c26e78f1d9e8fae5c500fac09da46cea93bcc584995b7eecfbad48503f37c5108c9ef8cbdfa2e17704fd8b39efc41e8d6ed91137108c3b55f7af4b79c3b825cf1b7d9d79b35f3ff0223c6caa68659d1aadcda2a28452060d930e71053e0b6e2db1b0791ff060eab48b81fdab221ef7e120d505f02aa8df7568425d1a597633da35f8649d3f1fd0cef0a809fb8b5e35cef85c5fdf7e293dfa7f93931ba06592769819d40a8019728fa73a1ba2e6c693d3745340ed91272e3a9775f0623640435f3f0262a138668af35836e858da8273504c1084fd08a12e8affe962517dbd0b1a3cd179377c6c26d788ea087c0dec58419ac806290725855f7a5b67273514e5b18e114f58ae4bd8975f1015fbc853519e1161f2c8d58a159ce1c41bf82f204f5dd3ce7e3ed33d8d723916eb0a0aa80938299130f1a29b0bffb446aaf524d433ea693ef900d76da8e76ad9bbdb7b4854b3f1c519be32921f5d2639416907cbc5bb0da973f1ebae33e48ad54ca0d038731790ca70aa2084958c2aa8739ddb5ed5495eeca38728b17780730df8e1613a6ee60f4c01246738c55d908243a836c184c92e4047d4407a414133bfcda31d74579f80936e0c3bb80ef4491da68a7e7838a51130168fe2419ddcb748ccef15aefbe73e6e4acf61b02315d22a75b57f73d1ef14be8ec481175c665f682ef0aa5b350add7c37d540be918e74c7fd47896ad85ed458a47185f2403248877e4989091d0dc326a5210a519b475f9e6610b87d2a718b65373c1fe13854978cf6ac9f23aae29e92767df3ba706d360da6612c8f963f8f01eda40e2157875cd3a5d68453e1da499f98f144769cf4a724dbccc3f88e49b4405688bec31b492fc2ce729db167aaa22ccedcdedf0db42d4070ec135ec18cc51e2d98ffd5e4b9a964dfd478f3e34b94aca4e7a76ee87186c8f6a1027d0a214c315902295de71c32d862b9e8d446fce89ec94033862f2975c05a023e08fe8f81dda29cd8423f151d3be9d71162224ffaf1cdd70fb41699f957ab5a4a412901da5aff2e02902a2be97f7df6761909b45450408e60e2f8b56341da78bdf6c1a3233eb1c5dc8d083ad76503abef36b9792a4efd9e690373d5da79694efa596d9ee59abcdbdd314d563be278c989bc97f412a570c4229570fc4f24cd5e9656d588ae58067edcf63e74a11951d3bd557e68476674a5666b1bfb6967bc46cd666e1482d8aa371d72416ef77af775ea4200e842438e898cbeed10ffb498d7ef13f4f8bad74375461096d26f3f3cb6c843ecefd91c37988615c3279c660339285034e73c250121ab67d9ff376e005e19080515d9b0f355cf1eabeca0c69bf82216a3542169ce8c8ad116fc36cecfa279214f1ee4b7b1530381bba7bf05468b64ee7084bc4679ac458ad7768a996802264a00895fed54376741fafa61b9271f7e780a50df70bd40cad1e8cba713e1ec7387f94915ad7fb9da3a6463a0eb5b72dac866bc5db8c3febf78161460a4e5eab334610291d9e4d6b2c8aca0f19cbc8d4ac1d2056a05eb2882c1214b26a8e59e25dbab35bfe2400222f0258e36cc72169e222b4443c931d9a4645799c87c1763a5b97be0ff92ee3f0d434463506413906e71b9e203d8a47f4cbcaff77070c205c3d85b6ae8a3ad25da41a1d680052404cd45637e2febae538deda487d933494a0b27244430f17007e722c78b867e3062b56844a538db27f08f286ec9348213871cd313df1c2926e2ad09b5d634133d8c7a44d409b96d590028ac566616a0a0606ec1433fe244bb43b565609332672a0287b58eaa48fae7d062ce30bfc17f9ac9b8f7e195ffb6786464ed65f435975ccd438baa9e98ead105989fabcccdaab5cfa4824c1bf3ea4093970cfd22ea48ee261be6dfa0d466cedb3acc695c55963135c646255bff6caffd5d2f2b1f513c1c0ddfe4dac2b9843fd03573d86bdf62c68c558a579ce09ccc286c207db820ad34bca83cc93df86866c1a760358fb91000514817c1f2d57d28611c9e5b219c0717ca5460310da75d4fef748f6b31718baaba58a3d0031d9f6a56f0a5623f93e554e74fbb4618d6a3933a265ca82a68d421430f24e1ca282c4ca1e14234809f30dfb227e4868653c3c63e34ccf605380d8c69ecf312de5b5df755f7c0c63fe33147bf9f91886b8fdada79e74c13d1a3da1611894e22102a5b24fd5a9fe4d8b6379c79ae304adc4511afcd3a0e0bd59893f3da50f951b2f1f37fc11e0524122f13747f82d7ceea3c577f1419b9f6dcda4dd88dcafaf4352c9c5ff830da80f054936474aae0ffe3fa60ca40e97e0872694f40bed52197ab8d13af3b5e3c37a7a44a147fd882bdd08edac123e6d27cb2d989715766040f6bf068b2bcac0b29202de485e2d37a47ad982319ae59bd7fa2767555f8d9a8b7c29a2b3169fddaeb0ccf632abdb05c65345a3aafa83846fabbc6f30ef868541ef2c50510945d1bd4223edeb3d786dcbbea26bf5d979e4562725e51dabf0a8c8b81396bf8961970dffe87b7e3b467553b7f0e6372a0190abe5f6ded30526cb9960cdc6ed907067c8d3c586161b5588294a814857adb6139615f1b84cec37e0088aec794923005340895f061a1574a8ffb7753511e1746400d6eff47b17812caa67030e526d1bf860d587608550401890bf8d978210a657fdd9bbbb05e3be626ed7e18c1d241bfe0d21c3eebe0b583eb26b8ff9f4c2d33195f30cf81aa4b5a876358119a3581ccfe513b1f55caffe210f0a8dc0efeefba3b99aaaf4175526a3f3afdef2e48ea8374e13725583b1dfae7ad26e17fea51772646e379a10e676cab51df6746f5930116e6c1a953780bb2aa1fa4b6f8712fbfae3b8b5d5d727d8b7bb6cf961ea8e917ec8a3f935fb8ff5dc5b85a8fccd570e0a893699541292138180cdf09634e3a20e55f57ab0a2a85e909a13a4096de20da93f0d1f891d98d4770c31ba7c7c232b0a0c6425f38257e3e9801b14cdedff0efa6e4c0982ab4c27a66d6f32047ed6e04e3821392a1ee9a5324455340ba72fa24956a6427857927152357cbe29c61db8f65c297abaea4e1869698d36e5deb073a95a4b3db33e0e007a7e463e44acb15d252f7355f9302acebae97b5d1076fe824f25989a93290ac0b3512373b3198a6f01deb7f52a5758082043781936a2256e290b05ed53395ba435b9a24cd6fff1483156325942a564693323e8e9815e1ad81015e7bbd1adbafde4912012b1a9b884e4dc953215cf335ab9a516eeb5f598be1bab3675860986604166836af6b20de6d5b56ab202ba3150bcdbc7a1b962feefed1575710f7daafb06978dd9201195a6f1c68eaaf9d6a70dea1bdfca9d2698174f958e0ae6695aeffad0b4d69c73c92d7c142d71b3510457b2c9a1061609477b7bdafcce60cdeedde2af708b2dace71f3356949b082e4d5653fe8d33780c3c26904012e4bdfa6a2c5145d4006c181d1fa513a21a10c38c18f4bfec7d94f69cd0d2bfe8f40ff606bb353f7abc6bd4235f3c98ad14441ba1b566479eebd14b4bd1ad2945a4aa9dfd15e7c7a817c7f732ef6daa52da26c663ad43f169bfa7e59a1020e7756a8a8067649d9d11b8b4511b01fdd1017dbda4a3b29684c12b65e891489b41c7d77119342c6bff1d0b47ecfcaac5b9feee34defaa435129c4bff0056312422ff9a7d9e80856dc36bdb277c1f7dd59ccb770a7077a57919e08c12c7a4bc32ebea3f00da60c12a775e205186c0f21e72336b4e831166f48f6d0312328760d26e6dcd74bf370b58f174d9f3a823b5b3e7e135323108fcbfbec2d1640015517f3637ce6524dc64aeca49b4e63499ac21565463c257fc806bec98afcfffc8687ee7b5da390d14abfcbaafcaa2378c22ecd93143ff4f184ca09ae20b921671c590fae8d563a9a381d4b5803c77ae804c8557b74767f6ac989433aac474e1a08028bb634d4d8139e38c83b9889e5a4babb9da94497e0ffe44de7fc0eaa9d52770144bf2277e1fa992af286be172acd1e4d533b1b92f627e3690e98a05d900354ed457c77a3f8b930c0c2469e4fd050e87009bec03f490fd095da41c147ee3699c46ed3c14b831d5476947f4da2a22dffb9a1291948694c2fc9a5a0368b2378898134d3780d84196fe4ffd645d2e29120352faab29598a31f0bc25cd11dd6bfe72cfff10108ccbd44ef596b0ada066260497a28bc0d3aef832af159673cc9cca8a8c615704414c58c1c1ac1d76ed67a268f59db567054b5dcd94fa04089f7dbe40bb1f1a6b08a335a3d6aff556702352e139d999d124b32e54142f7853650696fd5a37dc0f54dc68e6550020644aa4445dd31f015daf53b4f6c4f02835a9f73f77537a15da92109143c46844ed1590b22fbb4acbaefd843df64706ec4ec9582b81d7d686733c4b3d3d7cd6628a7babd4d70fc7e56ff39c90cf0b50598b86d56c51566ca1f72a2d6fcc21c624ccda8df12fc6689d22ceb26c1c3966f8048ec5d70e54123fd39a7c802288ab166fdbd986799e49a00d19d986da294e08fb63145420986c6569e941ba301961f5acca76205a65d26bb82c7a3489490f2677dbe92eda856a4c3db34371ad0bf9b56eac83ffbfdd1f1fea76f696e103fda34cd2051e34574aa4fa93af3a6452e8b0373a86281f204832c92be932e18dc8ecb16a31ee21d57d1404246dbffb9101470617a1b1c23a04fdf9c66ea15e7ef38297f820f38d6c1c05abf50f58d19b2b957606b66635c0890b4b1ab9e6811c791fadb05c5867ada398b93b4947756a62c065c197b3443b2af6fb621b75ba8fe2a99d84fa5ba78a848f75bf797db36c65975ad3d519ca15d81629693dbec9b1807ea990b077a440d98233b87e0c01ec7de6ad9e581262392d730e9a7637ff04ca6d47a392218a5427ae3960ed7c79fa1f2451ebc8cc328fa1070d55295f9b2e2e85e6b192c122b7c77b717038839dfbe6fab158065d6bdb676440fbd1ac3520a38bf7cdf88a80a9d45c0567457d10a45b4b5a2175f4055379daa815e3de50b31aa57ba32fa3a080a68e04556fda2832b144ee5571d6c870d1741f1d5cf13b7d31a96d09b7c18f67f3aa75d273619e532d2cb6f632a87cc1e24ec4a22c1652511225b921b02;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hac12813aa92d90f2807ab9943ecb446b584022eed9eb01658f3b07738c3a00f385b5f98a29505e69228ab0e77451fb1bc13bdbfb5ec62e0cb1f122907bd5b733e53358b1b53b344ad72d1d23fc08d76cfb3e041f4edfb532ae614be9c212ed317dc90dc827a142659fc2c20487754790a1ee19e8190a261b606e2488d3b6bd2810f246e1d1c3b6b24be5078266c8fbca589c4f28d88dc2ba013ff4383764dd30fd746f9f8f6fa25783e848d00f524349bb1fbec6a351a1293fc0abba6754455c4a13e2f17607b4e999d1c08bcb6e37f696c0f3b5eb8cd5064016913d0966833b8183faf962611f8a1c148d37ecec07b57ac1a88aff0f3edcd1f6d73549ee3738ac65bfa6a54dc3f4280958e8e074b795830a8568f768cf3e50abf4dd29e239c6c4ac2a2f086225fb18c48f78f8f4675659838635a11df3c952a03ae857260a08f50622f0b5d728c1ea5425dd41a1a1864ae7027670fd34ed878123ae0478de6dca3b0ccb6cae9cf026c9d2de96259403cc73593f61820adb1d1ef8d0bbb63ddb9327f5fb6a13289f89b756ef36c1c2b99cd35a35efeb56691a70fb31976f2042024252eb73583974aaf15249c570791c8af58c78471c5f513da15638686a5a6f09d096dce931e586a400dc18607da871e58933817c06ee3f762e97bfe34fa8d224d2f072ac74893ba64a5ff37d5e3cfbb0b847f35a8599fed27a01435111a79e3f2018a75f5e3103e2a85d55ff3cb434f9c087e380a145e18fdee4a39d371ef6115bc7868b63e0407b42ee8132c98b15599004e3f9d863dcd44eb9670d95faaed17e4c947a1cf70fd82d7ab2488b12578f61b55c21dc016e982707ad6ae4797131ad474fe3302c31b43d80b92c239c16169b4d9de78b8611e45cf6d531bea6a283b32418524f4da4ff4716b534730109e9f480cd82f912e75d6b0e0fefaa283d6ba8badb0d70e577258b547dd316f014091ecea82500348b48df823b8ac7e916d88a9d6bbda9cfc81a76f7956fb086d7ee074cbe4d34cf1a271a105c833469688f4f9fb474896e4af3823c12f6a80ca6602c9633b7cee0d0488b960b77804a3f94aecc840b5c207ca9ef7519cab652a60c6199c609a18b15a29421209c4a29ccbb2813a135ad9c355987170046f56cfc6cb38a750957d05dc9fd4f3feaeb7e1fdb173e9821278ce81726dcdf59bce7de4d5fe6a93856a4a7a05d46cf61c45d54ac0b8c6949b6b2732522598856645a4e3ed298295a870e1f349a543eea6c1c585a485a4c2933d3140728e58e32cfa9089c747756ef411502eccb63861b932280d83cb8eafac968598fd8583244cd63221ad0f78f403680128d6e20657e5f22c0edeb812445c67af41ef11708026fc72fac20a85558b8dcb091c2dee1d1ffd7b9a0e7c50c45ed826f4e48d3f64574028a0e42276ecaae71abf759baac1c539f1b2b12b8fd6ce9dabed904b8ed35f622667916d8bc310a97966d1f82d14cb2500689ad110891b14d6a6be29692e2c1a7d25c010a3123b7be4bfb9eb9dc85f6478e5e6ce94981bcfebbf189fe997e90b590b6641f864a214c5036f586850932279378d7336c3643bb50b91e50d9f5ff456edb0ed70db73bd5b767973868f0603ae68fb5f8e95baa2fe175d54b7590782d42c14d5474fa5d4f0a11e0115fed60ee17aadb2a4ec9f171390abd3918458b737adfe6168b16a12475f4d7169d7b973a1ef24b3bbcbbbec1c0ab4f2eefa08ee2d9aa4ea46099a1de095650c5ca0b360d76a6691dc978417453c82139bb69b5b2b73cbf36f908e9ae298ddf8ed21eb2d08d17f47c939a2db0b6bff2fda4026cfa3e0e8da3f91d584827bfd38306b14e4aa86bb0d7ba5e17a335e07d794b893041e8fe4a6bb5a81a6fad41db3385a212fd2bdac0e4942f845e0293d474a2ac3aef5b32ac972fc9ee1ff031cc708787d667195d5a42dd935e19434955b15df5c1b5a7803290f4515c3d29d443030997a971bc545cc3ba120a0b5b6c3522040557bea61d3fa03e2665f7bd1eb3ede570948dfe91c87e0d6fe53d1edf74365044122652dd576b71a98121a787b1916d1bf62b2aaa814dbeaa63f2e4605bcdff8773bdd913227a2838ed6c26438e2d67bffd4f2ce309d03209c1e48451277d83e4130c42b7b106cf8f6df76d38ca31e7c9843df46eca664573c6437154ed322aeed83e50bca074693d8ab0a77887d1a5b0a6318c95b0ed280b155b4fdc858b2a0c90ac7d8ae7e1f1ee30f214bfe2a66095a916c23b305bafccc46166d8cf8c0fabf10f9ff3cf2cc5d804dbce1c0e4aa4905d23946517107c93f6a2fadfbf261de2727039f04a35ac9e3095a000593c8379dc394ed9bfe5aedbe3db09fc6895caa4fb3fe1d54bc79414a34f3750b7e211c8394f5cff799a593c1bb7e477826d557850e4fdb9a32d10ed52ee9fa8719e898351ba65b6afeb99aab2c2aff368475c4af37d5ac9add73ca4f7ea859c261f0325a058904169467976bcbf703b910e825f1f7fc45b2fb5e66b301c1aa83253e415632f855e1c3c60bef10e0a43f8db3765897a2c238f648f4ad7fb4eecfdee8c2c37d0922c2d5a4b1713850de7be3c35e0828f52c1e762035607d711a344af52b341bb2df92c58be2fa7f55fa733120ca6c0b642f60026ad4c7703e1755af8e661aa1860713d5b785cc135c110917b5ed2b9122825913918edec515745bda029162ac92dbc20d4b5db3b6b2b52fec97ad03104e39d745f363d705c62267cea8e726ddafcac15f7429a67bc4ecd94c1936cf57643f320bacf29edbd7cd27b758fbadd09ece7d75cf1fc2e702ec42d45727c631a3c05d6ce7d1bd1c9eea4f2c87cafdbbcdca74bd72e80f28a15c22a07c7c93ab6db242f5ce32f06e6e4c79f664939e2c572e87ae922e67ef56a56a23cb27823376c8118acbe71a6362e478327132379a362c26fb87a2aa1c612b9d2f2a82e4b91b081dda571ee65376bd577461c71336edafee4138471635d51a8afa19c51f955a470891d87716cf48631c71771cdc2afa718f4cef746d947b21b3fc4ec0e7a60692e899b3474bebda9e2f5473ca6e8c013b49a3f5993e836e2daa34bcb4d89138010d978e51d74c69502a7ce116ef2f93393ae65ec67abd40dfd37721ccf80f0438b03f4ddc93d48814d229e20590a74f5c2cd82a4a87f591d390cad1518ed12e9d0e93dfec8903825ab432821fcb4a4d479d65d0fa972909af11675101205f428b86963ad1361a7b319ad9c89a52ec3ced051ec47703e7cf2caa3cef5cefd247794e056985aa3f36ee22b6155f13114e355b9b6a2a57774c7b89282e4a8dbd2dbd911c6b592eed35b12af60d3e6cd3f8c223d67ef8e764ffe49082651f8caf6858408cfd983ea70e21917fb2936c0037bc0f3321963c6b0f5216a714112fd91898b4dff3af422c2458f0310cff3da35de76fb682a9371d5fd60b799540eaa9340aae78618a56f9e7678fab14f0daded689300ea517a92553652610ada870ecbed6a23ef696d822d13c5a2fc793e7e111424664deeed5f0d66742bb1c3f74fe5f4f336d62a72d6aa1971581524cdc3949ccc777b906c1611b1b5db56142928269de2c95cf58561611871cc7f0520e6ee39e5bbd4dc3beedb85621a46f96b91ba4930202be909e905b0a62043ab16a6eef23d3022aa6e1ac5fca51c3bbb9847eda8dec61062eb4e306fffecd829892e3b469d30143a5505239ecd374d03f22bcad36b5b6fa3f389f700806df90ed4c869611605057a130052cbac6865c40da51c8da6270f4525610577971a08b09c71318df6f29b41dab486f016f38896cc8b0e966feb260311c29301146e61718e728d1e97e730c022074404c060899fc4d4f3ae96fb0a88ed7b4cd88863640cca1a09d2aee2d5ab49fdc403f8f720e2446491d300fc9f957197e98027d5f3f431c585db216b77ea77abdcc20853c78111a4a4a77cf906ff37a364b7ef0e7539d86c349ef1e1e977a0b42ced66926a4534b64344b74b764293db1e7e61b7716cd8206325f53cabc7a7ea3c856889ea6f91f55cf866ebfc03404869468d30a883062445a71fede2f8137c00b8b99a929089838c87814720dbebf552d4645bba1e270a317c8a94c02eb35b6ff827a4ed8fc917cd034aef99df0e7b4aeb429971707b08c6b9b960ec45c81f90214f29107f869351a96c4d63f83862a2ca0c7f8f1eb186dec207359d6235114b6945ee0b90702f0b0eeb4718269437329773cb5ad597748f77af03090b3bb201c8253c782b9a943eb4dcf4fad0e032ab79ba030fffda423e0ef621b8f0530212fff9d67239b6a8030af992fb8d63b5dbee78ea64ff62611b04cec216f205539f0f07be0b8c369f32882807a0d38599ff4779940861b00ab2475dcfd15de037a99f8f9a5a637a243bd5bb34c95716d004238fffe0c672336f3adb7b23a012f86b6e1f9ef2d67a41c1bad97f5be48132fa7325c0eddb4a6864cbe18891a4ad5662481170574fc32e6e56f04c4543eaa9659d3deef74d48bd24fac0bd418693953d7819c65c5a0cc85acb6afab971d9b673c5cf733361261d22035f43536f021bbfbb483a10bdddb6877ca8a4f56c42ac1b1b428c022fd98fb88341b359372ee7bbd1c6d5aedb683e3e04026dc0fd49fd933088cd56f665507743850f270fbda12c3c3f594c7e3188f3334eaa015f9abeac3a65e0c43e8485b6449ac1744f934bd89d2e5cc0f2df6e1ec4437c9b6fc1f24861528b3eb664d68c774da0a68fa7d5f4caa106ffbe62172205702dc0aa40f84b62da13e6113041a02309fa3b05b3240c368e58cb072770ade6d5593b610b9a288e14c39fdee09e588858d80e14207849a53dd215c21bb36af2a94f2d8730ab7f3a9d5e3979772efe9393470e1301a72b6be90a7ecbd0708220da8304f20557d114da95b7dd4f2fb72cee32764fe58246e3a8337e2e5c3d1ebddde17f8347fcdc5353e736ff1655d239f195243abb4864e5080f9096d6e8ae071e4ff8a60cd7a7a4de318cb59428003028d755b6fda2a0b2beb3604a5c960970f19339a1087f88a271e8b36e9c7d22f3f22fa4a1728305f018d4e0dd5ecbec5952b574642919baf6ed85efd720b793340a528f56b5ff3188632a7c35055ff7cc59628153845ce0f4a1a097a0594d92128e833b46f6a76534330c581cc5b3b55a6419937f43e8d9d30c1160b0d43fdabbd738195bb9a3e2f15f838fc02aea4d72998edda3a93fbd1e0059160f05871f9a5eb2232a3904d511d83a0c68d3af53b034e324fc014956e667ac79c883c54c2b1361a0f33228887265ec0fde48214977c7784694a5876f9a8ee6562eefd640ed7c2043c739bbdadc5299860e656ecdf11caa69c6f2006f2b7ccce2e644131efd24c4e56b07eeeccfcc4d268b9c43b923a8877d59e7d8e91480c4b442ca0d4d6f044c1a5d276d8ce56de73631d6accc51e4949546bcccf2c56baf5f8a3a6e054d8a3b025a59eaf5bc0caff552321322ec7de754a297ae6823fdfbe46874741d457b6c1fa874e7ef266091fc7c1157c16895571596e08867164bb6f35a3805d9a47848c3acc3cd3529b9d3c1baaa4d66373a798742e32e009dd5ecc6f3018815234c705d52440008f152835c61986a6d4c7650e5e4b0c587316c9583a692397e115d439b795e7a5a0296e8e0a960cfb4b7d6b836f912336964377ff8070c8e238b63a35f2b7b49062ba9b76cc27c9a543067c3c8ca827d3a326beb1d270a122c5081d793a34bb41d8f9008a8137da5e7ef57d087b8b4937bf79581faa219bb5ce6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h579957853b88158192015e822d7f3bc48cd14a13498694d144679f97c9f500256f7e430c76ef6d137b160b74d821bb335de60143c7b3a6063a5ebb2b3e233023fdbe9f1518665a8b8694cc425975b9a207697a52c2cca8e904ae9c11d319a1e1983e8a443ed50f8229e675628a79591470d9f70978874d7886a6e95171f6aa5390ac3fe9e7b67b8d2263b585c3b355ab3ba8b23725ac3ce53ede276ec6ace97c3862f39dcf9714708fe3a70198bc9479049ff373a01c16fbcf72267d8ada491bbc170d962d040568b0e05a44395733dfbe49dfd6238a069fcfb762af3d1c0aeb20d1349f1f2e4cfddf3d20e8ddf4118088d3aac4c12d71cc81eeb97a46d5111b9824c1b98e9529476b475620a70ecbb6606ca38a11242195b61b20e8b5aff91e78e9447747f1d95ddefea5517d6225cefb3264c751ceccd473ea8f9e456a8a055783aa3655c9ef203c0339931951ed6fac82767f6e7153242f3dfb9628981c42fa28a2bef5d4a329e5e02149d9e6c7f14491b98eaa55f23b691bd110a797fa6bb9b0dd23d1faac897f8e752fe3eb1b931624df1a9c52f9a59f66cff9ad39e280dc6b1ff51e6679f510f0b599a367ac7e79a371678963aa57e0b08e47d91bc26bc1d29afe1fabe1a32aa6c463ed671ccc0ddfc2c8084d3e64cdb6e2f116e7a3ad38d8f472102210eaae0164aa6312fe6588b4430d988e9470bedf0ad8fc87f3a4efdaa0cdcd865e5044c777ba19c1fe4e5cda36aa7ed3f1bd2c2b15a236f29d201c749fce27efb1e5beb9af81b622ddc324581d650d182a193cdaa84778563c9573928a3f7789314ec421fa5470b2bb31343d8c8e33ff8ed94e243237edffa4b2718bba016802be86979465913d2b9b0f9ed849ac387c9b7edf40ec65f95e7c9782cb5f2962f8ba5423515ed373e77151804df2cea1f4e96a1e61540396cbca7b6cb2c7ec71cc315852204091bf78646fcff90497bdc942cadef28276413b0ab5f6b9b5c626c4cc11339624485de22ac709fd8b1d7c7e95a08c0d9121da70254a023ee3bff34cae7e699a1f99cf1b3c39938fa9155dbd7dfc6970f6403fc1a5abe8a647dcff4c7ec0b751b535b4d41f6bcc6a4064e9559aff17cd24b904c0cd03ffb228d38745dac5f0724c42a17a986f3e6e797b754902c87ed57a317f50660f11b60dd7220740967f483faf044fddc7310a6d0a88787e89dc90cd1469cb0217da8de1717c4abbe48cc369851fed35315b837cc367e0318339573b98b5fe0b3c96426fb3136269b6474005efaa0323c4303e87dee2a36a807b7a981d895ae9575456d108375f23cc7417e18cc9c30a808c9a282d934ae232353252a4353c6680ea88f63f273226ebf97254292bf74df13b3848159a6dc0e69a8629557b25f835665888249acbae3445b89c5013c40a540b62cb6a1206b653fc9a86da7a9ecc5cb413e2684a4e9544b2de1c97356c8ef2ac8e47879e323654fc883f90965e53f9ddb6ad5730760428f4e67cdfb6f2f404dbc9d4eeb1ece0373a212e470912e52c4932d95c3525bea023c998be6d6e9c80b46b9fdaf6f0acad4a22c59abe7b930b2253216911614ffa1a219bd7abed6960d65beac64b24df21b51c7b2fdae3a2cc18414a2868281e4bdacda092cbb999056d66951446aa43dce3945794b818fdc6b739589f85809e3e018f9fefe488c74723dd7d130eedc50c192eb2eb2758f7857832c455de9dc8b41401c4cdff6007f20761f769f5d3bb73fa7ca3a922c95fc00f85b5c654c3cef46d79fb62f5b0574d1cf18c6f0a0c413f3edc3e37f50aa64296dd6b42262d0a883899bf90e9737831f4069c56e804845977f1793ebaf18a69e7500ab484a4e4993da0d1c06d4aeede6b0128235d00de01a239efca5c830986ea080a4b4767fb6b265e65c432ef61653d262580ff441ae76212f51c8463012e9e67a5c95592accca9a9e2ac006a6e6eeac926154c9fd0476516ccc6b2b2a5605f63892850b7b2ff0a1a3a9af1166b3cde050b0384d1ad59302764b1398a46092527dbc5719e6daac0d354a73d0ce52aa6405f9f67fcd9c753386ae08c9bd49425de6566930170df0dc18af178df11da2e591c8bcaff0ac246382706ddcf45cba65fcee02bd5e20419a2497c013e82081b1a68ceef5776cdd78a175425b2848e6f7cd8d8ede7dda4a02932d8dbafe3ddf3dee513c39a8c4261ef333eb8c85e376229ce09f228d08bd898d0a764397d9fdf0a5eba8b58177ff146646b93aa56274d4f8a5b37f0730d9159dbaad7efce10d9de433e47a0004a506ebb252504cc7fb0f29b2bafcf87596ed145474894b9e609e2ea584bd2ecf47242202ed29c654e977b77f4fd53046a00c3a31eb4c454b5c332057d44ce1beb6afd173b694a82f409084aed3c25843528bd22f568feb80eaa2535bd8a32b49658d6ca0a01dd1fd5ab52e21c9ed2c616351e7e8fac19ffda003660dbb5a1af186e4bfe08061c75c578ade08a2773788606b816a7787ed9343e1649471455c3f2c14388e1bb4949ed45c6dc84cfb00ff7b49c1dd587e816ae4a141b712c5de7257bdf0205a9e43a6d2a30f82ce20f095587c64939be34b5d41bf76a85d2d6aa60ab8daa1df48f6c71f7d1d4c97636a774868d8221a493c68ffd4f9f154a64f3fe6ff2d614d747cfac68f4a9eb314bb351502319157d901f2984bddc4382f79b7cf330dac7d83e145ebc490f68f068d29dd84e577d84cca9aac8d46fa15dadcf8b784bb532efdba74d95701b72670937273c30cc13638ed5ac2f1e6b5a242b1d4f36f91fa57e2cf5f393d78e6aebf5df98ca5a7388caf921bfe9e0c2cb37b83d5353387fbf59351ae1651abc917f8e678e4448aff9a23a3176a1985768c2ae651f5c23b83b42df221db6e052425cda89d24dc1f5a0e310ec9475791ec5f06e13ad03d4c918722b6c601f7e259e2bcb66a0635784a4e41702cf656dc5162af057c363b525388f4af8485e5fd7b4412dc92082964c4548c43f02f059f75ce4831c0847253480be4ab0dc1e740fe8964bcfd506ae6fc0dee7ffb36c47ba9c4d42010de1aa3590a0d1214629d6bfb0276d0b0eb1ac2d39f315e9ed520ff07d761bd998b28526670f3074412c926bf48a870aaace9dab23bd902fa37d7008bccc821a0e32a6afa7d8d1bb2ec306b9f458cb6042746c25648e0a6a34686ca13eabad231329b28d7cca26bf1f503f0e51241cbd6aa9807b6667bf0d123d361ed69f75c99df18d2718d770e7a36d4ac01e065f27319ee7ef3a1e94fd8d8260bb1ac16fc4c540a0a1a1ae7f70adce406d9d667de9c911989e04be3b8b22b06859a1cf2e567149aed24a3b24c6c3f70588e164a6af1910aaee7ce9ea1410a9619ab689dd24c2b6663d374f41e5b5e7725357e26219e0b71b64bd0606994019c5f2d0b0c74f66dad871fd015e5426cd5af0a2e3f4290365c352478fcf2f55e6852122334cc0c96602cced93d0142b9616fcfb4fbe69873273bffd5a35ff0af9e875c4e85623a4e2095d39bc01795dc82fa16feccd227439633ae8a9822f3f9bdbe9bfec916b8f5d11db67019863a146afa6fea4795ebc4a4287a4650093aa845307688b570ce374f86c828eb59f419e97b92475fc90ca6549d2c5c82a1b708383b8236935ea26f0de9584d42cf9456aaf88a1d9fe87fecdc5c59d6f49cbc863ed9191fcad69e72d0b0ddf161fde515aa3e8b2f5b046747f92a58f582fb06db451c27c559bdf2c98b2c6dc5f88e6198c92c2a45729d632da40693006b570c626750ac4f3c73861e760cc88017c615d8967320ac6c916682570277fa4178235c8619e0b6d4bad0056f957d9acfb86cc84ad6be7b6bdd331e197ab5c78c3c4aa93b56701e33e21dd290c4f4e4ff0504a659a58aae94c045d8d7139d5daef548b7941d559540741614c8cfd50b1ab4cbb180ade1ad95924f74bdf3c1a92fd348e361191eab8af66d654943280b268b871208672e74b368077930522497bedc0b2f2a4b984774053ea105cd3b4e76227600490a03acd448dcaceded835bbef80bca26cbcbfd44a172a3060f06893a564adb12f9c187f51267d8909e586eb9c846b58a19c8a79e0d55813344880b42217ddea04a89f6dc00a3987c9a6a6705bb5d692e59735d476d52ec4857b5cc3888dd886f85b2cc51e7dac7fc061f937d5c76659f3c9b39228c4e235ba024bc9c649021056d59fee67690d339d2bb0bc21165185db382374ea40537083ec93348fd7a71f23f43cc15f079b8438e1116552b93b255c715dd89e09edbc1e2f8b1bde5983ea7c54aefc082c2c8c06bdd8fa77b89edcd6f728e789b53e209fdfa48e3e40f08f0065a26b1d5d8575852f4b01595f2443a40b4b079a3b6bf527c5fbee4e53dba3d85478d67924556f02663514b93ade37b1a033de7625ccaa1bebb1b2d233fd19c599ff4725e70e26c8ede9143798bd7259c0ad060e8725b3ba76ffeee79a9a3a1a55a1f2904f452be226eef345740b97797c3f1ddb2a81ebd410e85fa9907e662e72cb91c2ddef8f8907e07eeadf02cb978227b33bfa4c8461794138618fed45e0ede3fb3fb2310352a7d7debd1491a770612fba41a255b073ac64d0b7ae5d2d7d23089244daf062cfde142c9a6785a1bc1a76fa447befd7f4f63c131407caf042b7c25eb59b255295a5aa7be3ed6f2621f52cc4591bdb770e9a64c1ae8b3563656bc9767fd00445914a6a71263c5d4f99658a7b2e010c5959031cdc8d0cc28a89d64b123b4eab5424996dcf3b52e5812761d485cce0df3ae771c8d4055ffc75964ed0a7603350de59cde98dd236ed50ecbe38cff8af46932249c8e090c42d9a6522cde6aea513f5e347e501a66d5ac4de378d684a22a228bf53b53404796d578889b2653f1d6bc9fca425a8d9f1fb5da897bdc97920b07e4acac20c1f5b78c961501e1a6410678ac759ed8dfcf42ba3c3a5a0ca7e67e87db60a54e43ac7e4f040288531d71d749b451dd0faf22610fbb293005313f87902299be9a41315fdf05b26551d4c8f15a6859d6640ca607bc427cc3de6b318f88da71d04501735273b33a16b8be471899520350fc87245d7f6a296a52244ce7c768f004c71859e78182da440b936b7888712338762d45a52441c043013c11d69f4931bfe49182904785fa8314b121178b6b8eba22c7dd5514c0a406c762cb84c97fde88e2721eced078f3757786de8fde32b0f2b5be25317e3d7c64f16ec95acd41f236176c799652960bb6bcb06f918a00cf1c5741fd66bd7ae381c252d75ba3b62e56bf48b0beaa31376c431706a0c0bce96c4b081896217ea731be0c28f9a125f62b27fba12c6ea4aef7bed8b1b213472b7cb21677f6cd1826263dac38531b02c8528862265c66d5e8c65b9c4206ec2de1fb3f1fe599e32fb9fc46732283674c16a109dba2e116e94ab0a391cee11fc85203c8dfbb64163696d989ccce5586201a9f361391c1438bbed48aadee5bbb5932fe83ccc2911d2414f5a35334a06be2466966e6169ba342d4439f44a450505093ca22ac075d08c73e75df9bbe5b28ae90f2920fba76d86aa5b46d2769f4ec7382d5e487def94909ad616c4d4d81acd818b3a5da6689f7c35a76e08da4fcc631386d068aac3c9a5587eba1807baf2c6fd662a36c4405c58347e2c989bde32b385aef9c693df4505e4973356903b342190b75cc6f38f7f83ef864773d379e595339d68a15422b1e4d54b92077e0a0436c0886b4a5c6c1e3e9c18ca7bf9d09eafd960b11155b80ca1e04f70528a6fd9be4a5a6899baaed3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf479b87bf9d20a9b1dab2f27a22ac4a52cbf577fc33cb3137df4f9ada165256695af5c1e59e3fe2ffe0aa32689a6a13963a2eadbcdcffa5604e299232891debe91e9d7f4c36ebb8e577a85acb20c0192915e8dc2b4aea4aaa20b9584deac8093ab2186837bd1c933041a1219614a003403b7641d26bf83d975bd1bec2e0756f3e5cb49f0dbeae70f968350a4a5103e95c1ad663126dc5e7189913fef84ead952e519a016c83b3d3b971f4e07983ef2393a446597eed224970247df6a85e60aaba604968f0799f93e0c2c503b662c8b2c6c5e33f5ddc495ed0de5853e73ad7a0ccc30179831a7b0dcd0454b2a84ed2c0cf15e51604227cf0dfcdc112d55bc6a33e8d2e4034161bfd4c825a7c6c9bd4308fd89ee37c542c8dae0d96a69404b1c716d801628185ca7b88f21da7abdde8cc0f82ab6aa75a1a43d2d0f7bb9eaec9c70f0be5099416c699866073bcb2511ed32f5c710b0619c3ca7bce4915f800ed9e259c29790572a956f608f16adf09d8ba49ebd1b28e4693b2a52891cbf3f773e28a0c15c572d13b17e9882e180f1c648f5a8c88d752634b36f41a0369ef3bcf766357611f1ac5d226b2b55a6c3cee08b7682bf593b9947c6d0a3b2274ba56012b9cded705a98aaaa714bb2ec74f2ca1dbb4113e50fa8057d5b05dec45f7917a97df2ad964b28608d01faadf4e6e53049b897a51493a16c828db4a3ec138617fa3d7db044e8893e22a81867088d8adab2c94e3c25cd972cbb1d935c1460379a46c15db99ec832ca6b41bc1a523e26a1022f09f3213981db0a45986bb8cb95d32da133e10a3de3aad7b1e383060aa9ccde3606fba05441dac6ad020262198f22bafc7fdddc0330abd9984e59a76c69b46880f1d3fec57ef8ed3a42727d1a3c4786a95b7beb8212126f4bd01034b553fb6f0871b1d6c74da89c1e2c4060ddc1f7062899d1e210720a2f943ae5f8c75789a3710c857ed6342f8ba461bbd51aabfc8c704d1abfb74095fd9f4cd7f1ebcb354d2a1c0bb15beac877a1bfc33ee60184582cba3dcb1aff396e3e6726d89220f0ffd116857d013ff52a95abf4c628c8d8e6a2c3aed767fdeb51af41e0cd77b4b049dfbb8a3804af97f020c4b5dc0cdc88d32a65a78431fea34f6f2c6ce8135d2bb276046492ec53129c27980f43dabe6729cc8168ea9bb89b023cc74bd69b6aec0b8a8fd3cba1787db61225638a240a36d0c8675e85103d88883e4171d9a861cdcecd061790f83bb5092920a24a96eebc4ac2ce784f3b7180b480d94e9b850ebb8d6e5fc583f13fda57bb6dd0c1f07bac9b4152554071e632fa62bff70a2dbbfd097d9715c37489c62e8ee4bdd17046e0e346e1430df789e26f58351680136211f5f853568ca7aab0d6daf5f48ddb785692fab092e6dc5048ee135bb8f9994cde33ba551446a160137b9555759da68cc971d3beae980f6c58e3d3bc2191ff502b9a4d302b835df78965e2f199f0bc5f77f42db3c09485f62151bdd9ad69e0af0ddd5f4546c74ffd984bf16ea09f89edc50c977a249fbd7395ef5470915c1baabc67bc9cec8c913fc3c4e0ec10874d46a4706300ab74785130a3579e9b7100a655433e67f13d38c2d3baac1fbd55af67aa8d33bbf38eaba618a5fe0aac464a51e5467870812cd9a64037dce3842ddf5419aa8783f15d2680800a46b26f7128fff594087bba5240471992cfa163f3c6ee08889b8d3b3df2b8a0455fa5158c6a39b78e549990c855b1f100430cc2ec36c58b4a3c19b2823af13ab6634051f7e229dd86163859eac467fbba4386aaf66fa01f149fe68077d38ec8949ecced1b055471ca0c3b59fd2768fd0bf9b8afb497ded394945052dbbb2dc356ff216354e169b3c3ef96d28c2aa61732d99ec098335325af6978f2304dcd2936c702e05c1a915bc94455dfbd87554ac3fc639fc33514856d0649f579dcf29d43dd92c21f4a89c430f63f6e49eeeb4e4b1a7a9c14c87ff3da9e3ae1271f3caa1a2d584a7b4aed26aebefac35f68e0d976403282efcb91f037bb3717ef884035cb94bf01b07dc0b6e3218c1cddeb5fb5769d31636ef38b1a6e8948d6e86ce2c62326bb9eca9184c25221ac41023483785968dfa1402e9e07948537518de534dc90b8dcc0e1025e2f4e1fb611d487b49c04cf66539114229c3dbb9aa784325be369ee2a1f8f0f3a88a4a8add9e94d07e71921818a1283d2708880bfa92e9e1e2ac8c6cd0dc0d476e1c49fa0f9a6beb043611199be7371d68075ad4e1907d298f218949fb51b294e045cafa758ece3966e93126714897af7b7b97075d805f0aa1e0967eec2126fa7ddc2ba923ece617d7b535e7140168c1cf1696ea6c02e9a9b6f3866ded415949d5be0dafe887dc6b6076febff655cc925540ad1357627aafd7ee0e12648d17a8e9a48777e9f2da8400507c8845355984b8527d3e85aa3bf73fd1454946a0107dc6a226d09497b4dcb4d5ebcfcd44cfc2a29f4b9ca7808e027ed0ab6c3641dcf3774650cb3275a8689c3ba3fc3c2af0810d4f284a0d9662d57130e4feb619568d3f3d939955d92cc3d0c863ff5ee2bc45e6460888a9cc35ad0894508ea56e9d701b490d7e29e46c207fa76f1c779086830829f03d7dec1576338e9b9a478c96f2bd7a7368206ee4237c4cfc03bfed9802e4983747fb95be2009f47d5142a723f80182bdebd078d29056631be2ecc880eceda30c526c17af43fe231f2fe4836ee5b45334565179c4f68416dea836ef1407b7aa25407ff836551ee3edca974107ff1c07d5a3b0d3d2ff7d69eb4621c490ccbe2a50519e2ebc717e97beffcbb8ee117d14aae077524e51f104d75bc2cb75f1b77a25f0c83a8caf6e0c53f7719cdb746a95988483d39337452020a343fdab63cd8910e967da2e8ffe13b90a4f6cc06bff08146b6578aadab6fe05352adf8e62aaff1bd365c25a15c92e30478f381f4614e113817d933dedce256454d2c089e9d030a5af06dfef47c6cac7533de672d93c72e0eaefb31b4c0430ba2179e0038600b8344efa02bbb964ee11af5612d7dd2da746c3527696c2b948325ee96dbe466da7c5e64d09a82ec602e9f1e71d70e413533963dea5dcf26a3824dc4c399159e0d44905ad77878c30c95da4a3ffa8536a383c3ebc098f4b0e3c2695b10fc1a639948aac774ac3accff5dcddb45e6cd60285b68bc575cd16d07f971a41f8d1f8cf38bffc4a38819de44cec3dec335facb3e664529184dfdc1f6037af1ffc7364589fb548de9ac9784bfbce2dc31a91c4373083b672f14246cd04785c2420e85849a41c8ea77577a170d7fadee1fe9dcb7c564c43d1d73eae8203e0fa91b4e762da460fdf8250542f6b8d96ea1bc8330d9e988e0fd390f6c348c9955fae744df344be6263a1c1565fa17c9007cae674bf2bb8835e030cd07bb79710d572f41e4ee513860d24eca8eb1b0f035981f9caa02cfac5ff5d2eaa76335045a21f7f02e5b07ed47a30f8b0ac648fa852e98217e6c9390e49136ad84d0413b91bdbd516b7904280b4891387b77359ede840e67d4528e3ec5338b9a9292a654d5b89a1479cb959f18f4aac26730a0948d3c7f319368af3123207f739ac38b2194c2024b991811aa72f115da18f7e0e5f038670677d37a042ac6032d6126e767257b1106c8a50e915dbbfae6abba6c4506df546cfce858c7b5cc149aa129adb46680ade621fd35834603c41f34ecc702ab75dd20e0e68ff8762978852ba44e706fb429014dde50200c60c262758d98cec8ba197ebbd0b10e7ef07b93b164ce0ba76b12a49fc3cd4dc902f8d45ad638465c55e5c1b6d95fef95eec55cac2e863198066bc30b34a749c5f4ca9f42506c3ecf41365d22d6972c7940a9df9f325c4940026b2d72d0ce7d4c97b28994f4192981b76d5ffb9d042a6806235928bff9051eb2ef3c892b137e3f0d79585c25cec784ea7100ddb2e862c8797a5b9f1ac238aa74f2faf41ca9d5b5ccbfee4a459f9f1ff4e65bd95f02a17f9d3ff463e4569a0272dfd08a63fa027db610166a6de8918e62fbf9213cda94894ba32a7defd09785d20d2f87a474efe021adb3ee5e0ebadd351c8a24ae07a35c18742506ad9d478632eb125bff111e9a1b7da59a89ff06eb42c8d7280982d59a0a3f6f6f59cf4bb50c016d1452dbfb519cb726e9b0252df792058a3799c217bbf65a3fe1f25279239d1a9fd12ac6fa6c88e6eb72dc00a31b8441acb4ce95c314f2dbcbd5a1acdb81cb38dc1dc81c3e7323f31291366e6edee827afb39bdb0f6e7c2b9e2f8a5abd58c98a62456af7667b06d4cb9854466500295f931cab0f9dc40ca2aaeff31d744b5eca8ee795957ddeddfa231260eece83c00934854c01bf4e1dfb23b9fe7cb0a0a2c2b43d5f5220860bd06a96eddd13d2ec8445e8bb27e8121c703ca3c895e49720e420d8f917a17b9850e66e5c22ce5bc0975299dfc38a8d6bf0656e64d63224d0041e962bb6f3ea51c1fdddc4b3bc533b64a351c470b06963b3461aa31874ecb41dd291ab93b65a6d7441c2e51321f95fdcf2540148a5da8653f8add5d8a21b23191af15fd8d246e8c6359ffed69d91fd621729e31984b016480397d0bcdbec32fdd0d5b23d0f1d0bd509849e0bf8c9b19b233282aa68ef85b1f108c9cf2fdf0303fa136b93fef644345c9d4390dbf44ab1014d3d2501c7c78e59f6da35fdfbd9263a586743143d337027579bb871b1cc1c0ef7500539de3a6ebaef613acabec5031c679963dcf5410a02f68aeaba4d4c4cc31e6cee1ca317a1aec4920544799063c02382e0016b1bc7a0958bbec13a2435c2f3480426b13a1aae74367a93d179ec5b2a877e907090b354bbe694c71beb5c363eb94857f76938526294f15cfe5449589eaf797b169a4b42d5629506f9c93cc549872e9062b49a444073a3a2c1ab30646b41a2d1baa91273176ff9345f6e156de58a0e902cbd645ff3482c6d7bd879fb3772306b7ea26498864e4d08895f7513760d1e3d7c99546a722ff05d9410f2068bd1087e6e20678db82acd39a65262aaa5b26daf4e7ef905eeedb3ff856682dfe1f1e1caa4f3aefbeab15cb34bd4003f1c0a8957e1a50971247c5d3f19f7c5658718976d57ca6acac798ce0dc2bbe346dc612f953240d6e1ebf4b0b9fd53da1532a5ce5da929497fc186f8b7fe9a5e711c17249a853d5219a07b53c6e8999fcc67787da5ef90f856a2a7709ac1d49375640cb513d7ab5d2889797e3fbf2ad89ba2c82ed90c7fad6783d23510b73615e4c821277235abca3a2a14513a980e2a2e7c7e2e7d0103a4b76bd5ecdb1789e2da383f493727ee4f931756d7d3b0d7a7e7fd0cb513efce0a82a35994694179c0411a97fbe6bb3bbe7b78e0450548a0d694e006f242b592add03cd18adaa1b4aa921134e52c9de81d0cf07bff4d9c544b1979d4e51f8d96e363b8ade9c4df4171eb5b779aae800f9fa4ca3221aa1a5c202a53db2ce31c245d5a86acb443d716be7f201769de5d7c6bc3d32e41865558c6d254694438d16606c051793f770f17ebb03e76a02dc493ac7248b29f9f2c1ac31d880d3e4e2d72c201cbf8fad0d8cc3365f5d36966ab904948f6c7dab5b2f379e27f8ca8e92dbcb92ad686a3a23a9ec8c65c90a2d39af4f8a99624ffcab96a53ec5c7a19bec16bb84b6742f362ff152d462e8f63a5b75f96aa1c9c4ed7a17ad330575da19b1479646d414d6cd9f7692267fad7f71c153521ea6ad04056ef8132ae566092de5f38fc8235a9ffc05351e89a2fe932e24a50de800a0e284583e246efa481ef0d8d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h74a7f1778fd532609ea9e36d0c1be772efa41743db96d7194c28e9db8ab9971695e736ac5ee19c319204378ba913adbe34e3b5de05f4300cb7c05cb90970677a6246243b42c50d2a6511fe37bb5fa88b1569cb7b22d272fea601211a85bd8fc6bc7dbde9857a155b13627b2f0fbf4940d286d83c4171dc35055ef766a146628a3bcf853b3ce2d29ca8b2c66bcef6f5c09c1fb4552fe54dca4b29c693c8dbbaf109d0450f1aad692c5002faca1d0664bdb449d5ec51374beab7830ace34ff9e0851e23cc4b4807e0e03b374fe8ee3eeca302ff9ce6308ee618289e77bf4cd6f1f378f82b7027e6ff861bccfa3cbfb6085d0ed9b92a4990eccba76e1a3939c3fb4d5b70ac5134b6bfce09a9475bd4ab33660a0281bc99e58dc83527510aab85bc177a7ea21762eabc2db865e790a4581d2842a44d6d3bc17af685e7da8abfe50c81478dca245f559bd6c18028946dfd6c349d96c49f627c73914f419506c4f53c5ec411390dbcde242ecdab7a6a792931c4438baf44d7efeb27f47f62704d6c961a3d27d8811cf7a8f5c7f31b620453dd40dfe04fe63dd662b20d1d0abcc6f747d99b047e19db1f23fd18e08e9d2f100b8e2aed1de69c6f83152addca2e4600c5f93af2e91b4519410ce9ff2071e3efc9f08daefc06591aa86906bc9ce9b57198f8306cf7188de9f2e074c41814fc4120c3ef9a094cd87888983ad9c7b7cff339a668ab5261eedccf01c9ed40c80466e0aa6b011dfc575c28a1bda8dda7bef47276586075d9bbbb88de2259b40a000d50256ac9db1c4c77949da136272e9dc99ab2500194b2dfbd8f955f951b475fd5ade4a01b033221e127c759af857bd60d4cd10ef97c0bb1c67ad11705562b6fc0675b66531e9ba3fc43c1cdac53c54a00df4939be919a630cfb7836f9de792cd8eee8cf72aa1659995ee91629cb28327b5741795df3f1a3a469200dc5a3f44213a75b50173203d1b266a6c6cb1f627e3eb31f530397e9a32f86deecdc6eee5f4564f7cad16df30cb967835921668884d93e2b9ae226abc6b85e6b1d0336d8e3625907c341440d9346b63842abfc1bf8285617b4c16678ead70e5cb25e9eb088ba19be57cf38b5ebb728d594614b9b442825b4cfa9e1007ac646966edafebb544a66dfb51ac266ee00de8700fdb502276def386158b33f0e35551398b5829e63bdbf99ec289695f63877d1a4fe0783099af0778a1c70bd43651e8d29d96bafa682bee8f03d70dab374169c12085e7d7fd44dd180519c5f40de3390f9a15e8ebc4fe40f585ccd703a9c259e39a9279fe406f233e9e6022d50ff65d4a15ec6610d9af79b51259009d1c2633ec2efeacdb13785fd43ab0672616fc82ddb1d6b918728f229e20fbf8e6d612e3093c93565c8b759bcdc9d93241289ccdff98c4dc74fd1463f5b390fb66ded0e664c1a0722cfd64eeb498e26e8d79be06d1b35ded185a42c66ecb4bea7638f85907070a2df63c5d374cee759d72ecf57f77a48e5590cb9388ed29a36a93174a7cb074772c35eb6d0c15dfef9b8cab7ed558268e241a927e78b0f5e66f0982b82341b80a03936b182fcd3ddff165feb7f18db2d1c0f53e70ef99b3bc71d076c28c33ded98d7fa60bf09ef7b930a441c56fbe51a9bcc9c4108e76f396987abd5159e334eb4a0f2581133570ad3ce7a4c3917f4017b3c32298ead43e4da3c7c45c06b38e243952edbbb6b7084c4b1b3ce09f447b1e5f371edaea349d3279b9f194786ff740a3f2d825ec1773b4d2eacbba97e868e61fe5597f2fb1d9857011cbc599e4d7e2c453ad8d55114ae616d95a7614977845a660bfb6e01def6c5edb0e4a2d870c4ff616b5f1d921cf81c43edb6194d95aa077eda5691eb74da0a69a56cbdf4837cbed911d42ba53bdb09f82473193fb0978276163c7dd951b3f2964106a40c7ea6700389fc4518932fae5240ec46366e8b4e8a297fce9a59103032d49a4acc779a3e3e4cb08d41a757cd3e7957ae98a2999d82dc778bd5cf0a1329625ef75791a1422e27525176b8965dec63b8b9ae1208ec2c93b72e6af21597e4fa4e06d732292175d47f30937d7c2498db7435a0c35a836c6c993ad8bb6ed72324e2d4d302d3df7159275b620aff23aa3547c1dcf14a54afb2cb9fb07992ee9b4c1f29f33fd1d7589460bc4563d404402ccdbf7491207945cb8b68264df46b820f6c7dea6c3c0d63d16bcc65f013dc825efbfdddd85294c1144483c016e8175109f22084aa9588c8099d8d54cdbab6f7ce1ff564a02f2ff07119a8cf3b2112c43b9f9a31dd7557aaaba96b300af523848683f2f74a79e4f5c8479e4ac74d4f5766ae0655556cf1d6b66ce5a51bd68dba7f218ed3426047409e43c6ee19924c22226b8f7b6c890e614535a8671757b9c6560a9862a40d3a738b27df27bdb4252ac3ddd4465ecc1ebfbe7dabb4128fd0c70e46b63a098b1ce617056cbbc077480de5ba470bacc016a801f42fedbcbf73c90bce18d8dddca34de66d1f60572676f0e452ef228d63394f211bba29c7436c195743cc6661db0f512f26ec379790eaf6909a9b7cb6250da1b879e3fdc93613559d02d093bdb0864f782fac4bf6ca3f36e128491fbef35b05cba65abab2856073bfa1c3d663b0a776d5fe15241bcbd8f6d1290a70f30aa301c08a3ae55764d91a86beea245e9995a77cc4941c631cee4f0b0e3d0cee213fefe53e7b89fe53a150c47b8001b700e0544f264a8851304920f944723820ee4c67e07a33b3e5b6dad421db4becbc58afb1c7d3655119566c401dee945bb65700f2d7d14eee4836d169d563270563ba11414b603e5c45a727b235fe2ca0b4b2022b05e11bca2054423d10e1b7cf7d4f6fccd2ecc23319e0f9378306867c1380fde356799453d435b0a042a592c46eb4a11867f1c719551f1e0a2876f8ad0727f7b06827a1e90a52e6cd8988077bb45a4187327676aaf096aa6d5bcde576862be0ab5b388231bef0e0e76518d0cb1aa59cb8e70d5905e654db29519d81302d0620ee9d69db66d4b2296ce23b053c69cd7651c4ecf2ce608896c892613335e3a2dc5fe4305a9c74caf39a2fcf1521467580100a1c371c067f57a27696ff34c5ab74156c48bd5c51f0e81927b95aecdd9d7915395367f5ac0fbeb844cc24d61d9fd8a80b74598799f10c13ac0dd364948ed64e4600f56e9ee4b9f7389da2696da25b6a7d2ff30ecdc0136c0374d0c79dea68b4a48f9f51f76134dd621ad43f85630474b681b37089d0d15c135fe310037291da92ac6b8106da6eee0bbd26f17de7b8cc817afbc46547c4b0ea5c7fb16c8370d7012a2cc09a1ee19808ca289bc4a35fa98840e157f5377616018d31a9649d7e363362e9e860e95ffb40f30642f7294c25a241329cf20f078b778d8645381b296556aa1f5c759df4a8e3b5252bc3e2f34dfd6ecc3b2f311435e9f8b080dacf9581b79d44c1244d2fea1b09b99aa95396952a55f1f12bea29df9973fbe730648982020fe068434bdc8196f750158ec467a189f5fea951346021014786cd3c8c2a5f9973cc50c7e857f0807598c40865d97fbf4b65b4a4fa409af89168c4da64ed3ad593e2d971236e70ef741218905582680eab8809d15cf12c4fc6be797b5a9f57dadde5bcc69198f859bb05c6a7bc12a6c5f86431736c77b96e8896442119edff70c10482212afc67ba2213a45940dd1e494dc87c35bd32e5b0495609cc0ce80ac9e45e067a649c34a95138c0e87adc589d7827670ffd071404e80676e18231cd7feef7d507bb5886ae0be1a5dec1bce2c57a8c693a76e1159a75bcbce3d06b16689bb438fe68e4224eb6b06973887dd4e7366f50956f1338328bb70bf78c34e83108436a57fb891f969dacb8b41e3a7c697bb99e0ac992c9318a19f1f2afb8d48007d40d8a49b0d2b228ea39f6bbe501be7303e40128fdd714efd0c7efc721fae5fefb46f03b4c065bc12a2693c82a36eef748a3b0d186d236d44cd65bc68a9b711619c81e60d84edc02872143e1cbab6d889c54d69b8279c4f25f66366534a304a289a1a1753450dbc8395a7615180b629e9ec80d85205d2c720adb3d26b148dd0d60cdfdf3221061a36ef764e1f8f140498f5c41dc0586d561bc6771e459d283f9d1ff555e2a7d64b0c8464073fd7fa53eeeba38ce6262ac8ece85ac3a7e5a5eee67b37b81078051d933cc6d47eb63c0e80fbe4720ef33d841b2aeedcbf24486de783ceb712601609623bd02b68658d74b65fdf9e0cec81f440529fc5371c0ec5525056d404f128593375970eca7c2a7e27b74d819bca208e61383c1fd22f9317ddd32425c681191b4dd74d40611f7e0408ba558235506a5ac03fdbef6052c4f774ffe7ba71293b2114bbc592f150655c7bc136ae20e06ef7179f97621158cfa23922ccda56d58d325b51959b54ec78b0158a74afde43773bc063a7c214079fdaab5a3fe2a1eb42424408f305bbe195c2588c110cd7b556c72d6d54be0c184ac74c163151df3f8198b6e19980910c7aee39dda3a16faa66fc219f85bee21539606f99a01561b78bab948b60266ea620c36e2a9fcdfec8e4f07d6262a2121153ef6167d16ced6fa2cbad875935a934fe4112c51f7272897f2a91724be92533fcbe34b0127980c867882c1c8c7cb7663e0261f26a2b2954d6d94d1259eb7a31575848b64204973ff26bd509ecca263e01c80a234f03fd82ef9efa2f5302460e9e48fcc15a393c4b560a9a91f16da90dd641601b65dace5b944c22fc0f3f6876c33ddf0ad9baba9e086a09e057c1f550a314f8b339c4bbf44fcd230546eb6fdc7a38a45eefd4d3232fc7cab4d2455a413a997ee4d0c098dd86db7349d20d740a51333bdd5c90d556b9ade0a3cf16eb806b55ef1e7871afc1cf93b69b4de6907c7a2c3733b4c93315f56ab7181ecea813869acd51be3bc0435d369c4054e73e9fa49d9a426108eb2b96def2906895bfa7bca98213edfbc0e37ca886253a291ea0e0af036ef9cfd9ab06910f8f0fa1000dd06e73c3a973dd96bb6d32d4dd96ee2f847d3fbc5e710a10de50bb3d35e94ca22740920a4df4bcd84525a63a1cee9b631858f3f74a3cbd5e960a1d26b4573a6cd874c33005fb210b4a8358af762cc96ab96cb359fe853137edf17945b86b60ec5244d2c57539444a7c887d37f1507764326a14bd7f41c4a5902e3da7afb5cbd894cab22600d00d1fb00731b7d2c41c50d39dec2118d7ada3b1fd5efb97c33829c2c27da97e499ce51002933b54cc0e8fa5ec62d341c2b4e3f39eef7f1a0602a2478a52018b3808d981d0629948e0d8dde6fba4c076ca2231a55a356e4c645bc74a7ac9257fffb43c2b01b47190c6a980ef1473549d7e890fd9dc6a6e8b0a106522ee94f2891cbea665616bb58d0347d789d5337486086dc8edec4d3688255a1ef352413abfd76fab7b26dc19fa40e308c3aee12ffb486d588db36c08f05b3090dd3df94120462863d03a463c816aed75bf7b8158ad85a2f9f41c4404baeaed561bb793146f1da1b48c11713172f43452ab8b2d1eaa6225cfeddef6890adeed5c5e676471e5071719ddcb1c21554582c29dbf73f93888ea530da2cb6f68849ff2373d95904ff970e9484d262aa4c2d2b36c5c57fb7514d00b80bdeaa355731895a9800d1cd1cc73c86cb90688e718df42458023018e55b7351cf6dfe5f08739ecde51e0a7448aa0f531f1e1b753cc73a1bc8bdd43c870b03fb455c56fdffc415862e2c1262ff3dfa8e685735c2518199f8761f31ee7d05a266167dcd4c1f68d35f8825140;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h56d8dfd75cd7f60a2655bd2429969e02e507817b0e19822bb90094f6750877ea96588c98f92501f2b84013c2a07255b1e3fd5c63eda878c638d27f9d7c3dcc8b667c052c8dd36522ee5b0030fa9242e7f21f1aac25ec2417ab28b375e46c314a5c2f4c636eed02206dd445801d8382324c7a2bde983887aaae27a7a95adc934a156759e486a4265e5156fd49294b13e778011625879ce72be6afec2dba31f7f08bbd6b5fe1e4033af04a9465293c187607eac15e40e362f88a52fb84589fb6d2024407d9c15f5aa5337c5a8761aa93a8c414cb1813313d1c204bd44444f2b362868f6e422c1b2c944b158edf77d4dfe542ab45838ba935dbed782016df1311c9b1d901bb55c30d22170798ec5d753974bf811cd64035b9e94585544b156f0abf7c49e55bd0d6b30e80ace9da852935229fc403cf5f13aed71ba4f6759a977ccf68811e5d3bdfdb552d92c8066f7217bd9f60cacec72616fc8ad9a6f84d06015a5990edb7c7b514bd1cd5e5b67595a0d08e1127088cf5e7ef338fa85dcb04ee2fcb51b87c166d05e2de056498764b83de2a21e3cd92aead4c83f3225ef3ec10df24fe3712b5321e9ab1b28ed454af40c7145131f62b249e3021eea55139863caf1122a6f438dc97851adea856d13af166f76a7de73f6483c902b04de73582dce8e70f0e6eded14a70437ddcfd2f3d8537d20716fe86fa6d7b096838a184fc973508dda7ccc3aaf46a2a2b26517f7969d67ec0ccd1560777605e19aa2d7e1d02cca55a760103712910a2c2b2dffd3097afa2cd0efa0dbb500e04b865d794b304b158ca65f6a03f8ee405862f24445160ecf59ef3d8bc67b4bb7d29b001898a14af1dd027e3c650bbe64bfd3504c30966fd83b29682658740b65bcc1bbd89cd6a1e453a410358cc7d55ef478616a29620449af11d8925d71486aa76101b1c267369079f6630ce24eabc3afd5d5a9f2709163d72b7456d0d278d2c8476e7dace8b5d1e2a394d1b972dc5d77300f665a50d0b39e10bef872e42378b97328631dbfafb133fb02852a0690f4969769cedf6cce7c6c942f6cd5c87d43c585044b9e7b958885fd36702e9883302697f6e6005c2fbe5b438cf1e8f6efe7d27f105670cee9ef971490aa2bdfac81967b75a2065e7251cfa373a03ebe3f1b6effe5c27fbaa8aac7e48d7e90f2ad8aa24c510522941c4268fdc5a28acd9ad27ffc11183274679ee66a53e12d6662111462c2de192257358034d253bd3ad2d3c1893f9da1c6aa7a65a0fca6536c533965e334e7abe4b58c83303368cf60ad0199bcc8cd559d358ed54f65776bf9e96174e86c9783cc5bd3e5847c534a3f91dd4c2fe0267a2d08037f97871e5332d78581ae1d523af8386e6a350bc533ec0f209ade98374b3cacc73d2e5c30414ff7d035e378949fd5532314d3a66020a07a4f7c0322c885feac58b95b5407f91b35566e4cf73be4047305ca5c47d9b310b8cd767f4afdc742fc3255009c4ba70da9f3c35b735675650f4e5b7da1e63e04355255defc4b583bed4778e96615c340c80afa18dc14298d1b49aa4c48ae1a64ad45097391311d999641b39a89585fcb51250e7feaaacefa7a384a7ee9cb1b8487dfd6de0d531a4ce225fc57083fe777dc94fd8b3d31cf8e3448eecd3a780ee8ddc86cff44f688ab6674d1508f6acbdb760597ff394ae1c0f1543f5e4d4495e06aaf1ae11496b850e7dda2154afce6e991295adf0d3b4c354406e32ad1266c41d56b67fa6f0856384c19512be885e823bfe398f173575b3440c09f64015bf633ed7e26b89794730aba81a17e8b36546dd2eb29ce2cabe78950b8c1e591a794278caecec6e74ba2db4f25708c4a0245a3d5cae149c24e1f916b849368b928b511223e98a69232a4df31279c9ef20a1d7578e995efaf61d376ad9ad4f7549c3cbc0a1ea7d0b77fe8f705b2f91e3f54bcaae58bd9384a72eb4b4fe19f41ba72051bd6f00922da77b382a1002c5f0565cc45e2578ce4f4b7807c10fb44f6a5bb2fca720f3fc53acc5e8b83a304cb92af87dd79d3670ee61c1acaea1dbbfcf8092f5e55d1d7c1760433fd7176a771a246f3f11ff41edeaa7869f271b7d0289af19da45fefca6fcb038718cbd9b084cff19f81c8ddc5a0d82d2b97c3864ef29b00380ec8e9a394f0ade5e862b6c9c1e8a77e009b95852fc4eacbed00deb14586fd1e26b36a140cc4e37b70160ccd06b3c69825032cbd514c7751a3a4f2946aa9867170f55564308a21b27c93a53f76e42c5e30b2d5768d9c1e3b140ce87bb70c2884eee95a1f358d91b2c756b2c76f35cb0c2325e7ecfec6b8cf8bed3ed737cfef381dd5d26ac27a764811205b2bcff02a9f0964af859ef2de379a9430e447df4f053be4662546650c8333dca8d6ae2d156119c17038f21498f865f4b629f7a3debb6be4e32cfd763af56810639fe2ba62ad702cbb565b0824db8ec5db20229042280eee5fec808016c33a007457a8eec7a32a61da054d0c50fd0abcb1f302ffad27eff5ae468fe91be69f795111b096fd2a602612581c7b5c572662997657d96d159265e6ff400ed06fe9fc6afd75d0997a6c904c4c0b5b12984053878a725447c282f84f82e6f4bac544c09f8df3e63b2514eaa757c30471efbe4f6265026e35be4b8fe1571c6a5bc63cfb57a0c6667773423bd9b4801fde19bd78f31be3dcac05e95862be5861156636f02b1b0bac088cb70591d4638de6082a5b16bd453b44a9c2e21dba04856cd00a64a43d4213d94d894cfe7ecac1b233b5d5c4a5b981df12dfc4aee3091d58c915dc7d8eb9a13f8d65f8a4ffc3c8a9f112e20f34c462c0ec9da1b214b07347d556190ff75fb8e9e8cc8b7adc4a8f27bb807e073ad79fd7eb9426f64219298a8fa8963f59a3f201f6452e505fb3ce6c92ffeeae047b137dbdd0989a4cbfab7f937ed2afc888daf33e30cfe90d2b086fb6bb22d00e43d200a5885cccbad8c2b92071652af95edb94e13c9a410e0a556bd148323178694f95c3829c195edabd6430b192836d9e928c9da5c85689bec94d2ee3137e4dea239bdcf80a8f74c1646e7e535625da1c8773d338a7a7663ff1fcd95aaf265592dc4055294a3184715d9a71658e541bfc6d54abb23d2d72ca4e161a9e99d3e05eb8b2a1a1edcfbd102a6938e74d82776d3e4e97e94c53a5c462e0109a06a48feccd3382fb04e5caad995a413b2715f705c647a1785e9eaea3a66b9bca98fb84475c62d8eb30dbc7e001cf6d0144ee302310d9fb2f549118d405760bfeb13a5f87d488e2638329cdae2f14816ca0b915d1f4c1731bcd08b5188c0a19a0c04ca2fa89a3879b451efeec773f8c117bbce17b7642e02a8777822b5b746167071572836bd3b8f9d5473cbbe4d2f4393a9364a44d50e345b29aee29438f06589e68f524b3f74aeb69f35595ff29c6380566a548278d786f05b467d4a5e92e30db38347c544112c79864f4aeb496db7ef900a774f9491d8f0864b5f01d300cb8d980352bfe882d34a55ca786ff20b6ccc65df19164d485f702e5125c3c1d24fdbe86c10a9db05771a502d18093180431e7b7bd219a53d55ff9bfa8b481d699bb18e6ef3b7e9902af630060ff9bf594a807cfb962261d221f0be521273401a00cd84f1402c74d99eba6839399843ddc7cd28da9da0e8c46ed13cb26ed094b439df2a585998862f2b387a0ba21707a101ba6984c5ab77b9c7fec9477c804a54244fffc976857716a924b322788a9770b16f9c37a78d085c2b2abec21e1041ff25eafa76f9ad3a285196af80d3969f0e54b6b3b2c00f8027a742b12d0fb62a478737ec0b3c45ca29e0210e2ba6d2739eba3b4f928b576dacf7522fc19ff24850195843dfcd77e71752afec2a9f2ef7d491954ab496d42b751bd5402172cde5fa26907c4354c468065631cdffdf402836c688951683929787bd93f7732024ddb8a0eded1c92e25ffdb379557b84b0d7c68b21ab84e6dfc0ba79a094bea648a69a7fdf929cc127430d20207bac399787d80223f417bef31e99e62a722eaa4106c76ba40ae9f48fb50ed5e0a562a23eae1b49bc3a2361ff03f8785699df9d2260bcd3925f938c94e9166a804a0796547d3490477330f5d12f0d09ec5d5f35500515bf7c280b9781a0b354bb640cfc57f2b933989de2887ce1ea6c357eab0c60d1981e788d6ef931af005582d7ce2b6f8ef59eb5092874d0a0b41365a511a1b91f675d768618fe3f683601e2cc71b4c31b5ff3f08488208e0a362c6091c984dbd7882754d9bd783bfdb2b74e6d404a3c6dc561abe3061f8340f0f080a3baa5871163b2a9dd5b14e87774e6892ad07d439d89d2b005ad0a4bcb98f7d7352e5f8e559923c767f261c427922c946965cfbb53518526f1fe933356199ce35ea79a6d11d69ee8820edba2d00171dad06f8dec0cb0b791f3ab0b924950f7d8ae24e0c8540cb4d4dcd4c4c546f36f6ee19f43b2670b0459fc32a8075279b70694242407d310d001e0b720502a5eefe80f8ffcb115f2b2d06608c39dbae7e001b3afadc276b9db128a406d1ee09d32b2d7d8bced8595f07de9aa16df0e1eec955ec3b711c19ac75460de1db0c82961ac908681d4875807dd4964c47f7b33f436a2c609c27df8bd217565f99ad253d6804b5181ca8e0ca2ec51ba0e556a3cd6c4757d6c9e8374db7b19182d592ea4ed87881c86517ff2f01d594a27c025f314f7fcd23e88f47ea9535df94ff528ef83438c51a348a83d14fa75fa396a58a47ab4fe7ff932c66d6c541cbb02e033bc9fc849ca4c056a145b2d578dd4f904a32d13fba712d70a778ae377316140697adcd138a1dce669602f473c00e64382a2addf834dd09702c555c75966aa737b62fc2135892ef9b8639376ebdac3e0255d4b1768a5bc2847b95d04a4f4dd3d04a68c7980c5bef8637ec8e88fcfcdf5493d8f617c62a1ae63cd21e205bedce53142d098da7b7c4a76ff1e5baf6f0843b05e9d8bbefa2d6b258fe79656e8828b3033c0e66f782b3e7616d0ad313f3e7a5ee6dc70449cb1995d80498bb30f736c55321f2adf4dbc48feffda3a29d7c285141c531b07c004bffa39a5d52445dd962a3635ab48eb5975663000d0b9340d14744b9b2ec31d23624b1b65541ae2074638aaa6ee5fd0aefb9e88c045041bc481067a6698bdca6b45f60d18beb06bc64ea4b7537ca1ef52393af8a950a2586665a689aef64955d6104368ff6d4a7e179b46c35ddc52a2bdb1ca05183fd7ad872ed1db7e702256f5a307e51737adef2061a83a943e0fa8d9447397bd596f609d2606b08e2b2a9af9d1475aa0f84e6966f56aa6a3729076c3ace435f0c33ebf24c400bcd202810d83885bba6be2f3e63c1a5d20ff10cb1467a32d6eb24b07abffcafe0d145c21e6108cacf3614f913a86722e1853a6a213f83d1ce88ee2d7b0a1fd06ab656c834d729d197d737e820f991f3044b5c425a979f7842f19c6b621525cbdb7f6232617d57555ca6c7adbd8669e660177dc90abb3422b4f3a4f78437e089b4852c492f29123a4c6b54da0b694afbeb7514a4ab4f55807f684a7047706e9664aa770de7fe699fc105a264c51f77c6c3a36c28f362b55d6bb2e25511a7bf482119d5ea2275fc2d1c863de27fa09038e99e9a900f075844c8c3a3d991ddf98d5670e7811f8355bfbc52a3c5244f9982b9b1544385f1c592e9cc8dcff1c6f34322f6b37f4e9d367157f2683f5eb4fbecf90b9cce1cfaf666b48d678e36c7cf851119acec008c37468a315643825119fe0473507c8c92d9aaefb92b6fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h6e2754d77ef1c0c2394e8b9c30e29b36e8e4c6171f66e7be88102cca1ab01c6ad91f59aad26db058cb14d6db905ab6f0f9cfcac2e7676e9e8afa84ce20f26700ac476183e2a51c76e8780c2cad4ba28ff5f50266b13a007bf783819b7ae20284d5fbddf893bcb83e85cc55feffee18391efdea7a40a2f95a36f7db033572382f5ffcd5d8188c1c573c4aca09f7f40914b377a92ae35a408d0084099229d52efb05febd3e8ef718b0c97653f01649463750e29710e66f99a5c32046bf49bffe169e25c987d83d82721735f87852fb5a5e0b016d758605eab7cfe0833269d6c958d86ff036d24ff15b5387686577e74cefd2629304c401493c39bdd3f8f0ca604a388dc4a07a8bb3b2a555a45f63e37ab238cc7dd68457d5e501986d0876dcd6c7677f4eefdb77416953128cbe8101adeb39cadf9e1c8d4e6c4d8d8a089fa78ea302f58307a23fee1644acc2cd1f452660abb5c55116af874f5c3b298e2b80b2abbb90b7c20e863db5c5a9fdc1bddf9651bf23a352e46821e98bcb6c8f2ad793ab5a7f5c5433503665dcac2fbec972cb18345451e88349843ca8df73be6b455cf97e655251790bea7962a7ac342da7ced8832d9ff267bafbe9641824b6c71d506aeafbd8afc7a4a6fc0303472896510dc345f979203d5fe6891e6675709aee9373cdd54f1a626f27ea9b21d0928e3251edce2602948f1053b12130cfd52fbc8b0cbbceabfb19e873dc55e1a441916b04e4104ed3d7b43d804490b3b020769bf03497f9fc0a6a1650e0d652121ae00c7d16543001a677faa5db9a5d9ba48b7569c5f76056c02f4715d5f1a9d3f32e3028fdebce88d10804a9985696ed80686bf4eb90ca6187720ee5c008c882577701477e3475c240cf15d632d550efdce1bfbe89cfc94acdf3da986040f35d25690e0161cf997c265f8be4ed1372379e32bbd1f6a13a69035c8933ed9823ffe4ef3e24a164a2a1d28328101bbe78cc22bdb36b7a8f098eba8eea781717025e43498ee423c53241b466d602d9bc5c1a2a2dbbfaf120c1a9bbc534c6e6ba5401b22574d3d26b974939a44081ce40dffdf4426a49c9f7e14f0a9fc484cd1a3cf3b9f14545e83dfd06f755cd8187a16d4db4b7bec7426114d68acda369aa6bde48619130054aeb764a7cd1f2c790ac83f47c59d3fb3ae93e451483c37161a3ce687ba04b970199f0118c69b4be9e92399c0e31c27c19bb41b9017add6d515a976f7f17136307ea78f8e9b56e0cd6cbe4f86d961dfaa5f8a2aee6bc32c67654dd90d1c1d901770062ca6acc927e94166184fe84e9c188f3bf3d9cf3223e5b32ac17382c9866b22d3aee59bb314ef5566693c6f224796f2fa1eae37b93fffe9fa2a83a30d5af8460f8f5fd8c650b8f478e961458102526cb84ff1818139d4f4aed68b47621d863501fdc1da22a73f7f08bbdab769be52ee696f715934f3638cde7f09516561e76f5b8d669452b63e5773f03cba47b2bf5165200f4cc730204e201884ab0a7efe8e70e1c6db28dc87a82bb7b5827acf935a381298c3675d71c3d099879a3b6714d2a48c317264367adb59cc94509630e4a75e77f2007e768bbf74a00d4773a15a9783d3d73df47ca20abc9f35b4fe6620cc3b2c8f055fe08b7e1a18e5a4bcf813652a0db1c089ab1d4ce67b1c3f4a07663789d01c391c7e9512c63b0ea97c3cdacfc39064b10128497fd4d56481e5f68f7f8f47affe9434aaf9aa2c6584990ae42976d77b230b2f3ea22f5e4d94190e977e89370926ec8ba5b712f4ac17aabc5322b81308e0f8161d4f7d736cd5d2cf34ad093d105fff9939870529fc7f694ec75624f07cbd0f0889d81820eca94fc841baa784d8285409e939e3db3debfa1d67b1b5d05a27e45fcdf349cdfe55fbc0a0dfde68fdabb4180028429aeee6b2d73b3082c7b713f401bb5dfa6b034e3bf53521cd3e2c0bf221e9dea2afd96ad58cf02caedc721765e776779ffc851e2e27254568b7d8c7b5037a8efe324a2f9c41ef2de9c2bd2f801f816ba91ad2e390e52d1832e7d4a69e70a041762c59fd1fd33ec502cf05c77c08b8252d75506113325378a150ac892eacc4eeefad562b70d6aa3dba704f168b65de2984292fcb1bcaf5e7f39b0737817a208c1663f7716ed407bf31d712ed5141f3257edbba2808d711ca61b2b1995345d8c6d341614b9966602cd72f82bbd63c6093d7e1ae8bdb782afb9cd741714f5e66b26c642f339d4d5bff5f0cbc081e8eceb0c9355d6bd27226bee2ea65c59c16ebd80920ab49ed90ad1c484ac91dadce0b62d37a556c01aca70ccbaf25bbb4b171efb9fcf34ce4b7d885d5ed9318dcabdcfd81a5f13f64df54b8ff34440b4917b37c2ab2fc17aec61ad01059200134fe8a40c5fa1f93b33a5ffbb10190895a94d4eec00214473912256252f2b6b03ee87b554ff33ff0407b2d2cd905d166e4e901218fb9c65dd2d626a98da683914d1b9fb8da0f4d2a12e4cc253e75f1ff157488723656bedce713f3074ff0743b7d7de91e932bf9c789b63d14f16bc1099f9521b4e51cdfb584d3df5f7d40185d7d67dfcec7c903a2fcaaa7756b4c8c7ed8be956e7c42b2438c7b224631a941cdf7fe2570203f17f8466c329e140be29e52298ee924ee9289423de24fbceec6f8188c58ec5aede30cafce6ac84993eaaf91664766f9b23f016db031e75751794bd3564996dc7ca7517da779419c888aa79d2df3fd302ea369e335acdce4935df7447e7cff5c32bd71ff6d2d3accd84f84b49c3f29cd2846240efc99beae4b3c65523125a90dc49c297c5b645a2cbc385bc0f6e82a470971425b88bf35beabd4898e63f112221714dc3b325f1bc33fbf90df27a353d82a8bb363aa1bff6fb6a79aa9a1bc7470a1d29fe1bbcae4cf40afdb81882ef674f8f3d7147dce9f69f9af2cd198417f89da02d00edc12cd2c587a4a26e1ea03303621d3deb13a38ccceea787d25a2ed37308b5cb53731f77ae3be99627e3436a98b830b77bd36e08fb0a953b600ef1e849b01a214b0a2efcc4255df2df8a02a8f22e023527b66ed840d4ccf4e5e478f79cff3c2c70cc1740c1ac397625835ce679b2be30725f172f9edc6fcd19346f57bb8f0f94e6bc7d6059e1b7e7a6f68d348023e2ed282d1f8e8703e4315582937b715cfbaad70afddd8aa6415c49e6fbfb8c4265d8946ca3d16f8df7fb0fa0dd2ab6fc455c43ce11e98b03caaa57333bd4c914fb69594480d8af88ee585937584ed444a730f6ab7fb3c19f1d986ef917c37ce045bfc26fb1f9b09401b505e6797851f562d2565097df8607424adac1bc0a1405041891739cabdb52ddc2aed70fd22b99f09829af7fdf09321cdb2388fa174624b6a2e764ee7c3311c4f5899c483f5cc1fef9403232af5eec5c52b36e37368fa5e926f3103fd3f4c1dab12d3368d44da144d0d83eb355012f494a9404fdc514ba84bef15c0a5e815d0d8998f3664a0c0b43f596d6dbae40dcaf46491fb2ca6778692cc2d4e04bd7459b9999ed39d9e861e42cf14f10ee997aad028008cc74f93afd2b12ab7dd03485b7984b84bb9c5f972f2635976cb9795ee52ecda07cb2175f654f65a2778de507e1cad8d662b72865845e9766e32540e07b31c9f229df27628e90b5e64c91112fdcf5f3208e0c4f1fe7234cbb88bdcccde5071fcdb558c6f2b42454ea8f011e8d4283121a7de781cf5f4df2036627cb189509e7dd900e9d5cefa2b65d8617ba449881f71938231a03dc9fc6587065d3642176b36744d676d63bbbee3b172cef1b1e809d8bcb724ea817a1ba8ea01dc204013e46c3138e4ad7052f818cbda23b91d1c9e46afb549362725ee1c1ad1cd17a5c5351e7bf93646db4cd66159826804a72b2ae1487aca9b53ff961ad46993643842a41ecf25f39c76febf6e1207da5d9c0ac81213d630c7b46d1f64137cebfbc5eb02b174a1cfd7ede1403f099e58d48ebab0a0af94a443b64e5a2de5030a1d5c840ff0bed55a5df42e2803e7fd7dc944010c8b0f3341cf217627827e266f3085b110c21efaf6f5566cc579a3017812c442bdb55c004311e040749ac65af716a1dbc7a34e44afb57e35f4ed67210c61247fd55b940b09a12c77e73acabfb60f9d60212fca3c8b0ef4bbb3a53eae80f5c580ef14778e6c12ca3c921cd9ad0fb03e0c95a9c4cf185e97561e91faf48b5436a8cd41cccb7e818523b72e6b9d43ca8ca00a5937d09718143ebdfdf87e5b8d2d83a25b2c21b3700bfad0808478f5aa370803a65d1d795430c77743a62b6ae65ad362df469eeb15215779f42a8f35352b03b09953a0df0a83013155df5e48371f0af0fa0dfae3ba006ab4569b367a85953b0ea4d85d43d03b4c5a1a35d43d95badfebdfc6d74a58597e9cecb99d81df5d2103c2138d498dc7afcb761e976c2d8f24e92fda4176e4a37738226d17b03c3907b491e420e740fb74b2fd4cf2f33b21a3a0fbe2a14a1339d800f168c0a7155fbe24eebe824460229ccd4e317f1dc07e9b2f3eb5e3c645015407f8b21fab24804724ce684170b0d67c7e8cd742c452623271d02b72214401dd15699640e9f5a2eb853d7208df3dec92d025e5b7131e009104ac020222ddf69d90ecd8bcc99cbcf6fc18b618d5025e92a73746bf260217a484242862191803772b705d68acd52648069532b4788dc6efee1cb5c6d8fba5f90f5b715d25328ad64bf5449c82897b73c2e5717fecda4730f305cbf11534bff658bd3475892e91f9e1a8bee59dd3c50b5df820bbe161931dae3c93970e9580bbd9f2304fe04f41b52f34aec0887a235806ab356e80b2ecb5245d36cc303cbf5ccc6c79538e90975ab205117cce9e6a8178a61c703edd3ac3d7ea211b587a16060c74dd0ac19e23d0831f6d0d688d02f9bddab1924fc7a6aaedfeb858635362b83355bc460a15d53dbc812430d9fa2637e1e27b0a0e109749c104866ef51b11f70573c824bff4710cceb2559cdeddb24e63279696c3e41060c83b5e06b99c0affa5ee34d7aef64c17e880531bf6adf86b47d9aaf4dc37f18590a03656b618c9686eae654ecbe7402874434a12f2b39bf0beeee4fe479fb462caf2a9ae88d87328357f1034c2f0d990444965358dc6abc7c36e4c3208fea2822ca7b88ecd342569e868d2191a971dd942d97505bd819dfb0f2cdfac36e60452c5c35d0906c46d5ab10c015e5c783cf4670ae67db16872cd4d8fef471426629b15d345843dd4cd5f28651100b2e08b5057d07bb5fe7d442639ee346f33f19809a2b74325f9776309c63a0a98e3d70548799d3c4ad377f34a44f7d8560ece9bd7aa06671c2ae56c29b7d64841f4e7810db1e130152076a4e30cdff46ab296e3a461b053f60569294a19042eba108b61cd4ab7d2aed6ee544e9121ceb5d36b3b7a15fb43e923229d71d44ea074240b2588605544ac3e107960102d9357473b23ce62182ff206e1a811582a91446fcf557568022f72ce8e709e691a781587b3292073a7cffd0447cb9c5976232fa7f7873b42c96d54d018462002ca95d0a5c87ef4c6610f7d04c8b6a39314c5fbb0168f5dcc2dec3074a837e249946720fa65ca9107cfc5b22df87efa9eab7eaabf632c57039ad29568be15b700712fe5d3fccddfd435a36876602c35b3579234a2fdcef0abf54d351d8aca393edeef21683b58e40d2f66db493144ac713c0c6fd2d7036e9cf123222a16763136606f95ea697665d341fdfb8fb1b704c1b54ba6ec7e7d5c5ece9002c3d5bfe11d4fe5c422d5823eb33cf6d12a9859e403c3733995c129533e57db7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h432da388204a1e16907b3dc9f43397db20a9ebb7727f5c654a5cc8b0ce2d875be54395a24c09083b996c94e1caaf82659c89d993187647469685459d24199307cac690ca8a7c08c26403266f107c759aeda9fad0139d434d9a5a8663911566d5856389caf85fbf0947283c30b042fdf6b37a29b8edab288ad5ab623330ec12a4584e78828f0fb91e49bb9e61df8203e8cc6855e95080874d234ddd33f6f61ecc0c4d95bcdf8775968b33eea95da5fb3f132866e65150e44e94f9734b93d30fe4988d07707f71b168d9c181feae395df9f806d6bd7dff5df00730f1fece65579f1aa873e17f79001e9a51d6d22b355709c20219bee491eaeac10f0315fc7032605d2148de67444bef2cbfe7901100b7b5ae38ada62d5e06c2b51d6e98cbe3508bcb73296d4cdb42e9889fb1002df8107635937951bfcf401f0055bbfc76e2846d2be9df6ea5dba1ffd051fc0e88d96b7bde2d90739df6cfc47ffb1536dcc6779f941b5f1bfc262710e6df2ca691686e4d10ca2b9de9e66aee448f05abda2f82fdb0c1bb2965b753d40e29e7aa592140ad762a649f7493aadbc79896a89d81b2a7d7d8dcccdb554d7473b5d908ef4b517656d93f9bd29072883e390d41335672a3a00758538efa1ef68aeeab3fffbe9460451988bacad4bacc03574851876d77a7859bbab6fe9aa31e510873a8cfb247e63e1a4bf80a4c206b1abd30e1f5a440fa1238f1512c01fdb76f9ffb547b5ad40a51a9cedc2d0e84240f787b55117ad07f1b50033ce0f29a1b9b118af0cf669971707f017163ea8ea7b253dbaa908fc3fbe7264854b38a18a942880453caa8a0d6763c7bfb4058cba41fa583db919940b15540713d970f6214daaa9b74124752bbeaab99c95b39975f07fa4559270e5d900944681a70c04bb780129fdf374b8c665158b14fd32018a00b3b445c8f94a1c664fc3984bb17eb6faf690e55b6c452030b27c29f0efa72cb6edd9ded6c794a205ddcebdee87e0403bfb81810101f725d1fc3cb752fc1fb6cef36b4ea9da0ad78decbefd1fd0f86b530dd7cd286dec4c207e94e12834cdb032c4b41eca41eda31ea87f73d9c986b0d984431787a217e1a20ab8b47b6f821afbd49983deaa512ba706f9907a41a420496c6b05cd1af81d40ef930fa6a230ac2020cb3cc54e29311bf6dbc7ee31d027e74105cdc1fdb15fe4250e5630282a0012c4019623c310bcf7cfcdb1845a1b76681e5063a0d04d3e9e8f69ed97c0086b6d45e46b60684b933e5df040c85381536fee9325724f0fb91b6fba363bb52e0000bcd43d58630763fd134ec5a0767ddf56e5d906bb9ba6665a3eee471af81f0167243ce516469887dfac022114ed65a82434aaefb48cabffe7cd76b449f334370d3a8b71ebc6ba1deefcedee5f3eb077f9f57fc5c1d46dc5537c9d1d27fd4115d51ba6d219d789e3c07c95143cedc28d79faab1a60300477c35d86b922a93c9ef32132aeb0bb7c89f6265131551dafec35ea14f1cf623fcea19cd7337b5bcefa4e7a44aac23289646b18a9f33758b124a3c6a43ba96f2e003ecf5e7a5a08df32205ead26700c1bf98951ab00122cbaf18d6c85b8bd8b1c07e1e4bc66115b016a33f99c544eb95a9e7e3db7f2b5a21c04bc2c4191467e1c6eb8f08616bd7ce44d58a293fda0ee21effe379c3884115214a2b15df38b20943f5074f9d5aac36ada33223089d9b74340f231351cd155eb144d7d90467a452209864495507c79de1c3ba27e12761f63c1aba1d0084fbca9b73e814cb8b18b6826f6d0c01e5620603e4fc9861e3134b1ad25e4c96c27d0b10f6411974b9344e905aa070e8ba5ea3cdcfbcce17c595e1adbce4ecc5953a516ffcfcf595770b3ba5d35745a23bc610e172ae673ab73d5ac34a8fd8819afcd039158a0eb3d6d93cb46237415a115a9fa3da2b58cc85c6f86818f54262bee046a85cb5f0c07f515283a42e68eb341a793e885aeee943372942ee0657f9fc87bf5c78ef17a8a31cd1588b0187eb1711d940fe568d47889cd7289a52236e52437c58d3ad9d945acff14fd4cbaf222fd6ab89388094de3f1fd6fe974a099ac883dfc1b41f58a293ae1ba0891522759230ab7c35fd02f02cb53a7b9133a894ca8423d29616e1529b41571c0000855383c793b41958ecef7fa24a43763f7764a63c7904cab505367a14bcbb098cf6693f584393f438c01be7ae0f5a260d4efded0576dc296777b1e36eb29358d5f665b699f053116382139905b7e035713a3b4798c42c661198ec09b545c9972b45315d76735ff637669b0523f5b38080d8351b29ae5c2a98fb3cb89fd98d69d0df45a104715ccc960aa8420aabadbe6a473b26407455c28f62a6ff50692b6fc8bf28b7f3f2fec7d8c1a3fc754e55ead41c530655fe105586123ae918b4013d25aae27f9c3d30855e7f18de0058cea4f45c32368cd1b69f356514584c6696fc16e5f75e3374e09cf51151f76e18212709589bcfada84e896fa8e580f4248cd1ddd70a73ad488361821985e93df095f31ce3ab2407448ae02bebea2bbb2f8047f491dc34d4720ec0fb446db5e939d77aedaf36a0ec4b6418e0a68ef1064c3a2daafdfddcfa9fb1401fe02f22100a031e8a19c7fd1f18ed061789c1157ea6e1a4642a9c025bd606188dee597666c60ffc4c10838ff1e08234adf06c2134d78356852bcec0af28ecf678545c2df1aa753a4f2420d499748179573db9d5fe6aab1031be24fe25707326ca7d679a932b74b4826b2e8184be320d9df5307ce5529668166cf204b65bde64ef3daadff83484631b2c30f1a6a498a61489e147b3d627d99c13f2184136a03941890b1f3c2917e48a9c2dd29ddf8194ae3085cf0ba7ed4f7d57ecdb9b7d6bdfca99253f87b0c515cf8c543e7f458c4a4d547cf9f03b9c1f6805b30cfc466b952dcf9ffe28c13020bf3d40822b41fa998bf31c0715c72b835ee392ea112669166577f7d8a449a5aab02a349a5f3da2ac7a68acb26fd0fb174e3b8a9fc4c943fb9b311b0bc6c893a749743ca45f1c6377174e73fb1d8055288680be87f94e0f0bcf71d20750106aa53f1df1669cfb59c0f45a330e3bbdcc7604a78f7f05520a2257955ac923dd8fa874c2cf7a7c4b94f135b04c4a1feadf878e5ccf9f6e6ed1e263b4521bd3053dd206d291d9b7b62b671bb8c6c2a8dcf6ea4607f5d889342b12b0579c3b360e7170ec66865358fec3836b8c821e4df143eb23721c2e4d50d48b9cb95999cc4630f3554691948f9c15cac7614dc11e0e223333a2fc2008ae3afe1cbe79fb8e7ba5aa4a56f21683c75cb6b4b0d629aca227b2f4e87e0d9079bd028dfa24ecc97496fb53a2f557163e321a2161108acf7fe561426470d2498b7719ea63308a7d827cb8c3ff8146ae8aaf9be427afc680553b2b6fa81e61b26e4445492af201e658a09f35a9a2b213f312c4a855536a60a700c001eccbfab7be7c6148148e17331221b6ed621a8a2fdcc523a76edb051edd1f4e1642a77dee85450e77ee88d8ab03208eb0bf449d2c7245097d5db9b5fdbe1e20f9ac0523d8bcb139d42f00c1bafcfd5e4bfeed0b6eb681b43cc1233d9c0149bf9e6666ecfcff853a67291a898d696ca67ab9e9e5c145b7e459ee608a26ceedceb37cb2b444d43447e0fef01e66286c272e368b705e7d60a9474d6981e061409194f3110c5f91550477e83c4ffcd7a77c04b0234deaa387b283578489a44b7191f6ec0eeb9c9a888ce3f9ede6c854d48fddc589041514b2988a72eca914655cd8288d24271e386c349e5658f57b605c923974c2057922ccd755dd35a3466dcca08674259f30ae3b9a7173d0b0e748c5f3375461a0b67fe30c3e1f434b60f437d77543a6769af9fc1559d00647f5a65e70cf0a01ec499c53c733401389143bd8d002a9aead38703bbc3c87ea3d812568d6143fcda3f23d7d0fc899f68e538fd9bf25ab6632e44cdc6665f06a66802f803bc33d21f7b4d627c86a3b744877790161a58d1e96477ce55ed132151fe3e11fc7096d5f36a6a645c020119032374b261eb6574c986be377122256c3152a4e4e33634197ee5605c91c8bcf0ec67477af3eeb7e7dfcd372f98352b70125d7e769a4f75c0d52357bd7eadb764bc9b4e350db1002ef93656f99941df019a8883e5ee25e6da81b155a05254b5372fe253ab06842fbac90d118afc71d32e9a12cc633f09665ac2749ea5503695c9c21143849ba2500cef03c98c1943083a04bb8e31a79e188426139809e846b7d583166824900cb0483a8ad1d2a5a5245b93b54622619c8ee57eec081d07f64e2025c7e9cbcac05e7cdc53767bbb1b262b0a240be14994f63e86886db61f8f95094f5b34505158ea2360d4183342bd4d0a2dc2352e0a4f790e40e5e80e4e6b16d1806170197ce8ba31dbd19906b03a34ede8261695901c24f698aee4cf4ed4726b91ca1005a2be1cf4f5ecc7e8541b6dd831f753386d2aea083f817c725269fd1e6f03ce924b4676faeb1891cd0cfa6738a3e051bb98b4d7288fd605500af862601170e5414e4d560ac291263d4d5fab58d00da082bfb55468603014b88aa21af8b93501e4e6d2ec55c7f194dda83825c5db5e196d7253c7ff2eb602be02fd6eb850668db5d1f6f0fbcf00678c7076d1007b8d8eb3aa3ca04c2bcf565da97e08fb7df632511254664c44ffa8e936bd0072251d7a53afb4618b8a88c9602854899b7c2d797f949a1c86283b1d3b1c4b868915b2a5a9ae980567d16d00f58e3209ca0a951f6832ab3acedbfdaa2349b82fb30aaa6637df7d25bf6460465bf689b852c739f9fea26c1d24e595da360238834684984faacfe940d9b8ec20ea334665489b6849b248bff2f28c28fa1b17815635d6b4cf17e6434944dc9d31da94f3c3a821eb5e9b2117456256898b8e5df0e5ceab6f37578243cbc4f22d3cd5f8adcde5edd9d341ebef5f31405e8e00efda1d27a84918d1794cc74257e727495e2af7637af3f8cf8d77f12b6f63845ce985b135fa3615be1b7bc263fdc7cc70b3c2d7ed93ac7a985bee722c2390b1fcc537019e3467cb2f5c5e521bda1a08d010a721600122eaff147c737e925cce741574d2c5b9d266dfe4a816ca8137c6183f8a5bfa178b98c6ef68be9bb4cd9743dae311e3c08cf5e57dd1f6232c5815718857ff571d2d0d99f5725cbbdb78e39603dc3f9ac9513ce6ca8e1f2ead50205d3c543488225b23bde7eab232cb445f86281af079035efa9a23ebefc77bb263cd73fa6cbe937c2c08fa3826b8420de595baab6be42319d6777dc27a6de24c14000efa026faba95ce6efc7b1315cd2268f36d5dc94cd000192c8594eca7ec0d99b6e634d02bed2ac2fc42135ebd0cdebbc0052ce17afc731d65f3c90f4802cd23233df3e58cae9c7923ec2a4a90a4c8f6bd756967512a56ecd9d95283a850316b364ea024cf0f20bc6c4b2997ca187a92527a97277c7f96eec2492304592d3d8be148fdd24d6840319e152e3e423a0665c33338dbb25f27dc88d72846a83d4b917603c62098df1e9e9fa2fb029e44ac4b7cd906a5427cc681fe330451cf719f7cca1c78df30d197912fa1558a06382a7cf113321f7f66500f3af8a07b220e8f4efabcc8caca9ae2b57f3b231c4a98cb771664072b916b4b526dfba6f35417da415379b281ee9c6fc2c6b50894f76f3de0ca1280577db14e8266841e5c352e00b6a447bb305a25711bc134e8654075ffab0aec70aa824e6d3677511680e3920161bcfb013e68606c9dcc3e6254782b35e8efa29a8e1356bca90234;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h9d4d9dd3f0b401c0b71ff3739d0102cd00e838a93ffade86289fb6d7fe0948524301a894e9c7fc21a21e66d779667baa6376c3382c3f909df39fa7d16593052c65836c19ace0edcecad7f852bdc972acca03301263b7aa41608c0587e656f438e07c3bf851fc92c46fdb61b7a7ae066b12ff162ce8efc11c043020000abf7b5aff5f72f5f3a272baee40e5e22e4faf0ca05cc1b5a914726cc61d32d265fd322b50256936108b4ec58256fcb50acc2c5cdfd5dd18201b9ca1ef6a3fa727a6547c3167299e7c85cdf1afd97b8955b2e44852c1f0244c5b2dc203e8d277889d9e0d2697cf9930a2a0e26c15f22b590097081ebe9fa2c818cd0a8f73854eb66aa52e2307aedb613ff8598f7be42373347cb273d0f758923b0f2e38f3392c53206bb852e71652a0773f24544efc640a3d71f50912a27c40ae06f2850ab90b296d49d187c9160465e43394ce10ed74696df812c92821ae6abac1b7905fb77818528cdebbe566709ae6105583b9da50f070e3842b172185f028589fdd17ba7a5f1050bac58e9baed216efc6920a2074f6f94066d6a7cd65602a8ba315d5066023035163031895b8b775f34feefd39b42d9baa1db1a8d068886adc9bb0f97926ef902e33173b9107f85a00b5b4d29c0d67a6cd7e1f93d95e90b60c46aa9642565009a8442466931b2580af77596cfd6aad9dd5b72a33bbd1fc4b01e57bf4e8bbabdcb0a54574bf237924ed337c2f224e72f021dc88283bd48ad9982400485013ba461f948b009b50d8b1796240bbfa9f9998046dfe761a73b029cfeec3b304989c1fbb07986c8a332e54d999a3d96d2c66f8732e6d9b3d8f975dc7fcbb892f2f257ee07d03f9324e42802919f0001388e5b702bc2a8957f0c9e515d8773103af4f726228361024ef3e84160932d2033b7c426a22a5f7ea0afbd317cd85886183664a97bf736e6c2031b79e7c32f0df7bd4fc2aeee5263c299f39c93e08821fcce7c6c6e545662c1b6e8aa264fee4c47eb57b9132344123a979041bc29d4b3fd974c680a16821a2c8bc9f91be34b5cbe3b61ee4fb3204acb9761b44e4f682e39ab6329b6e3090b1eb4f1c1359d49fdb36fcf361b930ffc0ea628d32d011fd58f5333795a642713cc7110a811a2af424ff12351bbdab88be3ffa2a06d44fb733ab00937d853792663885b5257ea04d782a4293cf594ef5727406690c128a7642f3a5c74adc00038d6d0a7f0b132388cf9d2707fbb4b05f14bf6ca6767742a395f1a62be986fbec992cfe4ad01a51413280cebbc953f3211d8672bb2f1e8cdc5c49ce88e047cbc0dc69340da44b5350ffd8c0b32280e2d72fa4f56e49f757401dfa1fdcc0e3bfa4c78ba1344814a7731b2f3f7bf09d4e3ac2361b77fa3813e5383c6880b3e11659e1a460d6055b3b52803b5eaaf3977de814f46a3b5b9030d7e2e2dae28a8b53a02ec6b56f1371437a143c1785ff3be540b6098f6d413eacabeea8ff9b1a32c9b5ee4cac728ea2564bb0ab05b6131187998554b9bd77935d688fc620635197176512b30bd8bfcee5fbe413cbd8a4ae8b5bd2e29bcff1d5a51ee1d28b99d006142ea99e6dfe8a5de69ca56fd2992c98ec5d6c19a0a68e1e5a05310ea4511df0eeec1b19da3759c605b51a31681b12e6e3152f25b6d84bc6d2098f79806f39e5d221e21ca4b991e5cdf6fecfad97df26c37ea81838b8e9bc9ae1c046cb2fd3ebf69de68435251eacc02f3f27df7cfe9963f1623f29748cbb857bf4d9456433092dce2e2629585b58478692525a5775bc4f8fac42a178bee163f61ebb0e95c1269f751b982f2505251f815765f5341a2f681ede7abc4e7733c1adfbea622784e65d013d49041e808da78ec10b6bb7ea64ce6b1d81488a066f324338163cab0f71cecd32b0232436422622dd1b7c3461a36d733b6bdfc55544422d6aa5673efa92781281dcfee0dda5cc1b54d5ed3c4e2f6cbb2851480fc8a057108ef554d730730a9a7aa1a552ccb1f3b2e5890cc4e8f41f358ce5b22165384417cc725cf1af2d7d0263c8f7cf05bac9c5c297a7333d6e76c5518c56959bc19dec2cfbc2ffd771bd508bcd3ed5d5db405e6f22140a87b7a25ce43d9b1ea1e2e0c6b8781d3d9223ffefd4730696f0b92b6e30262e2701f2e9d40b9c6c81bb82eead120dcc1f0b86c01350829be0d470ce12f8fe9fe423004b7e6415cd537badaef692ca5308b4b79485c1bfb64c441eb961f450d8a486ad01971086ccbab287165854929c85061e82f9705bf468ef5c3ff28336f7c00382eecb4fe8bb073bb2877a7b3ab39851bab8ed9450f46c72c95851347a8630a6a71eaa3f1033ef54c9c50c1a0575ae7323f0a2041101b0da913082c95ad35366e52aa29a7837da6944b99eb95fbf5860e5a2d72e958c7a788c4d102a091d8e5d99fc90a13b6c04607745a9962d3d9670e69c57c75cf1ad55664c4b655e2d72f3e14fa6e9294877662150003d4881595a8ee2e1ae0d2cc62853258ace25813e900d794cde0ccb51c26cf268d3bfa844a2258ac5e8a23b043acbe8d8c45b7efff0fa9a5d41c73bb609450f325d21d2344f4c813407942a577982a6211f05da0db0e98695ba3aca9af0a805bac7221c021eb438a017b41e6e964d9e07ca6fcb080702cb393adab2cccd740dab57a7a1e5c0fbbb8d407d09f78de229eb172874dd0e9c797e26251c9ac0feedeeb857b98d90c12b885cbfc098fe07f481b43badec679e8b42351d95f7fec9cd4c7376416e017aa337d8e7df685fad39caa108ca754e27805cfe00dad184590daf554241d05d856631efd4a3625f30ccb2e14c3057d9d6083b23620c70593c529540f040edc4fec55a12c3a95faf63aa8ad61826fd3ea7ce99dcc9af60ac794024359c92e66add83c9a89b1f83793d86d31153ff5ad7d9a4e06577b14bcc5ecc9810ef1a7d0168c394d3d8772560ccfd6ae1667c622bb8277e4486c2eecb086edfdff1e88027e060a5f982e73963282e73bc23ff2f4a04225a9c6b62d76874cd2b6bba773a7babcbddaab3136f31f0f737810d7db310d52e14416d77574997b6f50474e26ea9d57b51781a624d19e29ae9eb17e53d3a5d397a22715291003ad7b54c902813097b202c5e34b6dba75350f0ad1ddb953f53ef54d11fd9499fd8d099d7e1762dc089ae1f11590b08123f9ecbcd477dfbca6d7453b80f3adc379a7802e61074366948440ad03c15e737d85ead88b9486d13a84bf1414016b7e3969a32dd5c2ecb0b588f48846ebf0d8845303a0d298ef5bcced241f063d491565d4887305ae111786dfade9f96d6fdb848b9a2655e931cfa8cfe356e0ab0562a6007583d2dc2c725f84518b93cc0e08f85246dfff6ec8c34287470a22b09b2d5f0da28a2cf4816266b60d636fe853db229edbf30bf207cd60c5683778eb69b141f3f9db894c212744b92d71daaccb3b41147f3a9adfec6d8b1973b753526a0f65062f6c6c06e432920550f4f9889b05444185d9f71231c24105996b6a03f365360816071dae18722881ffc1d3823dab16c31cfa9079944e1ae5c376adc418be0808dfbc247c9199f376c461b807a3bf0e4d443d4b1653732bc7ef16b4fd1b929b0802a46fd1a484bf57cfe7ba3b8c1232793511ef1a3f5adda1686321c411db8c03deda86db87058bb384ac66b5699db8a6c614a37d3e8aaa9394305c37ae80277ebdb304aa97ade3c4cec793eda4a3faf4b6449e33799e70aeabc592d78d25b700fe5f623ed802667e83654351edfd40ffabfa1c8c84f3656622156129f72f745c9a7cb99637607f0096bc400a6e5fe8a730f3d3388b47e444d6bf6d87b55d19836c7cde7d9eceb6c427844847ebe181c00ad0e245cd044743ea31a7520a2a1893214a0467753baa1752300a472eb56a03b9c5a7d7beacb4d1c51cd7c95f802db4068d40cac2e0dc90849e76f5b9f093e57edbef3097698ec28ca08542bf4d63797d21e39e05f75773a6484c5d73df4f02d56ae484ea8c0431666d2121778030f7d839781a514de05c50fea582ad13024d6035cbd6ce78b3ea7ea485a6d402c6431f8588844af21f4e9bd5d00ad2923749a4193a3ea51b3c18f9093b721ee75d77da5b6ff571fcebb6cd1f326d20f391c8d6971a045ff30cdddde29602f18cf61b365ee511c5a53cbfff1f14689c46efb6cbf7f5dc3bc282144ff4d5943048c8f0ca5a582bd9393a08bc803b0520386b758bebceda803993606111ff6003967dad7b96312100dd7667ae7df8f2a0ff17a2b9a3a5aa9ba4162cf0ac664c432a99ce772ba885e417ff4396afbbc20b8900589467a475013b0c5597a6125d1a7f25d533363a6102440b2e5e1c5277501e3be8c26cc29f71a385ef4116ed045cfa15087bfdd5140122a137ee85f1a3fbe58a8c7e6e6966a9a8200fe6a12d47d59ad01fdefc0e6b2dee512ee25e4df7fa38017efbd6265438cd4e77ddcc42a65b42334cd755904be0b54fd83e4b40eed9af5baa53b86763bec9d456fc295c99c2871cc4db14dc349bb479ccd2c536044541f6e8d3b665e1ed5a2edd6fba26e85c6564221458d2cc27f475a8a4aee4652fdd1c6effca698abb6a59f659c00d167b25362dd4c48638bfd0703d4943caac61907c08bf0eb14f34dd91fef12b06236a1788b728a1d7c804aecd1045197081d53feaefcebfc550d038ffc3e392c219bba7ff9373c7394cff6972c2281a606b2778605bcc3f35a4d3fd77eb57ac137c5dbdcfcecf198697880cf7ec25293214b143eca318a66c2e3fca2d40fc8e77b274adb6748a5ec79cc3430298323e9787282265028d0318670f4a223b8c6ef628869b05a5adcd7748b6880bd747548a09e01149771a0363af66e01501b5f8fa468b6b247673fd528985f3f531fa61ef2bc88da5922cfd5afe5d07181308cb047af1b17f39ac63f8453068161397454750002216e00db3c869514048f79a0f36f8cec905647be533e4172b64b56f825f1b70dc16f2b3d04b050f2335ee39c35eb622332e3eafd85e3acc8129662e0c66b4120efe07bb647c64871039afd6dc0135021bae0ff3d43904e5edc579a934e0c1acfc1a877f07374b32f773a236ab1af37e1d4a96c6c5daff86b0081bf661ac26b24c59abd807fb76328401e6c537e3a184ee636a465c10ca156f39dd88e702bf97afbed86eadee8aba5fad4a441ea0b8d5354291caa293c5710823e79f967dbc6d4dcb7d687b73998ccccafdda2829b452e12687d32a9f3d75d800f81b736dc51ffe1b6da0ac47cdf77cf8213f3f82a4a557b4c1bf3abdc6931c406df7d8181f037e2ef95e3332affdf6abbcdf3221fc157eea90115578b83368d6328fb6fabd10d4466993f6262245d8513750e9a7d485b93cd63637b57a86135f4f8e4a838fbdcdeb2e1a537e68cd63f95ef7b166a1acbd6d601581c19f2cee701fdaf984bf8975fd8cf80e78fa69cf34313d62b7180edd9362fcc386d10d2b0f15134351cd3a2bcaa0efecdcc9600532bfc833d0d606b31e68699ebf60f1cdebd460441add9cc3958467e5b711c8910a13a1fcea5d78414603a054bcf516871cffc2d458469d1e452858dcb437ef3bec689307470e4b1e8d736b68c6a628bdd07fa454eb111c21f31e4a7875b8242720b1a18dc4999dfc8bb951da0be0d8c7355b439396ab65d088dbd1d5dd6404dbb4ceed6525de7877fd7fbd9ef56915aca4979f2ca082252e311ac927d3f6660eb6c25ba0f2a2f574e6b4e18f22100083a02db1e8f440bdc4d2f3cbbcfa34d7e0dca15243a0784cc099d93e884fe819677c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf8d7b757f9a7bfb7f8caceb134784f240203ecfd3e7410be391db4d837db3b418fabf9acc2296e49a0a5ff7bec4e64c4451db40b42fe3c98cb6b25796d1d933010651f0529e2ca6fbd2f113e771aae41077bd226c960d6060e20d8394ced98455fa1359946c8214ca2375f47bc9cd29adfbe56c14fbdb292af2230c6b40d82d69991c3a664fe8d7630813c4c62452c54ab0c602f325e8ad433d917a1bbcdcd160274b15b250e7bb4d6a6a429d674c455b68089fb587cef033542d6513965aa7404e02816537c431271490e87d217c49730c36679480c7dda39506fe546a4ebe7139ee66550883d834f77cbdd3b9097b316f76bb1217a489c2d61270d4d7953d4d3160ac960453385561b33a1dfcfbf7ab3073745441a1f2af1643a58a02ca125dd885150dbe527533c3ff5edda4e101210b31af01285803b512dbd25b2f206933d00d94cb1d1394b111ef02ad06779c2331f6c1a052b8b9707673785da166d40af957c1c3823cfae2aec12b03bc7d4aa3075557e4629cea4179572be5950b437d49bc538f925ff9cdf0578cdd3f317441ab2fea8cce77042bbe48dbdb4d54f30424f36da962dd3533394da2ff1cb9aeabfa584dac57712ffb6e1982f49dca6f62081ac9e247622f861f730ef22f84e77c6139b22b49b9082f8a92a334b90719ab22404b4fcadc745f2963a2837481477aa0ce1e1f6194959e18f66215e489ee56163767e5243a9f4c456f45d9a13cda5fec7977b2b9bd889fe0c26b5a7291ef3da6c217a79448788b36f08a7e87501d04501cfacf912dc2af152ee5c493f4337da1d9f14adc38ccae3a16ac080ad4897b5fd80b0a5df7151b6cc0b4796e888eccd63767c25c4768bfd96257c39ea98a8bb973225fca9c5a7e43111ce445b28a07e62a8346756c3bd9825acae312f14bdc673e38494b2aee0705c054ec8504e2fc0e1275e3dd617ea99c405418a941e73a2b3f9a8647d361241b4e0a1031ca53b70d4f550f6c3c69ee8b4cf223d66cc1805cc683a25673e1ee1b75a0ae9c16ac2eaa026c43d67c50fdaec27eea0f53552083428e54f9a654127bbc8e319bd8c5181ded6c1bda51e6e280407b6554c6f939b65b8e4582c310cded0633a0f200912afc11e39a419de03d71972a69e9d31af0846bfb822a2cccc52e2563d2c823b63f45dfd974ce00e7112f20c80fd897832654ba8035979c181677f080f7cb32b398bc911c40e1480be36c84974e1010ec4944db5ba654918c131d669ad6c7c94a14f0470cd3cef69cef4c262833fe0baefb058f0a8ba8da3ab511c3f294a0d6b2f0aef020d9135de231ec93a410afbd9bbc0c5a5dd15e6436eff8a9ef45b32c08956915f73d2c04187f794992bae301c4353ec8c39edd926a0b3247e43845efc364298f4e1ddc6d68dd1dd81145e445848b7ceea7534b4c90862b996d66dc309793f3f33ca3ea24347a2f0ee7f20bd404e04c67aabf75f861564075bd36ec1c13cdd0db244ce754689598aff2a9fa15d4c67fd3989294107c585853a97ecc5cd23890c3bebd27d29d3aae62f367853ae6263e4645a445ddcdb1edc276feaca5390d574bdb8e72bc26c394831907ed19de94f4780931ced2cb63fb8cf1d294378082dddbfe5cbd84a80236b34ed4afa1b88bfc55f94ac99e1ba013e9839876e832da1d48a1649cb64527306e37fd8c3378a986b7562853ea9b841c2b5df129d95f6d2f3f7580ece91dbbc8f70084dea32279e610b2093f4b36755cdef474c0b7edb67d6fbd22ffa71cab26944bf5acddcb2931e56b7066b23dca893f39988af8b47e00867d96f6d397bcb3555ec9fcbfee0bad4bfab94da8a104a781103a04c5d535d89567539476a7c1dc8534cc48ad9e9eb5efcf6aecff4839dce6f10bd706e29f39d9114e9180fb6a49ac75426635fea6bbe033329e713fb3823398e3686312a5c91f45791da665afd89ca76c73b7f8aef0381edd67577a01ca8ba8270f1a9a44705e107ec434dcb560198daf9a1960f4e3edd999c12f24144e7fd80238329c14fa823f907efe0c0261ba707e830c68a9efd24c83bd3ed1ef685ce715d930eb2ca4032dd04a7668e0429359dc62084b2c56c51e0cb347def9d9804cc02878100093c304608e48abca144c82726fb38d0320225807c2fb672d0a811e7e5d201ba35476a522d65758b8343db010f1a4ea62370d8100cae053ca8671bf5850e94caf20be95b7d7fe566989f3c05071fef3a0789f986bbcbb4c2ae3b76de2eb77e1ac787f44f214b71e9e1164dd4adc82d44423d47681079817e88886a3e916e80352d079625e3a6f6669a9d781cdbc61dabbd44157fc16e70b88584143c2ad4a4891788e0e0d8b163c0979d70ca222dfb11e3d3db233603c725a68619ad3484584dd3bf7fdf656b660b31c705852b5dbbd38b863911195cb46da8b9fc5c9cce31527039f1a12736b7b92777c1ae229232e1e8668cce8563eb3ec9920ef1e3f12361759c39f4afb8c0967f0f556de01f5e98e5e972e36607ea4d6add314dc85be877f96273e17e9e7a57c59a632f521d5bfd5562ae89d971599c7198980e57fbd99978a418d8594c7ffa7707df00e7bbf7d62e4dc0adf4fc57f77979ea807ca6b43e4cc5cf01a4a8e6d75f3f6735f024aba8fefb458eef6c9882659c2c8c254610ef2728dbbaa0933a94a99484be6d0defadcbf33fcae83affa5f7e795b463ef1ccf0a2fede2282c4e7fcc292ba98c10a3c18691c4d0f7fa2e07d1c96a874b11d1d2d170e1bb153f6026c9e2ff5bec342e4f8fc010babc1f27053396d05a095f51c5aa4e6e9c9bce48e49eea68e88f737dcd50fb598cb986b4bc029ec2d084682d6ecdd03623ca711b9b8be5f328d23db2b1f0519e0f39a96515db39d5981deb5e376742a87673a6fca2dad41754adfcb2a3ef8c68cebca841cd87ad0f65ccb08e5f9092a0428960f49b13b56421dace645ef1539438fc0a465426e6c3cd7c39aebcc52c51115a8fa209d16ab669fc5c5d7de0db83d83352be9b945157aa0602561339b3572fe852bc75041862e7817452c261e95492d64ab649145e13c20a4b022f06a6b35c30e79069eba0f71b1c7c6a37634cf1c2e18e4d4a17e720d102ae2051871fe6caa0bb5e09c1ec733816364a50ee3113f2af5a810521c69520d61de40427751a275ec0e564a331d098b8d167315dce7629e376f33fad0740b97dc19be20df075a2bf0535c59615427b0bdc047c28bc69430e047c4d288cd3c38bb20ec37e4f49098105344460c33422de192f6c5a08d5e0f900b57ffc505617d7c8e03e2f2f10530bff81d061f340f3399d3a361e79e45d75fc5dcc550c507bc6d8a0a5ce35ad412d93ee0861b14281cb4f59b0f33bc4c9452e7c8e22317d0dd647087631c61564484f8eebe2cee7477c56164551a8107f08505af28d15415476a727c34157cecd3b6e7c54300b287b7463e0f2aad1b2e5aaa0adb37baf7e61f8f174eb83f89bee25437e8c360ca60beb6f4f234ad930ee6d97937feafeb91b5d3dfd372a0db3d11634f51a40e892922c2e123b74e23393f277af6cf6646b11cb62f3dfee5706cb31e08c60973d994de9453650cd1d6db470812a9a98aa4658740c172464dcf91ca61e4d404e763b940fc247c3df7cae6c7597c36dcc88d61842b2637d5c6581683f0e608f2bfaac743a084b4d55fa349db933839d0798c1ca7bff66b94f30fcf86454c75affc5234db46c0ec8f7f67b75900958974fe54c313bf9fabb9c81e03124fcc38709ddec8a49067f52ea3628778bf767e6ed25da8c6e2b713a660e25de3aa1299a692e124d762b934f9089d25ae282fc9d999125fd7e208536ad7d3d993fd9e1ec74a76df3e53c51e70e2bbbab3df4043bc08cf0d82c153ce3a1678d29f2afde5c258b308f5e4674e7a267bb862c0929d27470603c61ae5f7b6af92e090b1514fcb85702c82e227e002df6ff8121031fde23dee27e9b21196a489262ab0c66b7f73858695a7c6c0592a733612bd2c5a7f30579e58dbee9eccb8aeef40420a2b5b2e1fadd3382ec2837cd642021c87ae2e8808de82630cc56aa373ce7d813668d9e78119cdc771e245c242706c2cecf54e08680f657cf6a4f4c4bbd690e7cb8f6daf0f19a4ba56edc458311ede75fc6972c495ed430770e5348477cccad2810782467af53e716a380734592ffca21d5760cd6ce1074a5c61c83e2791c8aa2d211d43d39ce54c76755bf0eb1921fb1d307d4730abd19d1a61a792cc89fd6c4f3fb35f1a0ab5893075c96c11b8c3faccc313adecedf51a74b1c1c1bdafa387cd8610959da7c5f1a3fb27a8fa027bd75115d9b3d71cc100b1571053c6c630acb8761e6b028a8264bce20ae17cf19beb8b5834e6debc2a8ee5a9983d261007fba4328d109dc9c5a12b046b04a97a3b9ac5bf42565f37eb21e3a5905cabbe4f54cf4d94e17ee4d4e29f9b7ceb851602d9977809dc4810701b6e4a61dd2118e72f72f4fcb0f9b217837581422e007ce47abcaa80f3e2e25c3f928507e434500c2ad83432c89a68e41c6646bc4ff84abb4ebece8b98630b41f77fa4192198cfd016ca1695746907341ad22917222026dd946263ad969c73757641958cce2fd4d9e90eedb0c892f1c41124343b3f97736a15b981a5859d03a2827e14962f68b9548a8e19a0dc907c8344d3d8cdfa39830f151aaff9b269bc9c61ec8d0aa8873ef20a72df77f55d6a37e41098d5bc400fc0aeaf3676dbe92e9d26934989e350e5d951d120043a6450a7e5230499d3cabde6d9c6b6cd86a0bd2ed36a344d66ae8e3e10b73f22945b9eb02549a6d940b280f2b1362c2d706a99e7011b31370c6c003912a077c6562597f33ce7c35e86c32ef51b359f913ac163e68fd9a941814e098b71a761ab3b9180a8f6d1961bef3f501b123c7d1178a0d5ce5cae63a6a4ee663bf86156b0692737bb442b6465b781a001fbcd0d03f84ca9ee7bd3b964f747e363a990fb6b634ecb092c6c3c8a80dea7e30e39a4c11769c1978134486482d60dde4eda2d0efbe95f89327d36dae444018a58f32a90e576f27da0991d70572b524c333876045002a6508fa5defab3162e57d292321e5fa5a5fe2a8ef0f9e38cfe7db9a0ab6f80a7e4b8946d70eab25d196a3d4e7af5a5255e9f4a4cf5a3d2bb1e4494e61052b5731812e6e4af02c9cfb23d93868a2700bf9bc8a85ec29f5e5ceae79d0f6b27fb6157019013c6c4984d9d96c4bbdd277934b0384b3c6867f94bf97b13c8fb5eb0b43a5056e7846c8d757f1e6a02d62339d9960059f59be276d4eae6aac2906f6ea84309b8fa1ec619fbe569a1e60e54242a4c216c54a273595938306e4cd76302b94ab822a62ea434f64680ead0b192532f6e33a7574cac96f9d3352d1cda02837a27cdc00d08d70d6d805b0bd180a3beb848a3151bf2f02bea62cfde15b80e46fa2eafcbe423c9e69569c6c67dda361b651096d63e32b085e5b76842e17c6358a6bad5379753059eb45538cb0f756677dccc5f5baf2b5f75d8826031f3189152a548b4ec0a2dd1d4f54b47cfbe11046d9790c11629b3131ff97a1060df9ed9b83f08a12a5ec0e2152facc734093e6ce1bca3b8408d79d7a15caf9211afb858868eda04d9b4ec46b84723e72b33e63f9371660eebe9fe387d87adc2d8209c12308b53cc015144991620496c2488afea6357407b21a955a77a868878ea75b79d0abf7f83ac3cd9fc5474be8dc14fbdacc10d0b936549e9776bdcd7e30f0fa43dcb4cd4d130b743ee5acee0fff78a90625a8155f3b290929ff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h832da2c1e81c0801c996bbbe3a1bd3a78db51a6bac6d2730fea332f462cb8d637fc2fbdee12e11f7cd0a9e424137dee2e559bb149d680bdaa7d4f575c75ecb89c02ec118c6ae7d6bfe9667fa469dafd78da5fb48ef3b6de313d83a58a25400a11db765e6f8cb308096206fdcb8a1c20091eabbee8225f8dcda7d6e0e647cd7861fa0d03c4752d2757d48ba6d3ab25938ecd107122c4989cecabd02cc28202f5ee82f633dfaf191950d67ce53854481b6ce50f7159604f1960f69a082dfe84d644909e72fb6eb491da279b0c147fbca33d0a02e0f26407a3a38ef24c7a501b43333c09be44ff432ab10585eb2d695df0069709526b29b21de596e5c86c9d7a410c19b79067c01d9336121f7b0db99db09171b493e475e3a32ea08dc9159915a1ea37fc18c2e4d60fb744a8d111398fd6cb68b8e78ea00a580c6cf99b1778b80867d0e52adbbac419637e0d3f5fdc80b954bc6aa4af012b4ab426647cf0ffaac513af19040812666660aa5ad01cea3ebb13fa63801c93c3a3be9aa2222bfe98dcf1862483d28a7384eefb04b8dc03d74fe8824ffd02637eca41a2e320a23e9b52600f2670e923c0f6b563cab65c9f9c83f9ece435ae20bae78d0bfe4aac2b93b6b6535174435744928a82c6bceacb4d2dff17095f2ac73cc2fdfb0a658870afc2ad08ff02c9a844a96e08b7d91905d45bdd1edcc164ff2f7aa1b6fe502023a556d36d9743a6b5b36e17534b3cfe54ffa4a09e2346ccb03bb077c2d5ed2a053919a69c4ebff1fdd9f76f83f5d7941ebd15cb49f1fb8594192726a6bb7cf9556a0616ab54bfbc5125fe6647427b2768545efd2fd1b6e33ec05a0c68848744e358bdfc3b88a902b97d791863a264b588d273ba35dec7444d28c2802191b6679bae9b0ee0444cf6187c66fce5bc56edf5b04a75be9a78d38102ea9305ee9e9c26007bd99290dc059461f8cdbda7fd545d89ad250cc17b6753cf5ccd55d1f5cc21208076327cb2c8b6feee70de880a70d16c2aa4d09bd8d007b5d6484fd8ee910528076c41e6713a9eff49e3352209d4dc497bfe90b4deac1d900ac3b0685aa190a9343bba59aec85907f736af1081f96b907dd0de6a842d33fca12aa9a6d7f2ffe8383bb5af70afa654094e12584ce5c51696d3965cfe2360cda5611c652caa91ac587acef08b28472856f973fb167adad1ce399d6ef95ae80ac208d371c90e3f323a9a9602baaa00aab1645a038b67644cc1b259c4c7696a5ad977d75b7af3513ec978da06e40dd9bd14e36093345457f26111c6515fe4e045feb1b262ec8ede0dd6d177399d5421fe921410e58ee525bda9ef8e1a0295aaaa6c169967425662f8b50c8697efd339b794c774845faec985f3296b9e54d60af7aa767f1998eb2740ca5b2c38f762b3204633b1bfac2689e374bf7f01cf2fa6a6ef5cb3c55ee8e93d4a411834dff195725058ca52c863b1c96fa2cb9be58ae861fa6f09eff7ee0c6230ed49ed1804eabe1106a53d61f2610463642d76337407ed3576fd4039c0db6293378312d5b71eef2f0ee771c18bfe52be8f1ffd31c4bcc19eb183f113a9158d2f16de2cf4b3307c6ccdc9bbfd45058bb05387ec8756061bd7b1830432d74422a0831f68ae53962744cff717c0a0e6a099443b04e5a552e25d817c892829392eae192887c30dcac6c074a15fe42fdc1f5bad1208dc303c0f67adc92bccbefba92a13f949e486e65d7052b074ab490e69505fd592bcca058a76fa619e740d0c984b5875efacb25a105ced95d34a517ee7c289ed3736048a4e2475b08c201863f39b18a7e90c9d9f785f060650630f3e9b79ce1614d77fd22c73dd0adf70a0de141377e32fbbe3e4387c9491419b4a1c9b087e9f8ac6b03c6b8da29c061eb4aabfc0aed53b46fd0418b53e3702078bfbe1b01899a7d7e4206125c20b8fc78751f8f34cb5b198f8a390cd5117ad16a8e66f8a7f67537e0e0fb7226fd4555ee93d5f85725312e667791a021d8b88cc4351de1a5980940ff2343e67920401ad4d76a93648747d177dd70a7b0f897f0825f04016d1aceb5de23c2c2ba0289f0d4277cf5a88848459b34c7ccd8582f26d924c01babaf9364c23ce6b3865ff04df27ff4737ea0ea630f326dcf3752b60595f3a56a9b6e0a94b0c57cb41890d1b6a9b5da56cc5a96e2ea003d54b104830d151dd5af62f81b9e2d009cf4fa7f7a4fd5534b3be067794efbe9b48d693ceb55f6e72fb3e102562446314c4fcda0a3bfaf89be17e9ae4cd50e4d8761a6d031235012cf3cc1c4b2048079cea1fddbafbdf3e031502b26c4db9bd0e1e9709471598221dd2bb7d5e34406ddc7826d21bfc4089c78aa6bd96887dfadc18879a21e2e8031698e31e810efb066ae1605eee78071d20f2877c64437574bd3987fbb5b7a5733188f8d3c697b3a5b7add984fe1a7098a3b1c5dbcc29b3073ac4cf3db136caf181b65e17b7bba380feb7703f2fad087dd66b305432d1727d84c317c78c99a68e0b347aaab03d9491d68bd06a897976442567e47831efd6163ee241c68aef72b395ecd26f2490c45c23ef28ec337f96447994e79eac49ab1e222717034b6880c74b094a39e35ecf11553889b6034e2d5f261ac56ff5c78c6e6e1d44f3225f9557c0a570a936af2ed836a67e76b23ebae423c1106e8530dbc8842fde3f039df5965a253d1d8c13a5c365de42d84296331ceac4988e92af16e8fce3941e8c00237e7fb9e3c38c8601816391b6a419b97c9837b2c83edd056a2aa22209654dd18a45c4d3c67eca77eb7ad4647278e591f9ed867ad797fa5406dc1ae1234aa1c3f2cbb24bcc130ebacfc918bd48fe59a91b27185fc4c561022582501fa6b545c6ae1d988d07766c9dab25789c40d394d9c6de0144dfdfbbec80a4cb876648daa43a661cb0c6442d702a057b86f66ae6037a9642eb3e1b60202c8093d6628d985661dd9dc7d318bc1c49e7ade9a23a3dad3f3a4663b7d5c2fec39d885b8a5973068b02885fec134f9181537ce80db8a4aecb1be8ff032b5ff7651640489b5ff960954c155ff193c925e645fd4e06ce768d11dec8797a1d8846ad47297f7d472cf359b36832008b9a253d1c44c0d3321bf744b0da1f0c6e7cd9494f813c878763ff254235f02064edf3959b420c154997032c5af61dbe71217649f1fe81f0e87c01d6f1687896aa2555eb8bfce9966eb1c37a1c0d5dc3d2d8a7a04ca3ac018e25e1762382fb0b944f8b7b220ff99af6116cbcb5a605e08d9ba04baf2394566589aea6fda2758a65b058105c7d8667c5c1cc033757b685c9b3636795dc55fbc67dbedc3db11d09b3d4458e09e4a3f8462ee1c6a678986a4ebc7c015312b79a532f733ddd0766ecbb6f3cf4ccb2453d2cc924840e8644d796673e7bba59e4f3141c1360e31cb7064be0c54db4a89e4183dfd928bac3d78ae9b83cdd954244b4f7dde928102219a2a31673fe597baac69bcfcab24581b94be8fffe396c70c85b642468789f2ebbc1615e9797c2df5d65aec3b50c596266c9341523017af46f2a0f75ff716906d09bc639879b10ee473dfd67494f775106b080490246dd2dae5607bad34353ad75594ea577a4800561bd36d5f2dbb0cfbaab14ae9a9fc8a7767a953ee6aff0a4f6b20a8fcc9fa0993807581cba8124c84ef6ef1a9b8012f4a84a48450dd15fb251c7352b49eab10e4b2bbf906edbfe357ad144d87ce5dbb76573f82c140ab5d31a3ecb7441a278c169ca40bacebc3cbcdfc6963878ab7348330368a4fd98f84d0c499d3b8d9fc7f98d7403b034ce5f3b5a694c6de85ad2f4e8d4edd6635bacd62094b171a30669dc6f480e1e012fb1082f7af6f3ded36fc32e010fe6fe01285573310e7cbce32d4a41d3af87cc5eb370b828c42044319106232dd865ccfa9a28f54d87cf969c39c14856889f55a86b3d072c64249d6546f1bbc46444377c99da223c329b03e369a991608e1cd13d026a7220d9defd0a617d7b40ec8b4047cb5f56697db0aa225b4ce6ad36cf79887bc222945a183158570b302324d4cd0e797a3cb573b103b93e1fc4de6078602cab59164631dd4c164a9252a61e3928457fb6af0e5d673cfb99b54e47620b4ae645e91ababed8a52122b972574b03dd53a43b0aeec20d719a4ea2d441498e5826923537d098100ff1b5cffea9d725ca7df3b95434c61fc89b8bdf93ba042acd992684695f259c890e6a79d7e233617e93d2d6d6a57548bebda4303d7ebd10a0043b8d36ee881aa7f7fca7019ca15249ce0c6e8d9fdc07823dc9d3b34244f9737a4e640b6c7edbde7a4bcc74549b4e41f186a680cd8aafdc6e975871f8bc085b96c3981a3689622e601b33538eddd5d1045d250e0b1a9a5a7a6db125b2397095d976313c85d1d68e157e328dc5cbcae0a32741099a47d7a1ef8af42ef6ce42ac64e9e7b502cc1dc6dbc7ab9d876ca9bedc0e736a7d5e51d3dc5689a45d25059c556389a8ef4991a765a5df03b879c70bcdbc152dfd38dba15d3c70f2bc988ec26044684b69ce68b5a82b11de47303e0e61690de2275cc8c1e90d7464a6c752b14b218055e3b531433e00c4c832b577aad0df5bcf247d3bdedd0ad5b7a81692b3e46805545dade9303e26391c86ce1c4539507de46fb76ee159e4c32b8bb906487f0a5068feeec63e5514b1abc444b7d0fcfd4d5a364b16cba706f523592369eaf61ceb6d9f07d820f4a77fe6f4e8d3fa5ace59f798dd4175dddd63395fb6918cc4ba435c6f60f4998fb4a34d41b19ebf77e42c1672552894400c644eba833bc464909c2a4d1c66fe7e410093f8e3990f3b9155784b6664cc8d55eb4ad5fb42bb8f0b7d084f8699dc6412e0a80553baab7cbbaca680cdcd7a3c1b23d1860c3451e4de04c5a4cc25f6ead34d0a29f15315da82505e19507fc8b36ca55ef0560a21664403d39f167c33ce4e121daa6b32f4276a2d3547c7b0fe3553ce5848d80713d9308ee6413c3d3b392ea11b0018dffed4882dc9af21c7ce53cf45c0f0b9389c2289731e96a78ca33e809873a1a224b3674d2f464ebaaefdba2c986748cf90753b86885839f69d24fee43e1d6281fac7c7285fe7562c98c8beb55b0a443cad9f19579b658a0c9f7ca7442e83b010325b0014900847763ac3de7c0be9bf9a98455c9f4c2f1bebe9a7e254d0b586c399e9998f1e2ef52d5753279e9ae2cd7cd4095304a5f86ad96bd1d2baf74287b2e2f4087e3230497f621fdeb46e4f0ee90543ce1677d7956040ce2ffde4b7428e6b25c134ed46d317f89644c168ba855d85e6be9b70255e16e304240d5e934acffba6ed5546ed6212f0c2a678148ed367a826e0d03f1c500e958f52da3498652992ce9dc59451ad22bc8b2570dc4b0cb356ea560309ad1724e8b65cc5c91f17e7e7b6fc70d08e597fe233eea17ae0835e25927e8b95fba25659082ab53c9f911dddfaff5a5bf5f4f4ae6cecf9db789fef8f5c731fb737e8bb9f60fc02ee941601aa0a7c8d7a6d933af0971c86bdd8c4a18302c5b3eac1ca19b2f905bb812f7562c70ae31c99d0d8a2b136f7fa0617698f35bf1520e74576f0c463739707f807d8318fdbdba93be604cd3bb7b4d8d01d0e9224c7569c6bbcf60d4c786b58ac7f07fbdd4023fdc3dfa786603a8cee4138855119a2cd2e4f97e4544f3aa7cee312c5914605a144ecca7bdd48989a971e8ea2cc6cc3bb8c69aebe37597caecc2e1c6cd2a63d369a24c4eed5581af7f70ce3312755e4819bda0fc5a1ee11187402615386ecf4baeefda3a4e37ee245d8c788f01825efd6c5d87e2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf4aac27f6186a0bac19709801bad3187d76ae0807efccb5a66d57f7404bc6c867dcc96a74a02773308f20cb19f200c649692841158e2cbc39f6268afd6885dc879e67637806a04d55e80c51b3003897aa3ca5cf99f491242431e7fcbadce349c55686c70dfcfbae3853861f9ebcf1b96a26c03f3f7d38e6863186b4bca665516121b62ee7717884296cb607c6c86b70b0c92070637d66e69797decb1aadd62edb59abd8a07318e80051507476c6ff2786672cb298990d7c40208aefdf1423933a17451edd4ecff17522b6b6570dbd2186a2eb6de100033337eb84a508cd77ada8d17bcdfb01a99661fe40a622f75cf9fa4d8c8361537ec27b4180c7539eebf9fa9cc3e5dbcfc115c17df76411621b6b4180ea78d88ae92dc3a21c0bb07616d315270788d276d52e88588d43ba9a4696003c2143b73f9562184f5524ce30fb537dc3d774953296fa24af22f882800eb031225c4996cb9161866261af5bb12ece9f2499995090dd870e179014135b664d006787f6d1561ebef57430ead32b3ae8ee6cc3ccce7ae600610b6c517ae36a52ec3e2178b2cd92c8ae87be93ad1770197cf2225d66588d8ca8021a3f10c129b2ad6684bfe378bfd5eadab6f09fafb4e2baec2c762ae3e744141c74c8f458ea4a6db8160c6f988b7a2fc65d3de520fa0e23568e82d5e26df1529f2f22093312de478df66127622598e11dc32eda424b2a0f9733a01fa9623897a28c309a212e8f9c74631d0c14f68beaeafa5b94d75e8c08a061b1cc6c6d84e96d1d587a24df75eca65286837535e6a7180e35bf5db5ac428bf4afb6ee637b468801785d6eb897acdafbec79dba5d75681c3a2de205c49e0e081fadb535e2426ee75cbd9686f8d70ed03bf794c87e403878f2c30b52156e380004486c16ae98a0bfdea257ce7e3b5681c1cf33bd45a1e9b19002ea7ba2e378027efb5253801426231ca4e9c557cdaac3696ea19b049a617d1acde207156669dd19890d54875b5d047449a217a2458f0bd73ca5285e595c1c7250ff4f7d85eb9471a205d65192a5d8c1e81e1f5cb9c4f790a27b0165dedfa03eba26638a198cb9d6321facf49a37ff06e6c2dca32ed136dcfd59e0843b749ee5f623e1791769ebbde9cc075680d22dc310056151fc9e72bc960230fee0efb0feb09b5a7092c7d03a205192aedca886f50f828fad59a9342c5788f63c79ddab45a3aa18a6833dc1438a89cf22063d6bd752b1a7004d4ae28af05196c88aaf56b92d5b97d2eff70ee97bec7d9fe45640b7b5d2fda3bb34388c08d7e47f924549ee15b3275b6237e2764e8c19fe0c5cb696c8ca3b4f34a0aa59320bf7693e9a94fa1a94f92d69f6ef116c1c84d9d7058edc4dcbb0a4e4024890c6f7213bbfc8d9970eec93be652554d49425f43ca569ee688bf245af7bc32e6a363a72be1878c15e3520f0b31eb491df84e2e95c845928aa30b1abe789f50fad5e8c5ff1f79a9c638051b5a88b406be6c774c5d5ef0bddb76fc3c682f4ed6e5f5c9f16e3ace2524930a52f5865b62ad3c660ce7c9b68444e3bc4dfcefc1dc65b04f93519d211d95025c8bde699570f7575465a088c4920515d860fc1f86407219bdcd726916b60491c51fb5ef413e8a78ddd253cbac407bb31255da1864263227c7514dcdceea2346e6a6422f0de5111ef80fa9c5fb94de4f8c7aa93f6200f1f37235f29d543e0a7351d51a1090939b19a95bff9c5b67cdb35891ef3c8e7d15868e651d1c45a8f9d3974b1aad206d93f5a0eaf700baa73fded9745b188ff19755550ef77a77a5abfa5122690286cc60cc99b8498071172e7ccb7e559cc423ab4e25db11ed526dbf4eee129ae0b6fe11cb86ad3fc06e9f6285fe5c4885e7f23017d48ab42eb2af1722cc1468a9f3b927d5de8be54865c504fba1df3a01dcf08a74cdf43c6b77bf14e5ed6e3ff64eee60a7b29982592cf0c9f50a87bd02573622ed862fdb5ea1255af8252167c075b4d674fd9905bd1731fba8bd86e247f7459a1bbebc216e6bd33e7e1956b94b800d495b2a4854da2545dd51f7fa246abca9560150cac0ea6df559ea23c1813ef7fbeebf23661748dae83b125f63a86810f6eb2f761fe8a77c18f4ca362db88bf4901f6062f65ad2fc1f1410e548cf91a88ea8ac06bf9e455143668d7818fff7d912ae78c117b32d20baf8175267e47b8275a3ad4d541b5e092d077e9c70b0fb9a9289e060ac40c1edc9438d087bdddb82c1db6e39758f8a4349ce5391588cfa122c9eac939726f7c43d9ed64693a92d49cf003970482e634b0c1c774e33c3e7569a4ad4a20beea85712df305f1096f956e3366c9026849f31600607109cfe3fe1dea34e711936d69fe1ff0bdaa577d4a8dff2f915d03a4f8d978c27b5848805fcf88d97aa94aea237557b0b67df6c495a8139ff09768fc21bfc6d42e5743f432507f0d9f7987966e9e52a8d6f081f9fc276279c71d6a81cef5aac5ae5f67f2abfadc17b8297db22d3ca79e47b3f24e61068c5050d3b15da40b6c16e0be7178e47574bcecb6692d0594b20a5b8e14e139df5885b2fb0f63103508c9fcd69aaaec6789da537984a1a3e2e75569c47565c46ce6abcfe63e0a5b51bfc00c888ecdb04457717481fd7715ec0ca4df81d43461b51cd0b21aed04d870f196e58da946d1befa5a93066617fa201e3a820a1b201cd1e9553ab8c9948c741da76a48f867d6e7c7e8ac69f086a19d42411e55ac4ebffa729dae589c220fbe9bc9bcec8ab8e079b6332a649f3eae506a0008635df62d847c36de6c2a2944afd66cdc938d17f4f565a450cdc57652875b0360bf67fd32ee2e1151e3ada168fe652d1fd07263ee9db81ebb78708423f6896b75dc6ad30cd2fcf72c719bb1dc724ec2cf00f868570c0129f6dd4f443db8b9bc8d73fbc0e174511a2e52461a42a74d81cc53aa744ce85ac8cb871ca51445c079324420730a6fac03124cdeea734e67f18c04c972705dfa04cf2e8889c62f75c7703ae26592e049377c3a1236d642c5f91ce1cf2f6d192f85459918220ea3321756c2b3b54340c833acc3f9b4f56e8f91f7e061c4d350de1bcd9fc17b8aa9f402ee8002cc0b17cd82da0633b49bb024d46dad7247a197747b0c48d1fdafe6e3e9ec2314667e8cc212cd15eeacda01656a7a204263b4dbbc64a500d22316db66e626218ff7ae9a3913b9efcdecc3dd873b34df6be49b7b16f99330f583f2e67ddaadf8793e5ab667c2c8526eeed80c7ae5fe8bd7c035423cd48b3fc215cae7689c0018bdaf80dfeb34af13bec41d643c599de43ffdacc39cd5e1a742342e451224f0f9f1092b9ddbd25c5811e24f28b35c72d0178c02b69af73a693b2ce3cbe4cd33a6aa9379b1e018454fc959bbc88b8164ef2ea9db1bf76c8165a7678f35a2eb7a3dbdf4ed5552e81cf492dd5f84a75109a69ca462230354c4767e4ae0429cd90fc386ecddf1bfd72e105268868733caf570af019ccfd082736207959e7c9ec78347b0598ffadf73511dea398017f49b11074e007191276de074c8702e5c572c43c56b05b8f32cd27ec4270d1e947db506f962df97ee2d5a4fa2c7cbbfdecf4a95c2e5817d41c0b93bbbaa6f7aba290483dd8b89ee1fbf7558805b410f72d61e31a69d8133b5cb2cd09b7320e647aa50552f7b1edf80fc85f68f80139582cbe1e0b28025a6a46ff070b37430bbbcfa8a46428b4035ef9dc941aa332ed00a7e3a17eb7f8b579aafcda8871065251f273ecc62b357ec9e013a97de8958f5845e300ba24574261b28f993c6f894824e271b8921cdff85e8cdcf81c6cb92c09e89ea587973ef08396dc3423d8076a87307b0a72a8494636061f96dd80bd66f7cdad12986de9f31c4723ca7b1bd9a7c2e55cf2e0d7e62b27df805f19d69e80485dac11071574c1a78a7bb31cfc485d4d12f3acf658a6f6b69e56264b1d23cd10aad2ba26d05ecec086f7b8cafd84c53bc2fe0253b3c074e1d47a1aae013f24de44596309a42234c8709ffe40a2e3bb2bb7d3ff5dd360f709a8ec471d0be82a87cd704298bcfa4d60ba13b763d923c410f903280ba3c869a5bddecf5ba2adf1e8783de84f7a56d8dcc0c8a7af676c430107aa34fb369d339488f3598a9fed71c875e39b8490731947104f8d960b3e4aba14fa0b7eab09ecaeada8f25170624e012be4e7265cfda873daf7dee4f3926296444da748f7e55472252063ecb3172cd6d77e4a24f00118e2e1399a341f16eb091255d903d15f9a538982f371b25f4e3db52f7749a4e45c7856dd10eb2a5e88bae072e390681790fec19869864263be7831a77b24b0565631d7d6b192d992dbb49575bba0f02cc653d62f7092a251c52a03ecb1ceecb42ebde58b13fe5fbecc6ad61d882289c9b99dcbdead6b9741591f74df40ad357236f5d32f5373dc74ad3b6ff25f7f1765f0213a471c4bf047a3ab28c4c892582aeda255df153e1a853fb3820ca0b2c90f96ff4fc0ff7c40e982d5842dc4791fccc56a9d4d768d49b2351bf7d7e3500df767e2f0e081b3da27c43418c536bcd5f97dfbfbefc1d7b6a0bb21abd441ece8df1113fecf63eee6468e588d414ab1b2294ec4b1480c3f488269c3395cd80ea7f3c9832aa8b06cd096381f387280b80e3c7d1bb99e7c2e398e927b5259d51fa675e7c3c5e3dee89197d143fb1a29be70e2413e9f71da56c1f31b23513bdc9c11cc7c5e2238ec612d60dc15287a7cec78b9f32bffe8a6940d4dd50d5438795d227e8d544235317cfc51171a968c164c6739ffc54feb583445ab5cb7710512d6a703615d080029f0aa90fc7b3e4318d515c604e8895eb10560a9509f61ef27187d494aaa8c60948adb1fe8f3fa505daeb246f4dda1283c0b953687f4d2137dfda63678c1035a299e9f82e7649b1195c8579a180a98896d64b91afd3ee2f94030c7526abb5221c7880a69927ab127acad5ff9946b421d4287f7b7eef4f6dc103e15b1a3f982fa09200dc2101b07f6d7f0d947f5a57c2aa2c9edf2b79eacf9bda1509f51f9fa90255291eb479c0be91e5e475e4af63a2c2a963c8727d324350b3badb376ab096c24010acd56a11dd176cb8aa3aa5794068c4fc5bcbce1a5e8046d968fc883166d3d9d58dc33dbe64f0d7777ccf3930694bad08c78af70efe797f75e9e838da70668f84054b46cf3ef85339778b4b245b4c8d9bbda1c5207160597d7a6e2d1a32b42e739810b9d4f15fbce4ba83c2e9b86c89c08f11e30edf45c513a94f9737ed6af25062127a21945a21f35a53537535f263cf8e9d5480e033e3f590ab718267d97742adaf4c8dbbf5e606c935838e0499cc9ccf14a1ca641b6f687b9e79049b5a2a1c54a91b4a17db277a019e23826585dbefc65d774f400e7b93b3ef88b6e948244d836766de5f890eef6640fb2247651520b36edaf2073a71973f4da6bd5002e98786c74f083e07f5804ce48dbfd9d187ee760f540002b9dcf3bbbe70b888ed7be880478074d87f80247b681f86d5410486d3eaee4a42b33378847ed5e135669e099f168989f675919b45bf5ff81adfb466820315a81213bbbf6bba7a6c6111cbe53e92c9c9bab5d53200897c004e5c221d7081fba8ac2cff597241c028bddbedb28945bb1219be86685b07fc436390b1e1b57db3f4af298f9b2cd9c20c600e6433ecc47bfd28fd6bb116dd3b9afc2bf27a204ac2fe60a0f456e5b35e5b41e4cb9c83f138ecb16b10245e657de790e80b73b9e26adb66c3f5a28b7bfc8baa6df97742f44f2acb97d7ca8108ad126576ae8dff2bfa8e0fd128559da155;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hf3378e4b3894d14ea5360fe680d3589038a4bfb3997a8d3b24a22b0fefc31805dca26665b307b6343e23d921939f4478934b02582c2129606634f476752fa7169aa76e388389db2e69176c152cb871148a150dfe1670c7ac3c6025a7e4300e4044d9d5a05b13a9ea1c124d5e819ecb0789e62c47069a2beb76ff11019c9458c8b34686f1a3c4fc7104dad60bb5b74f0edd847263c627600f1b4620f45f23f2236932fffe4e67aae019fe5df9e18eb544a622c848b93688e35d61095aedaf6f081ad4b985953cad36ff2b123c63672b1ef0f325db2e5eede4951b53c266aacebab41e72c45ad702d1720d030fe41e320b14efcf227aa7021da1743efe9a89da2cc07df900635eb92b7ab31aa516ff031d5e9bae0986c9dd7decdcdb5220644ef1cf0bc22de5801b9d086f6c3fc3c2f1e249ac6cbc8141e7bcfc49bb83cff8cc3a0abaaeb3498e22c2dd9cebd14111d002d7c8a6c8abf89469d07972fca58870c4cba33a44ffaae812e314c3cdf7878a001289d43b79ed47b277c99b2f550b52f4cdac9dcb82456edff9b3487aaa3825c3edce867f1f295c85386ef8706540482607f622a415e7a227d514926301db9fa522f53c7b63b53a7830a976540c5abad53623ab71c85f922d598bbf9766193fc379f36d178f29dce2b269195f3f0e37f9d1fc4bedcfd4d404b2651b3f84549edec1e89dd5a1284b6c107f01e8cd413a7ba20a0dd413466e34db79baf241fbd2e2150e86c8769f3662829c4267be1508db4530f9ba97505cb1d404bc4fb169c32756f7c7ba3050f19e1b3449bdb6286ae22a6c842e625129c8f57e266d227df0d75e83211a1d40c8270604e19c64f7022141f8930ff9206fac105250c3c8a254d46fea5f196728210d469533d3e2dffa70f227979ddad7c25a0cb6a47a358b2a34c9f600074eaf5a5b755a56977d555a183b40094a0d4a8696e74e72ad2813ee5e78271a2659571c7914f88f10e1bb8a9880cd1a423ab63c2334f0ad2043b53bddccbcbb59881c1a570814e81863c02c4dffec2dce9cd5113ba43f045175267a3a30965a6a358c7004476d02db9c81572002d2691466dc2e4425574d40ee11a27d2f39c37de72408a0c439a6bb329bfc4e1297772fb2d1f521bc6589b95a385be21eb5fe06282433992bd7ed71eca5285a217188903992fb53d40fbb1b7294b2269d36839f610274a025071b1dffde927c9d04b086ce389c7c5b85cb6638d5c15a765d0e9b843ffcba4aeafce5bdd9687cc9202fd3c238d761540342f942079d3af5d7be53bb9d73855d904a3feac1e6e072e3873d2ccba9bf78c053138c94b97aaa59c3fa2e666e13169e0e31f1374e8230d128ac90197b5d98f121d02d39e539cb0db928f6b7eb4bd1f761ce1b153cbbab31c5b2226d69dce8bfbf519680fea1c186dfbbd3facc49cd7245d42ff078a3e6858ae67fe68a9c98c5da9cd596201bcd2358e59df8950b617200d00e72851e4added51c8367fdd196488b288ccceb895cb7096ea69233be66cfe4de4fb53666bb5aa0046b40ab001f6c3e655bfc737e72d9724cc143cceab08786972898f1fcbf2ae119005b54a02285f611053e193d3fc9dba9ae78cd15539c2607854fb83612cbaf790752145bcfe41a222bcaff79a84353a893a396309f437d82e87bf67208f9b17f720ef54c8d2e3756375ea55a300095b2ee100d6ade7bdc122866b3e8e70ee3d5ad9ed048811940e1e1e85565c9a041f6fb95c6dea8838f8c027ce4c0a64ff6bbde2734b79146b4840ce907046c776ab6f099e23ab103678ce312edd0c80ba7137b558e5bcc3a7dde3fbed3ca7655561c44ef29cf2c441a6c1c6f0b06e065ca5bd231538c4a6b62948179383850d33b45d541db193278519b2c4b60d9de1ee478066cd46e4504f1eea3ece03679a0d5e48b52fc3210d31c851331e7d093a2288db81687e67a5303a5d4bbb03e5101679813ef95b6de6fd0421ca260695e3d26ddd294882afb7ec3b009a201f879da3c4e28743b00999da993e89d916732c93bfa0310dbe32c541ba6cf2d6811b1bf0d8a09e1df8844cffbe22df5a907b283ec17357728ea18715a5bce0419c1d5131fbd0e1ea837a659555d8a48a7d64a984a7a2dde1dcccef6d17acba56ea3fd06de6c6c04c6f9ecafc9dd8b5828210eca8c246c3f1f7f2e9db2635bb129898ec427f3dc6dc4be03ae9ada7bb773ae9ee343211bd4640b31eea5cc4967e12da087361db6ff24e2c46f3e5b29fb08be3d1b1069f3281935380d6ccf1a2aea185d0b5ab89207ddf42ef3e183d0ef6ab0c4e7fe382e015173fe24d08a2137f6d087ec8c699be7ae4a940a7b5812627754e92548ffd61d638a82e60dd98d1c5ad96786cacf920928ef5102b5b88410f083e03b70c21d205c5265b15b432aac8a29e222eaf685124bc9ee78b8e0548234255006a471a73fe01f0cd31edcd530dc5375b165198280effaf2d061402b5d39202084f4523b857c5a04c7e80da68c117dc8b65604cb1f62b56563a2ecbe55f39427f57c7121f11ca3bdc0f79cf7156ae62821f56196d330ff2b6b79de09200f1b53afbe7bfbfaec8ab7ebef66a37cc082bb857ece4a5fa9d7432851faff5d41d2a3740ee9ebfc139732cd6e75fa980920b6c334e4677e1cfe4903e2cb5826d0e083abbc6a4345a22a06fb2ddc6541f0a6807543c380945bf430d5845534b5b56ea02de072af8d68e59b9c36fb7240c710ef32af83ab92b71f55b2e1e3b079f29a85846aa9348e0fdbd346aa46004ff7d1407de5112265ca1fc596e1cb5d60ac887eed544c1ca592645950e3f52c70930419222c7c06be811ae35be63650f181aa6ed19069b8cb153f81fbfcafd2957d736f6c5ebb93f3686d580a064ff1aa9df502cf307e39d666bc406ab179c6633ac6a66b8a9ee7c0a37f558f020edf80e73234dd0d50b69ae85552c36dc874ee77452bc9cde34c80763a76e3e3bcc86c76401062ef21ffbcc5246305a87bfa0db8e96b75ff26c66765927552225cc66358fe1270e48137f65c1b8534b046e610cec061ae76efbabfc2b4d1463fdaa4489c624008613a52acaf4e2023b5ce6a402d5f12209ea801dedd15c04e2460d243222256ada4450fedd8c077a136b829054469662999779d2f2507aede648d90ab803789306568d57f2fb45aa4b499cfc8e8f4fa651b585d5929638777cf42eaab819c238f965e306c14a4672f7d03b0ebc2471cc55074b6b816e4a2851618710921d4788cd177b9f2d5c3e64fe82aa17fa43e06c1aa6b8307143be8aec2ce7e0f455df3ef48a66f544460df8c35c98f1656aa3f7010975f3942906cba041c34de059d1025176fc5e7a8607ee8afc2096cb0020b3d12c9a50edb43acf0de83f2e0c0e2b945860e16ff1995526f03b01a3e63387b73b5aee66d72a0c342a5315348b99c2038175701516a1f54f920d99b1da13923e3ed7c4d2c029ce69a60444207d91662d85b6a68571abf18097f0503ca4fc2dbe1caa6b0609a8c1b380939c88e058edf929f7280dd70330db5fdb44e0002dace5c96bda7afe58ea3035a12b2f8eef26f7949c7c39dac967fe466c908b2ebbd313aab6138ca2b06bee330b88aceef4ec1d1b5a5e8487ded38101e1d273fc85fce82fa6d5065a30a59a1c113a642236c8cd00c82d3d0795e9d1e9a49e883ce1d8d66db326bd6198a9e36cf85acb320eac27fc533adbef359334ba1349bd15eebd26709a2850acfe851994d403d7c8151f16a4ecabac0da5a3f3af0de8ffb50fff80d0665b87e44d8b4c96b11b49d71124f3b50309659cb19db28d35810c0de410666b25afd7afea643c106bd3fb0076e5f3e2bf8316c89ff859a4d3dd9c63f8802f541bd82b096e109ad01303241fc600f0e460f2f14166ec03bd9ca8f0d96fe5d1fe108b143e376d127e84bd6eca9526426d5c68d1f932a0102dd1404c6202f1bee17438c653f6cb3b084163708d44e644e6a1379b8a8c76c8e299cf7412a225e86eb0ecf65f9f923535c814057fdfac4ecbc42b75fd9dd083bb9a77ce2df1a7f770cd3e69f93034ec2b9e647bee489bd5d20aee134937a631f4aaec4fea1b92739459c8a6520c743ca071bd3d31f1bb2d6c187f10e5535c5ee8900efe46d995c758a49e4ba8d0547aa01e4fea4610014a88457da7ac5fd7c5a3ffe4ae919ffaca087dbe3e2239a29a62742ffdef793d32354608c16dd5ae262a64492c2dee1b419db669f536916fd29c1d06fae0e165c50afd2f155c3ee746ee178394319b82743bece11cc4225df771c4306e8d0c5e5df2e055661ee9b77a9e7ec80112c188d2fba4ba68c74dfcd5017ec31e02f657966982e600d80042007788e6a6a5e7a12b14ad456752a672d3c5c74cd6bc4cd465c3e68b48784399370eeb5924ddc2f8932c58c62d04e9ed61c9fd7a1f9543b6f927e810480549ba30d1f436b07ef06f0aad31ab37b0835672a3a2d7608d8267073a8f74c96965f2b0af71ca14e290b013f1b8fb87f41094bf7d8803548a37b839b32de4acaeaf016218ff324a75aec2e01979e4ff345b424b569af6f66e84b5a187474255c1adf1af7bc63ae25fdf6e10279d4479855f397ca9f3d3cb998071bca06cb0eacd8f7805e3cdef0bdb9431781d067e872b2864fb0aaab44dc096a3a53b0c9ad27db74da6694d2dd2e4907f79e262b3808bd20e18175d84fd848578f773dc35e729223a8833090eee85e08fb6c622470f1b3e2bee87d88911cb427a4355f05cbf853c9ed0550f8d48164b30ba33668999c6424b4e1f5ab3b9d72f03c959c0be60c343c30f5547b0ce4bc695361ac87547dda94a05186099fcbc7fb8bab923124d0abd750051d8dfa7f1e28d5a15843d77d5dc986257cd86c1a670de774393c0276575fdad1695dc9fa1ac7730e911a8199cac967ebf7df74bdf10b3fe088a000cbd17373e4ad2a912536acd5358270169ed2a6c4e6ebc398d509db3cff5b1ff5c9c20cd6b6ea4144e530b57c9e1607be3843f09036f17ab4be2f563c0d66207b48c78da782f0e1d863a52d325f474aecc9725f74db645d47a6454e5d5b39b723abb2f34f553c3e973d7b1612377b72c831a16a9cb1d815e838f40b86a05205acfd9e49104c6c663535dfe1892fceca6acfbfc8c773f8fa82dcf98775f3b07fb6752210cf6fde00b69be64b27101cad7829f070493fe07fde3e44dd9b4eab7cc92f696a1f8e93c28e0189772660ea2de6c9db3a91ceb6ffc420f9e96b62c647ab1e2b9b780bd309e2227576a0e7b877ede993f8269c730209e3c38c8a87f8fdaf0f237a01bb2f0b0df6dadd8e7b24fab43d655e5ae0df01862c8d069f712bb34815f4570a93fb2d804fea776882d01bee6856331debb8c244eac1e1c59f0695088e26a1954053e4afefac03d2bdbf4ad39d220e353a26b8e638a9550d0aa21c6d3d3e7e707d40b738bd9f4e048328aa5b0cafe63dc5a1eba1ec8d6827786dbaad8deeae0bd5dda90a29ef303a86a28fea556256ed74eeada1e2a210bb92a96b674663d7d2488b5a8075c8f4ef45087f0cd363b3cf4b090fd5ae6012c3d321129d0bbdb5a48840efcc8e21afd0394816ece76595733878c1a53ea49fa738b2aa02c46510cf4a3c3f2d43ce0dcb115d19dedca742e069b4c9f76027192895b1a755a00fa161636b1b408559daf9d9932e9c6f174cfc3168044a83226734573efd5557a4451b9683f9b046efa59e7686426f333eeb7b4e4f7249fced2025c4143c3800a96f9d46a77076a7e7ad392e34ee305e03a0c1ddd8558e14477;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hb9823bcab5f161cf7499c0877d6e112a410e0f6fe8463c65ada46c3639bec44d0b4e3065b2918e564d1c9b8354de75a4f5eb269ed573c39571f791ed054f2e828e21c1e595e5112a49c4756495bd23d73c7aa6e13aa5f0b14999cb529c1a15314dd9e3c4a6aeb867c7238390e8b18ecefc009216c7c4aac92de44f3d1865ac3ce7e7aa7c0552f8fb89a6221b8c7867e51390596d52efa87eeadeba0ba5bbf74d8cb85e9f8c71e9175ae476514236d8e8422b944924178d7f02048ae3265a607d375e208ffe4cc11d62ce09cf1bed55a5c24d85cc762d483b54597f8faa863671a511b67a3a95c423c403894a87b6b66179da61373d6d7179aae805edd2e5b2b6b614522cd7941b1f3d7cc3183fc11ea37f5a069156d2a9e25b2e8b69ab00f8113c1516375a9d3bff1e4b22c4ff2f52ea5913d04da533e37046bd51cfa5e6de1a02b29e0ae42c63a2489778288fc9bbd06202733a92c94945524a5a4d6214242ac7da5ea70dd239721f210f884f4b7ed53b081984bd7151f9b0e859ab18e4ddab770c4d0d69f1509152183fa04a73115baea73e2232a5cf89698e8a426aa8df3c09ecfeb1a45365be47a8ce2c1d81ddafb77fefd7d8b449e51f49fdd0e2448d0c542bdd77423eed56b972f33fd3d47c720110e7ffc965a08c756fb17a35f67ee22acabd11f77d37ac67da5c80d07c3c719a95c106a5095a38551c8054a164ac26c9e6cd536130fe54b959f933ff19a964ff9a08c33a67148345c2b98a1b7340cab483642119acfcdd8dd059668ff44d71a5f7a280d15116f6d22926b02fed0959cbe1cd276e191a1a1838468ed795c5eee18b006a033a86f04afa28569ff56dcda7c6c3fe39de61a5ca6e1b3e5dcdd958847e7751732e79e787acdb6a9ee6a6c3c5a3aaa0c379030eeb7def5d7a7a6ac95081532687a20d1cd6b3aa02545d35d2ec04280ba707ff14894fe76f9c29bc4e210a52badb9341a6d5c17b0b07f2118551bd990ded785a1b500fde90b2f4752171be2648d6247cf16778044d7749dc37d85c93e1f983c249794915643c211ba61f18b3e97e292ba13ea69e4211cd742762475426de6d5042a1beeced1b25ffc06d7d3ab379f61311889afc97b533164bfee4d6c8e2886c642488a768e2321bd960f09c514a738d22034e5c92ed95d9a832c846246d4eaf877abfba8279e3c171bcd9c7cb258682195c12084c9de5c2a7a2a1e867e5979c85efa2b0667f6bfc2b836d153145e3c42856f62d48bb4e9010accc81a383cf177f7f8ffe644224037e821eddecae362aa6ba8e24b81a5ac66d29baba89c1dc7274a2c622c7c71160953ab0ceb33cff7b552eb9536d02e0e8997107b5120eb3e7d9179669ba222fb2d99c7b7f7d7f411eb18cf80373493dfda4d54d4bcdac6e2b3a5e68f81c7e3b2a749fbe01a878b345c073ce15553ce5dc4ff2b687bf971bbb0d081228df7fe61767dbbbd908ee6d31864edfa0c4cb27fd9de1a2988f0fc2f55db5b3e18515ee0da3db282be3556d9ece04f6e1ca9fbb68eea4777590e81642769bb523e33be9b5934eaf598f61f2aba8abadd14d9f3ddabc78756f0237c905a463dcafb300628d91158ae84fdb6b6958fdf65d3750808958abb6f4f9b4bdf2994dfca454f41a28d9d480308c2520c4c18c342123e62f8a6cdeffbcaaae44dca4d2ec8c666e0a2308224a5be460d63c07a06154eb9f844a349739dd0eded0bc1ddd82feb7556cbd3440380727ba55e70bee650993d4a8129053d56e3d9b696eaf41deb805f5d70bdd9a63966b6b5fe8e34796b817ad5da1abb8c47a709e90907252ba9274cd8349f013869c8b4cc0f48b48de694f7041a185d1b5480c56f4d600db28996341c51e245f7f1a1506e53d7c3c4fe6017c107be848958a1c11d60920d0efc74bc790390f0f08989cc7ef18423a1247d9b31872883c8c349d7886e037cc54cae7d7f0d8c77cfb89b2e71ed90b306f96edb23363646fcb066fec144bf8702f0490a9789865db9cb6b969d9a146dfcab33883d452c1a33291a587ce48a068c3bffb2eab7d2d11c1b829a3f82d339c6398a3f3a17d2db36c20c7568db84d2d274561337bc22f1e7888a50455ce0b1c04633bd5a45e043f158debe01883fbc74dd0cc8e3e36142db35b4694906e6473620e5da1ad61d8ddbf52d2858fea02b73203478db51f8720593524b3608c87af05537c00cc58eee6e4190b0106bb0a97281edcd3f65d09dea0998ef2284157999469ab66809d0b133c538198d1f059904e885154d20e5e68b71fbe621811fb1115e7302b30df0b9078ba899dc163a15e988ce4a75e21411fd72293aff2e46b3b7462237cf84aa54ea03bcd85c67bae6c22b5a71402a6a01b8ede76ca8ab97bf18ebc807f97163a7beabf79c254e8481f50636ea4ed7984163d8736cab6d3a7824637ae7275bc4d7e1df5edc6ba37bd25eefede33058e28063d7991b1c0f524e4aa8cfcabd954ee0af262985dd69ef24ae30629abccb8a7b9cdf26777e7c3d6596a8e64ce1936f6b7a636a8454ef50cf46bd7c329e5894115e12a1002ae36498935bc171c7b4db569b7e0f05a79a2d1a6f6a3228cb3fa592749455bad1e94cc7feb87d74e7db99debfc9f03037bfeb97e826df91edd14bfbce92c0fa72a03be50259e0267dadb66f283022564132bce2c47e9d252c94f58f075eeeb5ecc135611fd7ceadfb2f4941659d8a48fb07575215a19f6c0c694a2b98720ecf61ba0f5d5993919f646fe00dc8070a135c98735c338181d0a6881bdc5b48f38138d19834134bfebb4271c9dd873ab501972dea389398f28ae107d77fc2a6b2a812b08f26c4da048e0d103501acac5bf9344226ec30d91731f60f442933dd201109be9211f7b102c8c72ef15dfa52b418257b582bb1c7d9b02d23df9855de5a8d23601db34120d26fae5297395b8f0210e6156954429ef988f66ec5108d5148e096f9d30972ffbe5dfd541a3460678494030a5b7a3f7826bb72230ad7e078c875827c00916b2d9d46921e57a8fa6e400ba3f2059b32afe907bd74c5f0b2e24924b96b809859a244ba0ff47f8a3609ec37523afe16f6e747e306c8ece28950cc6610c00576fc95c2a7092a1f01a84465193e28ed265637084b2eb5b71e7b43e71ee88b52fc915995b2f53670d8b6220abe20752c1c3feef606fa154f1219ac37d958947bb0789f2f7bb47946f357357e24cf6ed039db13c838fec168e6b0e1ee171046094a487542875722f8fe8a6f0a211598dedf019eae9fd9816d110cec3da6bb448f4339139969e9911811524b4cd5d5665d5bbea3286669f425de28c28d4012543064ee5e094f3bab543938058bcf88fe394924ee0967b34746d2e21d9e4174944a47956b65de9ff59c8a09ec569b6fee8151f6fbcbe7763e40a8fabe3355a13798fda8d4f7ff9c03e4d658a4a95c8827b88f9a26569861ce909707279b77c4bd008df7a2c17fe1c5693b7e9aab58283fc3d5724cbb2606d8f660baac2b38ec7f42cfdeb45921963b0f1ba14f6a745a241ee86ca43e72f98845b94f8380b505f253d9646962ab6fbeae29bae8ab037ad5e3647ee31dad7f793f6b1b209d9d4688751655b77d88b654a359948ce324889cdd93d3e3324c56dce601e34e79238884e9a1a618c7bcdddf1e7c39b54f09ba626920d3c5ad49a19d9d4e1ca5226e7c6e47dc606a9ef466adfbfc6fdb73e81bfbca25a277118a6043628fc6b46ccb46b33aa73a9906d6ef37b7d9442ca47d8bf195440a2d38dbc449805b753ef3aac323d3d709dc77fc44ccfe3191aa6016245f540860aeb61bcfc97e63dad0e266629f4075c32b3b672240a66f8845a7756e912ab2510435a3aee105b8585530d83fcc3af05024308afc9ee8c8fed44447d01b5cf929198ccdb8bc3a2c60bff96c5919459db43895a6b42e1a06184cebcda6a545261cee956e6a4d502968fdb4893b099ec8aecef52b3f36b7d8acb5a204490261143656c89eb50a255f5a2a8975aabd2ed75fa0ed7ff31962da2542fedf27adb65163ffd65d4a1b4dd404aa5da976362d78c53b216ff9752cbe03d9e01919ec7cf37e4c706be5406bab822f29986e81e828cfe4cc0205a95bada58d456649e3f325f2029f3d3ab99a3ab10f7b441892d4d4cdef7edcd9243dabfcae17d23e6585e9e259d2efaf13c56ad8af126e1102fab9d2eb9030c782e2eaec7694fc604a367336bb1ea9004dc053032b2c23bdc4c38f5348796895f4ae7f099d138e7b430c6f00d134134ff758fde5982f12262c1d9673ae4e649d18ceabcf7aaf0c3ea9444f3bd2d810ee1afc8aca7af46d98afa58c0394009c2fd1b71c4f26c61f036da226c40e161bdde683c575a0df61fa2f7d15edfea680f620fe379e299883bebc92327a2792674c938dbd4a2250ad766b619d30d1aa0bf4b4317a1b1b43a0fc2b1cbc8e4c1ed184062a6693d2351089e2aed1e7863b90a9a0d5a6b4bfb27c7c842a277313e59722410bd9c626f000d2321645e83d4d63d872bf0c51f497908216f55f22f20597f39208f1b73c2834970e2d86d308d837831244d3f3776d2a454e2c537daadd78db15085d748474e7081ba48c945f4a78cda0d8abeff19a697f260cb298f70a4c881b25505645094bb732917cba9d783422da91737e15a877c9fa235f5c23f2502a270d294a81e82305d89a08949031063b21080924a1494e5463a22169be80b1e2228d05e32faa63ee40a34f3a315f784f3fc98ecc438d90d5e8915700bc38fe571a1faafe8454ad09c44e1821092b0edc9a3b0d6eb8761298745ab11bb3634eb18f6d4f3861a9ef22c733051ff83a42c8729162f87ff67055913acd71ebcad88c10c9874b24f1313e1e9b06e995756aabce60ac436dc9e0cb224fb9c0ffda2e3d17e93e517c59e63a35d746cac29fa039b599ca0e5de16625c4ec334e11ff56d04092cbe689b35892627b67dca2b4cd2d369a5e8cc3bac2f9caf25d99d3db61bbbce920e92001d4cab325194d9e938b5f4aa7cdeb05e5cdae19c2ba2687f757fb67f97acf45f8f01c31bf28ed0e6ea94804bdc619e93407c4af67e00bd51d942dcb237ec2be02aa69c29078db6d96a41bb1464198163d1945c5291e80a96e733270d132ec2a7e484fb1605756da113bc8253819f0cd8d0f5aea3823ad85c4c486f3745b662de955adb7862262f01f30a1df12fa5fa03f0ff70c2b0b7d823ad545a7fd7a8ea4bce45afcbfbb88600b44b749b8459700c839b2b297778ed06873edd44008597ad195cdcb60e15310e0dddc166a7ab01bd0a7fde80cb558d107a4f7d9db7f4a41ef695a4c85ee578497ee9e26443391cbebf9677d2015afc242f8102d1bd4bc4f4f50b6bf27ef0cd5d20af55f59222552156e1205a8172ecfebf2dba5ac94b78ddb215d351d0ac6faefdda6db85a67d3dfe9b45127465e1d1afa0559c104902d2216ba88c0f6d671fc4ce9fd0f7bbb96891f13c0ceadda0a4774fb5ecefbda75c200b6b0c2b75187a56f9c3b0649c1c14ed9f1342b4956fcb13ef544cb31300dca78b0438a05fa44aa0127b9dfc85c03a6da9ff96af6ad30e98a9582be095410f726e7e4f560a63c819df82f28602ad914a1ff7118f211f2b08e0c80312bc2f6241db785fec1246cc2186a277662e904ee05b84e41a9c7374950d03407a2ffb63d83895c3d0dccbbc7d8db56bc212bd19d60b5a49c58e1cfb626007be941a86674b87569759b6e60d74697f901602e8d8c94939295e1c1c16dda19ff5ff33d645c3528d31f3601ff378348dbd0d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'h331b80bf585af0c02ac30f177f8487ea5157bbd1610751c2d9acd3ca20f244ef3a00df6b2e8c24329e74b46a2bfe793b14193a5287f9f6ee8748438bfbf5fb587f44b09b580f48cee75059968ae5c327cbea5eb6bdc483c811635f9c67d07f443c23804d4d50e0f5318df70ace0029bb3824327fb2d6f3b52ceb2178c20b1746604d682c1c83ddc5da27c3ce12e622a4394b9b9bb2bbfafbcbd28641eab66ccd1a17833fd21773084703ad19ed052923d6749837bdab8cfe7261261bc674578a55e773f90c7011c883267c9de7abb0af61c80b7db53a0677089e5535e322925e137e5c445aa2e88b9b5bd54c7fc9a1a25b5a54d6ab6eeb734f7101f1f510a050850141fb02eb092d25e1d74c28730a84fea98836892e5b86418936bcaf4d1f6531a496d59020c5f3ecc75a3d919ae0a1d1a9f3a8c7954ea2bdd90d392d3c5c90736ec8a3f1458c7f6aa415d05db7884bc3d884a8db847498c4c39df5f05cfe4f953d4acac78b2c1b0aa42070fc9b13cbdf7eae0afb69f3e29ebea479695d38f4eb0508d84b1d2c27c06111e3b5ccfc9d52a99d3d2d23a9badb63da58dd9a54327109f469b451f70a80ca2dbc8218cc8267f8e40ab4838bc241979a83771fb1569b36eedef5b867533e35a7ddd09b21bd88be4500af44c34ce3133b9cf52c9c6d9e6b187f5a1e6595d621d01429202b4080c2f197f9009b42dbaf045d2344c8a9b9bc8d7e8edbe6b5a229fa75aed763be72533552cd27e55371eb167f6dcd5ea2e0256a2b6bff02b9ae793e5c4eea5dd2d7287739894aba74dba756facaca7f94b94d22048077be9ffb8be4d6b406ad05b5244d1b89364cc7fa3664c6dfee57273e1fd8a634981c2b36cba13958abab18dbfe807b6f4eb6a6c32b99fed02b4998e6126d224736c7a9d3c54ae13d5414aa285d811d777529be172607230922ab0c5d19f8cff380cba0dc3c02c8265cbb06128ee0a421cae9dcaa12d91f808f047d15eb236beee0697de1ff918b62531a99d67d26f77425731280c7086e280c0bad83bfc968d9bd4bd7d898aabf1458d76e7c055b7b564b7aab05fe0450c0d545d3ce1e367f56b4dae6679ac2e7206a859aad9c31d4a30ba4848b261095fd4685b6c8658bc52f81c4294a6a3b1ab7f8ebcc61b3fc0c7a53b68e55d6d7d7277eb5eab620640eb211a96568489c09693cf60560b06338a10bc0b43715e7cc6efe6378121cdcf2e1a90c792288983bdf4df86a5c9e8a6da4255405a4c3d48d51a958de30bfbdc6d5887d21d577f81a33a79dbb4826a3f83ac5aa68006d195418c54c4ea089a04ab128d53ffeebd18bfa907299f0356d1ae417a6ee60cd296f91fe7dea7d78ea66268ba156d939e5bfd834afd18a683200bd41c47c988cce153e275eab69d7dc470ac4e0a0f4b146073213aa8faa2411460bec67f4686223f732ca65987b81dfcd86ce6a64c0744d7f342d30ef76992910dfadcd383ff28ac7180d7205b97b26191f78d715d4159979e8e556a05c63c2c136e2f88e3e529c6196e72020874b9540aae70a3645ce685c85b061218e7f3c320123ddb6a9efc4e58900205b7a539346966c864645fee6437b559ec27245e63c7089f3ccec7a03873958b91d4e507bf509286fc4b244f812bf68391b56676aec84ead068a6ab02276ca19c8aa1d3fc5491f264d4edc49aefe4b0b5a4fa5c5537e53035d0f005314da39d1705c0a2c25bbf3f115320f09df243fcd83c8ae429747b66577fdc545dbd8e36f6aecea0701356af67facff4064c9e4c9f2b62739e6551153817e63686db303b17cc293ff4db47cf9468c7dcf0bcd7bcf5c1a34b6362055fe72116c066533e62cdb6767f20ded7eb948689adb83f424a5b13d83619c2262816c6dd2287f34946376972309526989a2ee10db23a49488b97ec664ea4c320c8481277598e685376c86e73849db91e55f07b8972d7d7f9ae92fcda42bd5aee665059b681cdad2a14f638c67ad22d9d2cf035427505f8c83318e12fe0d4a5ca2e8d8a2abb58b2314206b4e4b82158950478754606cfccaf87a873d7a41137dc1fd33fa899c29eeb075e5f65e34668d0ff007f5068bc0a7b9caf0ba88846891af47d6c723d08c1a196478c69d5d62a256f68aabab25456efac900a8b96c3c3420543b87273e23c37ba264ebaaae0d87b10d365c2c6fa2706d625c7d91efe2c46633c7de410662d193c194fd07ed40fbfbba0527ef8ec54e5c3a655233adc2a7e11f261232df8417be5e72bd8ba7641a7a0a98cfe1164ac80354f761ab80f396db8fbc750c09e2b3f56a1ee598efbd100531f1cc1def24316703ddea2b1f88e72dd58a35310f690787d5243338c5066e5a4af1be2ba6876bc7d62651f57e16be3cccd5fc1dde9bea23dc6d7d2edb2267f256d821ac8adb5f1a698f92fe705036440b869235a4142b19ab758fd9a8dcf566514b9e1a4e5546ece75d152d39f1c1265dd986e068ce7bfa585c9e4736648be64fd8cecf6d55f206bf0e8248dc7d5183b525545e24ecc242b74b99e032eb979e72e886bdcb7283409b3cbaae515c428fd427ce432ae7a0ae40819265583edc68e64c47a06a930a9e028560e19ab3e5da2b7c7b1b2437cf46d9d11fa5285c9d5a919b1a77bd610a1d3f03edf4b5edfdfff5e2ef08492443f1356dc927b5a43ae47dc871330304318c6e39491e715a34fd885cdf214e0cb8b700b5b238a5634b3ee8fdf6a92366c75562d8c9737560bb2f492f649078c8f811b6a3c2ec574b94ea0eee1a71ba31d6a12e51c9862b013aa82d31a4e2a4643ef435a6a288dd2b1c3cc559558da376453333f09d5cbc0f2e7001b1822f4a9264a724e04635ffb83791b4d31735596fcc017d382b9d83bf2096b19c92ca7eb9b93ca2d79f2ae96aa19e39a80e725e5f7deda3000fabf393db1841581f30bad5923fa7e69bda59aa31206607edfecd5647237cc2f7c8cb51f4f1c02e9fee9501bf7326efeca298d536528bb20e16c03cee4e531facb8b736e1b565931d2d5b60920a5fd7ceff28574e7ad9b933ded30517d7e4df04c67f793648e66f63200bf4a5beab92d84974defa93acf6437bc8add04fda53a1e63d9937cdd4494fce31d4805378e147c135ec414c4377c366a8820049231491307704ff1a8eb826e7a60796966c91385999da21b42f3181b12f3a68b227558c2e578406c2d352fd13f6d8d1b159a2f41b29579f597d849b36c41123349f39a0cca3205ca302751e5d8c79b77da4ef6abdacd035c4179f7fc2dd3fd0b4d367f5539917a6914c3f1e47934cd1ab3b02f831ca3d6d2e584280be15f1783466c75ec62de93ed549c3a0e93e57c9fde0c3703e377ecc31b51e0e61dcc0e65044003a3954d7aab8e5e786cc5585adedc346620f2d18e8f1ed9e552d6ded7765e37ccd66dfefb4187198452e8e5761cabfa9ddf6d4b6e3fdf320406e43bdef4decdb158fa3a4a0c46d2008eec1a8baa9de47ac936dbb9f60d9c5d6d6b68de0807b57252583963482ffc6cba2af953d8a2a77ed77e389125233135fe741e87b8df9e400e34884809bb88d5dee6f3efde37de21e35447d953397764fd6a226a8e8dccb356d91a74e65b85cc739c60ce35d6f2d8eeaf1716109a1b686b79c21c71e00ca4aec8f5a40eff219498bf658b31b977e16700808e602225d70cf4949529c4f8c96b368f16f90d8f7a74bc0ae28d5ae3e013830bc7675096fcffbc38b06d94f0e8aad78491aad9fb59c07bdca72a077b46005e172d4fab88a6288a791f4f95f00246d63db9a94016c9b12c2abaa7e14e71cd61b3386845b345bbd5d9d1cb8000c836792bc9aef8ea331e1575c22ffc51f41f33e7c3e3b070852e582c96155847d3e22641089044f857252a89e5e4e8afce7e9973f04e302fc1d9a792d11f7e5d22fa530ccf2237d5f396bc44ec3c7c13f6bf9083c0d27d1cac6b46e1d4d409e5422f6b21b29cbd2e9a5f0902e0fc095e6749566501aa4efcac511a16c87d97478ccded91ec5c6a59216ff99d2ced2b2cb1f51668d7991f53c309d51e03b2aed817f8d0f16c5bddb07e968869e029263eb56e98a1060c12e60d98f5cb277cfdd25ea76f253cfdff3f941b1ff4c72ce9e66ecf2b89e93461898fa119c92b8d215ad0aa4e3c825f9bb225aa5fb17e04e2c382c9e276303e7ccc6c25e6c72061fdf747177097d70ffb5813442491d2f16e0bac5a225caa59c752c95c8314abf6967d91fed7e045ce6f300bb30c7c6baa03c1785e2879361ad3445b51add05624b70e7a58d0817eb65a32f4a07ce4346d1508a4ad39a9ec91145ea28783bcc13de6aaa3d345883ce59121501ed49c4b31194c3084f40f7c65e8582214da043006be2558e2d04f8ceaccf7c7530d619c54122c84834408151aeb4b5f960553b64acd087a643a5c81d1c2ecdb304801091ff83656692dce469d7b92a7df290ff45299363334915643f18a175c3afa1163837f0a154914f50d5419874260cb6417c7125b6eda513497028a9cddc6bdde502a059146fdf2db597912557feb825bdf84b1880bf0db12647c39c1b398eb3b8f3ce88e223d94adc365f0c275bcfc67e62d055a9f9445997a9039dbb44213036a0a941120be760df6a0045c5b9ce6462a8fe9a12ce2b51508a0843b0f13eba4a8cece412bedb8699ad83e3dee6c53a6d93e68ab261b0000a6ed353ec88fd8e9e6f5a892238dfb957e6c00bf343248d24b012b92a37bd7d3300dde6b4f14726ac462ab393698e9b2f03f314448e0c391ab7e30c4ec28e8535092f6953692b26e69a368169ac8a0e654734116592ad9456c7365bbfa17631a080839d14d935a76599cc1713d45aefb70822f44a4fee8d06178fa0696faecc5d753e94fe709f1954b1d974c92730de63137bd59af4b2f272b8cb432a84ca149ca787563cfdf96d53ec090640a0e2e8c8f5140bde25b49404bfea453b8ea30143e8c303e08d9b65f28ca7842655612f4a62f6a471af3dc33b039db58fde34b68e555d69710cc62f4303eced81e6c30560d8b9f28f9544954a1bfb7a4aadf4daf0964cbe71430c00e2755809b5c098323ff5c5ed378834c526c478a26883f25bb8e93e655b9fcb91d4ab49b431e0bc1b7429381d63f0db380355f2dd306a0d4c8eb8030eadddf5a10bd84a2ad86e652f5acc8806874106a333c2378f99b3f317defcbbbbd9889225132eadeb132903a02b49f36953fd54f5a80e9bed94b25d3ae7f22da17e96f34e0a2b91808355beb9b487ee4c27f6e2b17672b1c0ce4b4b48ae3baf36f9d0aec3c3bf3bc0ec78eec361e70438bcbf1ca5896dffb2c3063ef62590ea3ac435ebcbd5ce7b3fe5c43183767230fd513f026c1a6e2d6bb743f4891ad59f17cb2da54293c4e92217dd6380f79b3020fb869e57b2776f286a5264fc602cfa1291d31a7f6ddcd2fb5beba47f77fb4ea82382b86d9eaba7fb4f828c65248705d00a15b1b0eb390fec81f2040bf30ad40da6e07a2df9d263f729ac9fd9b9410dbf36354bcfe38eea50e1606938e237b07d6e2f3092bada688209f044069307c41d30a8d2b65ce98ba5d8ae9c4131c4b31a11ae742b9c53f19686801e50e2130fce610e100eafc8d2f1efc5dad8c4766b0c8a9b411cb8bcf65f4bf13ffa3b8776fa903472b51dcbcd4802e40b5540f2a7314b1a05435ce9d596c67dcb8e036d6db60915dd914eb4e9c9ecec5c2c0c9002557140f327b480df7df02d9d84cc6942ac8f7037d3a45ea8314751a8ce8a3f6816ca972291661be66167c7461f7cf05cfe31c74880720ff50a476;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 32768'hbd1f9229a0818a34ccf9f217a8ef3d10acc7c056b3e944ac89cd526c20157196bf600ad7a081d858a3b9321d0cf6e6d2d25391822a1e2dbd06a51c4fab01d13be77400500604ffd9be0f240f86e9c31097f011796824f83c2eda56e7052f5d1175b0dcbacf7c6776a8692ed575ce20a021e81226234969dc2dd09e99418fe6c6ee0ec6a1fca55794648cb4919142f1f53ca71a811d294835a65f8d220e919387d6e08b2d72274ee9a93c46e13cf3487543e9ad81dac80afe2d624519da8b68daa6ca1c74dc525fce896f618f0edaa0f200eeddb3c8046ddb0453a4fd7316e1ffd5d76959b7130fe5458a7f86369788ba3b4d69f4c722cecbc15a6d5a889e5c3dd0eb500c01f86109453983ebca854c2e9a36fb969f94332a639cc4f61694b60d51575150e434f57eb1a25b373e555f076317be8531d6ef61eeb8f559588abdd6123f3669787b9d4b0f6d3e055983ccc9ce2a663076bb785437e17c2adb33a821b2039a2bf4c530946afbb545f078a5022d1bb455e4dc0f59e4f289bbdc2c56dc0e6c28e403cfecc84aba2b1d9ee171ebe89569d5e1cfc3806b02bf0fdf98fb9fda9177bb0154a3791293e29344efaded52f499beebe568e2798ee6511e35bc7d980c5ad093f453cccc64ae3fa4c9f9e8779cfdf182d6980cef15e257fcd32cd8fd63ff14d718ede1d324ab541e961ff068bcdbfea3eb4eb91b329f213592fbcb692b41d5fea82fd725ac30673641be570b803bf6bded7c08363426c52999ea8ab7229316ebbd4bbfbf836f4b517f76764516185e6e19cbd3788d855520b255cd6f5e2744ea3475db61c22c610a1cb5eb548578d488f464154e1e07e10f65fc769218aaee5ada9286e4dd9f0375be334440fb8605d0dad6a84ffa8ca745d785811533ea60f096d3c5c16323e6f60083103b25ed4c723993b1868029e90def7569e6a49ba48f64082d31cf57c83e90a34d385b1082d96d81b78c3cbd5ba3a6d92ff2289cd3bafb43d7e1943e3b30eaf1f2761a0765943026334a59e8f19482f58f48f197f9e3001c0fa92af69493ebf592297a5a16ac414d8c07a8ae52d3b49d62060d4367d3e74a0be8f0763ae2b6affd7b2d1a4a9249f8fafc7ac400c40faa46588b6428a377d6471cea1dd40209edf64a40c940378325fa3acd84f4237311b314405a4ae17bbb5de31652655111136fbc068d0b13c2c105c4b29094609c1df215557ce9413a3d18c8a9b7ce80001f03e00e01a4f8c0b174147dcac7ee033a9731770c90c18462e56d227037e9f9cb63841215a25d9465eb269e80f4de9d42390cb9c275d72ac99a6f1f31ddc1fdd3bd261ed418fcc43d4715baf1393ca3f6d2af46b869cb6e6af43ca6866664c96a19c6ac218c7b0f3e9efaea8eb089cc88b0ca57ef68313df10b2352b26f17b007e7885bac0f2e50c592ca9481dd906740a412a36891424cc53838277a6f9179ea7ab054d097f11c60cc33a878ca9d36f6cb9ca527e6c2dcceff1e269b69ec344084124b2a6233cad54e476218223d1713be0d3425cc3782c5380201744201093deffbb1b1e0193520bb125e1c67a2b490075c07d96c0e76e1c88ae46f3dad57d8a6ffe1d3f2bfc24ee8651909cefd5a4555e9908e7c328bbdf25dca11bdd82ff2f4c9ef2ab9dfcd8a967a9f8200b9952e6fc8d6fb3bd18657b0b85432790924208a9f52acaf0bdd8a7b001cd5c6e78ea73c3af33fecabf771540c40c8bb19e543f010f02d6704cc4b127cbf0b8e24bdf78e59b7bf4bd9403a6bc9ba7bed3975fb4a428fa934dd2d94d59813843de771ebc1c792d20640fb6cd31b063952070d7c044343239107baa155899e6a9a97c8454eda64be3c7842c4b7c364264d8731aeb0c960162fb176174bd5b55d066c651ce374582ad31b749b6e4be1ce737c51d7691f207cb935ac903298c15ef9b3af6a06817412a6e558481ab609180349de4c42b2984f27a0ac1282c71e0b245210dc2d1d1b78a1075384a488a7b75af1157ad017bfecad7289463bcaf780a5b3ea98fb5c9438d10e269e28aa85e0b59c6bcc1c67d86317ccda72170204724b22947e8e06814324b03d2e5928be63238a0e757939fc6d6768fe24de8ee7dc7827aeb55ed7a6e9a0829e5e92b47666c0af7df7ee8639aa91473e9415b99f2df44935a2d12ea6120fd42096e823729ce74ce9a051fe548eca1340687835adc8cb02b16b0e79f33f86faa4ed6c85193a07bafc883057f1e567fbe39464408a56eb45854b0cda027fd397a4703e4a3badc29690e40b9b8b86df23d3ff688e309b0002978f57066bf9436306134e12e7bd514859eb6a21ee1b255a96b4631b407f4c71e60c04867643cff9df5d74d7322e99d7199fc37d72967544d388b6285e65e7c35c6c5dca253deea0b277ceb860f1809a5b5fb59a96e6c70c1f778b44d0d55ff6b57f8f9ffb95a5e5fe15825b2a77f7cbc1cdf547c118453f8cf31f58f4e3ff04c6ef5494c64300de30082e6c0abf71b018210c22a8ce327fa453414e28001ae91c651b63b862af1b68083d776ae786389d11f44b0e027a59d3cd3696e3063a6ae2bc501d41d4a887022346ba3766e6b16e89c9535241887e53d75c51fdbe5873e3f5ff001c6f4673b6f277e9704c0cf0e2fb1d90683b03012233a16da835994757f4ba6357c39897024dc8de8080ff54db4e51f147767d359da35b0c5dfe78e76ac3e51434854e7aae75f733e3287e3077c72bd57244d8380eebd7e69e56291663989e210791596d427600dd9a3b09feaa85531a0b8131941d7d2a653980d033be3863cfa70f5325ba4371a0ff3eb9eae929477c68c5a101d2c1bbf194133648c9397338c4d3540436900657aba28a4b8a55c220b550b18a9ce7b308b719f6fc43ad97274773145d6dffd6637d6cc5dde59e5a735d771e0e808503dfa77c66242f6c88e3d271e60dce303f311b3762e0628608c1e19b2cc18a7255233a525d0057ca8935855e6f0121ae1009af768630c5cdcb7cc5277225c936d77b536e41aa1822a2c9b2e4a1f829f5be20a20375da44545719029698bf2b0c1b021dbef0b20bf5c38325e368116ee1a196664b111fa93f9d73258477344ceb6f66f1cdc3f73562e0c61d33af60bb40b1f4e064e8bd92d726b0714dfff02504698a23a09caeb43fd7d4e7b160cee742b78bfd34432c4caa87de4ff73622602489f981d55f93f037b3c02b33176ed4a95243aeab3d96817b825a1de666f379ba7a0966b84b37056b1042b2cb66cab49f983c710172b7aa21cf9b7155bbe45a8a47c95c688b3449a115c717b2e446d760f3614a4cb3b9c93e01a36b5466162bc455d9afb6b93bcbc7df254acc284067093f1940b5d7d7d59a0c0d0dd83a5419d14c880caae8f390e15608d97a1da03b97b6061e07a859a5d00ef8f6c7367a5c2fdb63a34f5ffc92ba22d3589103db01e142770354ec87b558962c0617904921c22b5ba9a965a90885f251433dfa56451c8ec3919d30df9d485277e1ca3f45f5d4c9be54380d9c9e76e1c0cced5f7c4e296396c3e143e02744d82cedd127398656ed589779374af95720e8d6c1ff64475922ac74306b5a0b47539b7507c157676f6857a3c0878fe1678b5f71bb3a2283cf01c492cd4cec740f8cbe1861343bb267e8652f45b3eb8ded42f7ab30945ebc8a3abd1a920552f7816c5cf33d51c248412a98a7929324df161959feff21087f29504b2468e7c401d94f77cfcbbd9d90dbac1f912f5b01976b70016ed843e3d333e492b4b8fd8b7c21da1201882a580c03312bb62f8cbba91e21830db77ea1d54a2364e81e50069363f5dc9bd57a42d21eeed84cef6e72b26a23dfbaf28ecd3794b12ad7f1972476ea72636796e71ea58719fa58261a354b4cdab2ffd6f54b50bc6a2013ec4c6a06b0ac20398aa716bbba22b94d79c8cc174dbe79fb2952c04e6694fcef14a291b2c5417a3b4b3422d5ba0dc099289bf797bb351458911c8ce87cd1ff7463ddcf6cbdedf49974838aa8317bd536f39e51349a0f72fa0cc727f7c81da3fe36a01fa86cd1c51a5a497e3a6f5fa16b6dfa2d699e20d3088b16763b1eb5cb15ef830ef92d2b102c8395d0e8a2ee912280b8805aadeb0b21547199d3cd05856a4117d285d955a1b0b3c01947fc63aef6a467a02f1077c09751848efb93599c239e04c6c84441840cfd97d4290d8b70d630fc496daf8bf49d1b53ff3f85a2eff94e99430f431b723cfef9f876ee17cdd41dff2944497b180e8c79c1c62f444ed4b93d9ed26d9d313bb548bef35348289e6fcaf85a0daca62f8ee11f01f5f2cc6603ebd627b3f6acfa1e9834099f4b098e3a90edcccdb641db40e11c9ce2c1866fe1ef4b22c9685a88026a3002c8aad84866e85df79af6cee885effa13a06760a53b52eb0c66b0d598fb149764559ca1b818dbaa8f631042629dffcc45952756492ad0de32bee0f15ae9cb5c836830ceeb71058104d06d7e37f06f8d48183d3d5ab3097f67570ed40bc955e3b96fed6983fe47ede839a0d8a0b4908a7c702de5c54ad3cf61f8cac21fe7495a6a2c7b8ac6b82554842d71af521ce5334c99d5218318bb55235c05a8dcda96387d1e5ba6c61401aeb2a34d8ed3253ffcc6d43e880ac27047afa1ed50da7a2d2b0a8212f455a4b82bfc0d828714dd174bf31716bc835c3a593aac8a06be3521bdb823344df0fbc5f97e1fcc4ba50ead453c65fdc06f3dcd01eff8bc82f85601d037e91eb7bc7f987903fe059e9b89086623ba34dda4476e3bcd73146e84488b9105de30deebf00a53e703fe8e7f1fe22dfa6a24a5fe944b4fa57769c3f7332d7bb85154b8c7dcffe01800b43aff54a061647ccd15eaf6b4d7754cfcdfe36cacc3e73c51c139fe337fb5dfef83146f9b6ba28fac9a07853890b0c6bdc684aea315ec4440e1599b68b69238992be2bd14012e906ca2b5f6643d404f02f2832026051a1109b611ecdc3dde7047242b907756cd77e9df289c9c14dbff1653893efb4cc360e83d852597714ba90b5f4f143d85f760ea3064e90aa1be95a2f6a8ce8b0d2155bf0cc65ef349a239b4acc49ecbb89235144a95074170b194af95543b5ff374d72676c6b30ee7211a78163ec9289101145097d8e484a5cb5471198b69d7ecd0321a3e38b2912eb978e5f35b60dbb9c7f79fb532cbb17bcca47f9610bd6fcb4f050ac5726f076e60a5b9c604e8998bfece596d78b3ef4feb782129397d4a108fda2f64213d6cb1cb6d3e46f1474e79214f6dfd640d6fadba119eb72685353d5c585dcde719aa460b2e5c306c95dd102208b94dccdc938b85b343e13b8821c13bffc83befe7dae180ae7ab4c0ccbfc34bd22b685cb16a45b7d89c68c64f1c2a1a3360953cff97c84eb3d22a1fc52318602bff3c08fddb33da9dc7bc29999296c83f61fe71dd16e750b4413031ee35988e1f17b8a7a8ac95c0cd0ae570b4e52802765e5556ee07302a0db1c41eeb6328c48c72e751d19e1b06254c496a41afd19b4bc2f53589e72dd11dc8100ef82c7b98f2a4b9afa7d4d7ed3f7b89ecd83a3939a1ceb0e1c5e4b306eae47ca5f4283c9290b2620bd730caa6552f875cc052942a5ad3f60ed6c126fe1a759c0df54b7a010c17a672fe97a576bc09438add60f09104d77da5325b4b2dc681248f4678b2d64183c933e549db12fae724fa380b7106555752ce97d56ee98a1303583f070299612d731fdc25e023d4f9aa33d1b49503350ede6e836062e39509df8e77ffd83d7be1882929051e91950aadf0fc88cc11db4bab4d4fe617c9eef;
        #1
        $finish();
    end
endmodule
