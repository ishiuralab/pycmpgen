module testbench();
    reg [10:0] src0;
    reg [10:0] src1;
    reg [10:0] src2;
    reg [10:0] src3;
    reg [10:0] src4;
    reg [10:0] src5;
    reg [10:0] src6;
    reg [10:0] src7;
    reg [10:0] src8;
    reg [10:0] src9;
    reg [10:0] src10;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [14:0] srcsum;
    wire [14:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d698b7e73515db3e038ad94cb33562;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1208ec5ef113f21fe2725f978138afb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16cf2c358a0b9be62f94fa3309861ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec8d95ac8b5c297ef98634e9211d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f85b42bfab22fd6d57967f418a7d11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105023772b036eddb8939798617b66e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56e9b41195446e59d95aaeb48efd4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f71cd60b398242da47d5eb91801fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ff88e2b6d4133eea64e4cb77d226c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a19a31d0ab7bf0a19522bfce94362;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d22e7d4efcf3b6e89ee2425b2d5b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6aef2d07bf67fa704e1bd740e09e96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170d0c3c058c7ff403b98fef6438254;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a6f5eac279bce9ba0e5c9630acdbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1158e13a9d866bb822167861bf651a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2b157a0ecb17f5bd08e53b41e06f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac347f2f17ddc2a8c580f617c37379;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb10fcd8883a50704327053b76244af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1ee03f316510e3c5567c5409a6452;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b4ec01dec585d6ebea18c05ea9eca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbfcbae44d9a9fda041942587456347;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h127c9aa6de03b7f39de5c8bf3c88cc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126af8cf2a7b2ff4ea0965a87528e35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2823915b4297ac2082316f5a4bb8ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a1c1212ecb27aed7e2a491f3f464;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1132e05d20672428dd4f0a46c9090f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90f14277ad05b33b4db78d1f2503b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9b87f715ea6a6e56408bf4bcc10a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ed979d993cc89f1f8e86e83135cd1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113953a2a101fb1038c24741958d96b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha060800a8b7a60ec5f33af2d822d3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115651a74393f4a2ab5358badab00bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c9d815ee3d328199020ec0642a96f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184d47eeaa3f536c9c0e809c68a15f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf955bde80df023f9d56f053f7c0881;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f82613df36fc1dfbd5e45883786ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f0c18389d7a719a2ecad4e3f35a34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152ad8dc44a0a3caf68b3b4b99852f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfabb4190aff2a7ec4fa82fdf919ed5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf971e34220361bc3ace59d0ea931f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h508b68f644c950b0e2ea24c652ca1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1029e55a2239fa27e814e7fe657dbd1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176781af4987f07c3fae414e7e1b734;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60dc97a6c1da62738b2dd86b19a459;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78a75c43b4408c6109d2cd00b1dc9c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121151541ea5170c8478ed928cea086;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2073c23c8a1d358e92d3ef1f52033e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169dafeb163b6cf4fe80c650c4b6cf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f016d72c085079dfada02c81ad30ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acaa861c04ba98f0fca657de52991c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1799d6deab75951abc0926e6abae6a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54b08aff8f9626d0a2d7557fcef78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3fb0aefd4fb76877257ba1cc146cb4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e40c3bee66805777bf8bd1139caad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd805a4ce1d0ce2b16fd99d2b937db3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1790f11c414ff49388dce1929e8668c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb29aa912365a12ec912bdce0fbf86e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1751e74d8259c0e9ab3580aa68c85a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188e5b30001203e9a3130f29418ed13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b0144656e781a1ee06a899a7ff6f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cc0a2f8a3024e979bdf45293367b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7779dda1bc168c7eea5ac04b450f59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf517b3ec5f626dab2ffc989dcbb3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c9a0963567e1e8377f995ae945c3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dfb2f63f8c95f4eef1c0760c15bdf1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c943f0ab67e008f16972edbcc3737b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bb688641438377303be46d1c84ce8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9855c11878ad573b60bf9a2c69581f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d3c5e2624ad76561c13c2a97adc97;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf338390a7e555a51a01c24476fa9a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2743bd0bf83467f4b51ed81e9d755;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c140e1c0ed92a46c213f168ea9f8ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc90a7f2d23ad1133b04bc67027dbc5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16451868294d741409f0c4457f00eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5403fcd1f4ddc0d2fa43b3a73423a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f3f120fa7992466f64022e613fa5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11dc3e02a1e755dae4891e2e55c91f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha202066db546fc3640df2a0c1a5378;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22b665474749edc3aee55b256d4556;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b97f4ac60a073e8641a1ba4ea34d46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a393bd5490b0731dd864ec76ba059d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb35bd9ae8ebcba52fe62571c427dd0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32981b6b7723b095f78e0392dad5d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58b466c510ee8a2f0b0979aefd0655;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31df33ba385d1dcefdfd541603fe04;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c8c35a720ef86336d652708020c83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c88f21158725ff38a86cc78ef48117;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64f565d113278cc542321ff8178a64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6d8b8eaacb5f8b8b7f3f230edd53c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h229fa25d455cef6151eba6fbe268b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39d275ee92dcd2562f7961557216ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79fe3b119eec2fb011b23593bb12b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2231426e63902682848a0a3fcc93e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8dcdbf077cc52ad8ed02ecc28147f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a808d2883cf9b459f37ed0b0b7211;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d7d62cd56d2c5624351aef9091a81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd90091a6a16d38198cc0fd4089d396;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1513e9ac5fe34b8ea56d82d6fd309e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71ce094d051f88f81f5ecdfbee0f48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea82aaa73d071751253a50b9ef07ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34deba05d6303ed9090095d1bed5ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110f6f08673fb10676cf2e71d79c95b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd52df30bc6f73f9318dbf7bece4cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd99e8b043164555350111df800e0b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h38ccd645bc8eb8edc47831100da2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa1715e74d10e787e1859900904004;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7b977a426083bc2a0dd22fb20659c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h551b0b91ca9a839c1eeebcbcde09b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ccc50395cfa256adad991e20c1a63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fa45541481ceb5a345efa2b95da6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14430063af051eb5f43eaff5dc83785;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3c392f285f53a689dd6ddefa64645;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25f8bf52976cfacf09f05113448605;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1caa9f5df08746c33f316abcd50085d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a716ee110a4377e3a6c33746bcb78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189f4dfc581040d64ffe7cdb87fe6c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he55a19bea139d0089d1cd3bc19de40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5be95af61ed2e43c543ad10855f2f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50ff47dad1ebd36226dbf8c9ec4554;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e796865518918cfac16d5ca271150;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155605aee219c6e3788cdff6a6fad3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1dfdbc7b8a7f9f48e8122ad49338d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f96cd3e1a97bae4b28302cc2c69ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88c79aedee30dc757b86abdf25f766;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff63da5c9bf34366bfd7b07daf85dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h502f649fc41391c97f381186d96d59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189f0a81b52821fc83a34a9ba4abeda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h341604ae99248d2220c0a2f85b9b6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2e8941b71292c90070f3a4db4d3e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a009447938c007811cadb295d6a870;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3420c8e0e6a055a91666274c81e1ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a00db5665b7df35196c941e496589;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90a1686af52c8645046068deb61c4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1953f483457084e60da9642345b5ee9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hebb0a4dc53dc801a694be3fc28e1df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163125b994cd0973ad2dd6dce51aea2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9b0e58ded223e4c1ee137b809449d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1559e175a75d70c74e9e34fe432b8d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de92792d31474c48d8c276b66e8f00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2bde1c9cb7675956fc64aa7d8de96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d41220c928ed4ff00093ff1df67154;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eedef5fca4bcb6ba5eeefd65fd4f48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f64a2c2f3aebb03b684655acdad1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182fe4ae1ad8d58160322c8078cd8ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1552708fa34e21f065f27c7e51e8619;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f21ad3978e104922df88c082a3fb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bc01ad58cf13df615433901f74f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1007b2502f978e2003d637b5c0ec2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he804f700ec989e11cecd99c3aea100;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e44ad7de12cb5819d1401fd17e16d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7cc56528b67cef77f01359053b98e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad21f204a19c5e3ff89a80f3bbe531;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b73a05c36250d9e94018adb49c75c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0deacc69366d78529cf60807f9a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e0d4b3e275e61625abfbcbb772ec9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12776ae4e6426b4988cf6c2a11f5522;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66486adc912aecdb9e4ec58ac28a6b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db44599cf0b775075b1b401e7406d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8aa57a849a5fd029773c6f6bc1fae2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd690d6226fd93355cffb65c1ca53e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103401eee28209a57f273ca7972b522;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160d0f3f8fad0a90cdbfe5bd7e606e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19514c1b93f7fb492be978afc4ac591;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43602d63eb1fde48626db8d4007753;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he632b6ddaaa8345167ce83939a8a08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbe05f264fc6a073e8fdccbc9793a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5d5f5bfb2357231a3f3f62057009d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec67321a87f21a4564b15478532654;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4f908288b2af77c47b326d25dbd3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h456c3585e79ca808bed2cfa1ea02e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf81775a10458c7632acf675d1aba1b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a1a046ddbebcd7375efe5ad29cc3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4a3eb8659d7735043eaed03257d8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b3092f7376f27936700b28568c930d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17eee08bddb6a1fb6d6176455eb4354;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1954514ebd609c1a6c09ea35707b767;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3a8d9cea48ac915f0b0c30959f07c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc4e3fba926edb646bf48627aafc1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17864d3746a983b5a38d2e056f76398;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b484a99cc263985293bac84101f044;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f6b508ee7331ffefac37eb80807244;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c801cb9b6d41025df17fa1a85d7768;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe5f6dfb4439aabd1e193c03ef065a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hceb54e2ae22e7a3f92ec021ea77c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1024278afff0f2cfe1e97b4e63584ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acf96d7215fc9c276766e8093e0ef3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb062c67ef39e51fe4f205ebdd794d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19345190be5393ece3829f3ba4eef4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8bd34ced7182ae7cba6b13ed05dcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10bada89698a561c784312cba5a3434;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e3fd762a4e18c2c3c6b03c71894d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b17cfa2e6b7758907148ca34c8e5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b44ef5d8a5ce9e8ab4b19cdcf4b2f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87c549d9397b722342de26abdaf8ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1608b8b1f0286e94e9b514ced41a15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b11c7f406c803118e65d10295c4832;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42d1d70d3d79455275b3a4ccbb958a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc098a0677331f2f2f16e383543646c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ab678a61cf035f57d2b1b3a7271f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha55e702e48715820145ba0a44af1bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc78107a5a0a14970a55dbf4838a87f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120f9d35d08cf4fb8a75c28b1cbe20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90123ea5fa0084923bddf441595513;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df19de43459ea54bb63ded41400629;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h479a87621d47f4e7babe60da5a6e24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1801d743b1c0b35c70ad25a239677dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcf7a19ad62921d9afcde8142ce0b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf9638d5fd11531391809680e20d63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18112ffaba884316125ad03e920e13c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1303139a995415ea1658cc8e8b947ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e4594e16af979147374bb52f6fcff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d8cc396d0ea7db311384a1121dd00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa16578ecf0caaf89458504dc7b542;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1911ad4ed28eee5fa0ada94c82ff0c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fbb0a95e922f27c75a8c2fe0ca5ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9767ac75ca07c85a2caa6a547aec10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b2be7ea0c6c3467bcffc6616c159b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf85c5c62d1990b46aa044821645354;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7bc7fa6cad75389e40eecc780a24e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efe47d3e750e0d9f8b4937d475386;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1537fb718ee2c89aeb61ec94cc8816a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e15340698e468ba7699a8f913495d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h969be4861a200406bfcca1716effc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43eb718c5e761986e81094897d9f45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75e17957ff3c8ebf05645bbf1d25a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11af550dc04f7892287326c82a121bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d7148824a4b86d043aed2dc02aa24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22cbd4c58d087477c9eb39ed4b75bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36a139a2feccc64fbe11247865ceef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139e107e2ccefffa58ff1d90347195d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e2ec3e3a2f8fee0374e29845cb2bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73de2ec3354127cbc7f3c26e05eb55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19341c5d03ee4c120b970dbed1b453d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h607d587f006c69d9cdbe9b1c420ca4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h434733a54d5b53293bda5c541d8310;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82642bdd2231065475e554f5031dfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h948a8bff810683f915b851a39fb424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he121555231daac92a7fe2553ebee14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d23a432cf7e18dbfa4c2f92d4c4e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10be3e79b4722df712283d8426f82e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e851ca566ac87ccc79ef0116fc66af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h101046f5623fa2fd9914542c1002817;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7a511e82fab3ab29384378bf48286;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec610b19d5162baf52853bd8eec41b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2a5dab89d5173334c111a5008c358;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3545b26c17f024ab20575f14a8c55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157df2e53128f1e8fc4ef6045e54bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1feaf473a95b80993e8b27380bb4649;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1639e690fc72e03d0dad3c865896e49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4997889a35f67655ecfe21d7a10e4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12978f0e2af197b780535ee3b5bbed4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h942f5e67937f34cccf72f76426f87c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157caaa6e9b238a6d851cd639da7d80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9696ce506e370cdc4c0450a2b4c519;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc47e54e065d3a793bb2b76ddb179b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he61d26e571b8a158585e09356b31c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a9e0756aaca8e73291fd414b3a5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3c903c3cfe58c8d356d56db24d133;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h356e36e2594189e514b47cf6ae387d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecfadeffb818c52be326ed5a9fb2fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bab6172fbbd5eb4591e6dd27fd6b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a6abe9802deac00b0d4b01106454e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heec7c65797bacd77545b49da78a475;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a7984c8a9452c37a4711ac6926226;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he30c126ca0606dbc5452d91e537d4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c2ae5113832fb206a11b0baa00a22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f2f327c4cf0995ef0283c620ad4f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h932a4e515c692d3e1c6345602c3847;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ebe336dc361fbbb186eb7a7207d95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7f14c624767d6fba00cf734fbd8f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h230b162fde6066a756fcbbcc6cf4f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb417e789e486b91f6796b12bb3ed14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144bed2704bbbca6404d1f35e61d9e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9d81d1f25ae600f7664a56b7e99cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133879340dd285e56089471c9ec10f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10db61656dc2f95cde90199b29a207f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186005eb634e07bb0dfc07618fe4efa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdd32cbac753001f954e50ca9847424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19046167b0e197caf21eb0751031185;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96886b0c43d62f09bdbffaa3b7fa22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161663da7b29a6147348c58d29909bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160a33a75f52ec5114f109461ff93b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11277d34363102376b0bd5623827b44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79fc9a7fa7be9a6e87db342654bc73;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115172ac4fa36118195be9c777c0e5b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hccc34f2ba813ba29e9642a1191e21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e8bd50fb8ae1b1b29e64757c6c45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b435ea9ae8504cff58dd91d33c72e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173e3655e621ca2da3efefdf0272285;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28b1799624cd0931a2c8ad3dbacb41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e856d832de25c561ef946b5422312;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdaa68c2e2f1f3d5d7926936710d1c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he95948172c44770ebbbee22a296d8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18359dfea87a053fcda61a5f427cb17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb95a5bd2667116b627d8bdca2a0240;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1efcfb6eae6518a5c2507407abff6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1372c6feb9c2e3fd8ab8c828bbd29b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h127cbcbfe7d9c13dafc6b6bbb34197;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e81aa558944dc60de2384bcf542a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8e8c130c39e8342d7e6d93e283b5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb33d90889be47ea2801a70b180624;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105d0ab068c9a12373d2aa07131acc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3c1e73fdace807fb032b9160f0829;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce23c084af37ed96ebe98d7ef1c32a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d4edf4ddf0255fc2e7f99a1fa0186;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e6ee20a734a38f0dbc338ef9f50ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f366f8b4410173f9ae04b127f312;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47fdb68525d0466135b21f600bbc59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11bcf16f5138930cdff1698ba1a8a20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe23fb16542deb50176e4132d84520;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h953299bd42e78e0d81ae4836b4e759;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a29dc955be67e54c624152a8b283dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7340f742a782e4b4635abf233c4fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9a9fadf7c9df3ecd9f67eb8942be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7361b75b5322e11093d4c6d69ff0f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8b2f189da70a2a49dd213bb5181ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8af2e7acf84ac2bfb605a13e63eed1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18abaa4cb53ee994aaaea03d7824b96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dcc208076ab65617573c8569cf8283;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba1062f6af3ae3d66abdea79963e0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a87469308fd852c064819fbfb02e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c48c9bbb8a9928fa6f459ea0af038;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a4040cb1354bd0cd161adcdaf9615;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf792b4e5287bee7d51ec6223e0fd47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18820ad5b678e7c5c8f723e964a95ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb359963159fa218de15aa537d7871;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125cbfe7e4d69ef67a28c2a9d693f04;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h484322189474a1ff65d160e3a40f1b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30c6ba57c2fc8f2e838ea93feca6bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd698a666c29ae546cc767f15f1f4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18296bc185dc535bd9165a725c45fcc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5acfd9e30192b94cfbd5739af8f4f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6b907801e1b9604d587686dfad821;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fe64144fa50fba8495d7fd92737fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a745297891eba210afd51b8708f53b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6aea6406d8ba538ed6fb129b6902b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8a36e26cbef8bc5af9532deff07ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8249c368529dad679869916163bd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he60890056294119a1e213c65b85a08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8cf5bbbe10f278578efc4370846d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158156fc9224b8c626cdd209eecd19e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda6421ec1b43eba14eba870d16705b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11093a14c008a68f9e3735baac726d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha13967d5ec9152fdd2386d122a2511;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8889dea4497b6a87f73da6d48c6962;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1611666400e8f7a9ab170f9991fb358;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90334e380208638b82974c4a65a4c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab6382cc093fe5112c0e98bfddb04a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde697e726177d0feabbd758bb39c53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6c7009a89c4e2741271eb65cdd169;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1c2bb36b5156c53c3fc4431ee12bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcdade71cb840a73913cc4286385096;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2fcf81232b205f90b502d9d9f1e5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134b01c037c38905b7d93676f300506;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e29c5b050ae16c7efe1a3f28b816b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ce91c98a9da5de7168d691c1de26d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfa4b866cff0e9a2a757350518534c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd308bd1eae4d9e09a00daed654fa5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16da0837a23fbb6f6716d625ce5c8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1698a312b540fa464cc92dc6ee0d10f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e05afec75bffd2425f323786d3aa41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1958be555805fbe5b8fc080e434218f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107c8ea69f3186d3c400fbfb9c712d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1123f52a65229c0f12fe56b979b9c62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdcbb98415afda710422d5965d76915;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1753ca3f82618b8b2e9dc59520c7f5b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1185f0f300079519da8098df958067d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb2c30216b0f1e30db39e4c84eb9ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2654db28722f06abd76f3c7b89e00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d1af4de434f2a2b98a98db515b1fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1d12539daf3a041bcef126b0a0adf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heabbe9efdf42790f3ee18cb07cc845;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b872a60882c742894f9b32d5a4152a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d983d0158452fd4f16d8c42f8f6d4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2b6f31380b60282891c0d1ce552e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117b5d1fec296f3e74dd546a5934ce8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e40c7c67e2c9defa60a3b35366056;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf2b02e6fce9815c61a5226ffac58b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d889842fd837d6abd918e7f75ba7df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc63e1953336ed524f8fefb9099698f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fbf324e97c6fd4004cd88c6ad237df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb10cfb9544dad5154554aaa2043238;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b5d17a999bb47c5ad2971c624a71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b5b3097604f346049e237b6226f9a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf0b4e7c5d5564c195bc244fef169d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164eba8f799ae25f056cd9493226fcf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h434aa9c4b2288d684ecfb8dd84eaac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52eab142bb3be7002b78b80ea79512;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7dfec734467b5284be27397d2b4759;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd6e8dbb3df081e9a4b78d260ec19a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59c62ed43e9cb5ca393dae752ab29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea5e8c23e682b03222d93b341e5e8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e53ceec31a03819f227014334d568;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5952d882c4db5b88b0611789edc427;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadbe43bc5fa03883464aa097024aa1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31c18a6cf80dff8799d16676dfc3e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde482305c82275ccc67451e4726bbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124c99e4e173495a49f430c9682b3a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce51de83eb733757de56580e72beaf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acfa07e35a79380fde7162bec02d86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd99e3920c17681fb6336341b27ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181f0faa88cf06cbfe312696a8c921b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h172a6cbe93cb9cef9943028d3b411f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h311d88ce043b346a746574a42deeb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13439c455d08f5e3cbac093e2a57495;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6976e2365e81882dd6474957d515e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17133fbb3d87287628894d9ece6b166;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aecc1e22c86810c512ed35d7d19d26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbdd4298e80d1819066161c9615b759;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14520415bba30612636b0d190c3d52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d25bd589407fc9cc206c94b7f1da8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11651d15539b2db436851242cb470c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ddc8c6d3731af34807817c00e443;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he486e0ddc4e676065671aab06ee834;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb37c24ef2524a7914734c7c0360513;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h250df7e81f29c4dc77b9c7cb3300f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f4395c89a05c924dcce9c8fdf0d10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1529f2bcb5e3f483d553e8754725893;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30065cfc4b474d96620d8a6ab5a3ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0e189e5fccd1e357ffc87f1ee5e58;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168668ce0268b17d7aa80d42e43d457;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1257706853ef2197f581936eee0c86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b63687037c6a79875e76fa4709c95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d040c0dcb1c2d021319b3fdb1b823;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0f2a5b6dda48a1e6281920b87b2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1413a110848b5f3e254168bc39e8951;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107d8812c2e5e7218c568f193ddf00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11070e5fb2ddec2102cbb91c1d698ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22c08dae3d987a0c807edba8eebcb5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h137091f04a04a227ff8952276e683de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h999b9a043e5c2f38db924bb9a878e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12530a3fac04058ab5f555d34e265ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f64cfa5eb26b2dda5e5b6579d09033;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ad52f023da3aeefdfec7dc1420745;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcea8dc66e4fb12ce57aefc475a0fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16773ad280e2bd5420e46d107886544;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a3af0b9ba9f2f9f6e0752fdadaf27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c51bbb366c8bd80ade5c1a6cc291c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad13a17901cc3466887fa966d907fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha15c7d01babb0629b4c70846170a36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad1e87e75ac44be35a1ba63f0a904b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c7294ba6f66f989b03d68297b9673;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf214dc130fd2eb5f9255a64b3737f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb1ce2c795db15ff60a741e20d27be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167f20e9922dac3394491634aa79f5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce7e56f8bb62454ae6e1cba16643de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he192f7fff47b83f5de8eb747a0b7e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfde16755cb3747f630d207d2b619b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173a9480e4e55e02a40f2e9fd4d2458;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5140f9d088b5457307bdebdc5acdd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186f8871099b5ff92f158f92e2d0b3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47f1d947e172749c8dfcbbe749515;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e58d752e5230ae4fdb680d170325d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e1317f648e9da5a06c60121196dfe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f49d491c0a4c1e1916dd6c7564a7a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b85509521a1935dc4b0a6eac74420;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183521e588ed35cdabfb15fdaefc1a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1540a7346e732150c9931bcc015b7b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0c9776a8d425a79983565b6cc9f1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b7c329dffc52c02def95af8b0976b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h165dfd03cddb101af63dc8c0c91aa99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1918a18bffcac53270ebb120d5f1fbd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10235173e99d42b892749d5fb0d1e5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36fe57294ad21e10f9c448d20e25d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72ad84499c783463415117e26a223f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha52534023ac126f1c7d4b0dcb945a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3cc6cd8727a8ad2d6df704c6920de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25bf0191bb17adce0abf1bc18c131d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b93c1d5be219d7834a5a88ac09e5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162ea7ef32880eb6b9d0fa51f9ee3b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c1ac6cc5fa0482a131ba6acca513b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1843b71f1951ebb90ff6b022c817325;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f29eeccc10a4dc22bd72bdd6a6559b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11152a4dfea705b500f2682071cd3af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde60d247bbd3550dd854851f99c9f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h221cbab4404d8148c3223b0b6e9d64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h146ffd55a291a23f8e6f13a65a14282;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h177c3bedc5db3b0a6fc52474f934bba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7298ab8a7e355de1905ca99533104;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151199a7c4050819aa3dc3ee2a7a27c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cdf3f09071edfffee77e86a7c73028;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2fe1b31aaeffaf9628e84ebf8d374;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3c0846044268d0f5533f638433dcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e2432e89606c9371abe6cf7578a28;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc22b81573e19cd086415a9084440cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1662247382ca9f4ec0676a9eed20064;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee9a6a6ed613f099f5049f396882bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadb80fcdc1af1e6e69a8ba226ca5b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1afbd9acd9df5a3db0ee4470cbccba0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0f8c7645521826d74ec36ad1b4146;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1712b7caac5aef8fb7968231664c629;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h137a5ada0213054f1325b5b3419dcf6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c02f6c8bde7fc0b92f026a51e1f19;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d793ab8a090a0a9751f360ebbf8ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf43d2ac15d89224732d283495ef941;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f49c431f6e972e748f1ad99445e65b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2818e3a2e8632ad223cbb9842b552;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f13b3c75cf1e4fdc2a36e5d3e4cfe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he03b81174b37c94cc031d2d1efde51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0c59ebd7f982fd7c197855b8ff4c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9756ea6b0be9cf9bb2d84deba09a3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f1bff6ad6cbf290d6bffb70339811;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1493944498423d521a3812b090780f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce0a47f2d8528d708dbf2353b97554;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ecd4fd82054a43d3092343ff8838cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf126f13f3ab23a3a1f1727d1a427;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18202d78dc02dba8bc0dfc63b76c9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1392f01d9badf43ae0338e27c14d263;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c2a776c1746bcb22252c75c5ef869;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8a09855e9b7bf74bb8b645f23c125;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162b631ec3d0a5a317a9ad22ef75dcf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18869a981b02d68c9fcecebaa34ef82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176193558134a75ea37555b279ac166;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb41cd14223dbde4b5d1308888da829;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32e7fe4723a219afffd8ca4e4662b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1c4fe6af7f3a6b35d4b9b8158b58c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcde0d6abff2f4bfdcb08a196b1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d14f043ff20eecedf46052fa6d219;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h836ef9283932635aebf5d5c8722cda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75036e91878e1a6ad8b5dba60a1405;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16bf6269777b006d6978de9ca3d4f29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10344157de015c7982c06d4b7250522;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16aac0624fcfcfbf26d43d7069b2099;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a247ee7fea5750d81a3df0bd1a058;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134b399fec5e8ea00bb66eb4238b3fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a107c9e18edf23d93e3e8a8f68bd9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6f2ef0f5418d8538222277c8bdc41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb76ce5ad43ccebb69447e8697a1982;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdd3a035db1ec7d269979abf884b562;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc35f764ed044a696da15d4dde5aaa4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc90bd72fa029bbcac49aaf5c4e45d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68fa6bc2a405bbe9575594294e98b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9e214fec103f6379cad6eba5819d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a88b09d0153f0b4f09a4aabfa457d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ad734f459f23fae9811c4e12b1694;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27aadd0c1382acf3f4b993a8c29d7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4f8f814c129cb3edef9af3edac105;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdba52b04d963cb0789f142764a7a06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d9057908a22c14d28cc3f15a33ff9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf85fb57fc49d86c389f9cc853a14c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec9ac58c812b3c1064dfb03ecc0245;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d0c5fc148385125156ba74f887341;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd356eca44b0dfbd04fc8af64873d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a61982f3b8edb99abf5d4153cc81de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ce41e6cd7ed571f215cea0de19dba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134c92a741c9e3145ccc7d7fc61b96c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13339461de0ca851041d463e7c128e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117ae5ef7b565416aa5ce397126081a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17430922c37690c5385a07152f34e12;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a39f83dbf45573b9cb8a19a17b2d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h265a8a5a5f1b4d2ac914ecd9bb4fcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd619b70cc3542eac81ac22c87127c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he28ddeaf303e3d3385fb5c4ea8e3e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f767fad2c11bd3ce0a6e88060aa3de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e87ef6838d4c96b9485c3cddf22e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h278f40628a2a9fdfc106c11a71404d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b015a0533708e450d21e5ed3f21ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1743ec3607a46ae52edea9ecf4e093;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bc42271d233550367b57f0323d8f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he46006ab7198b0757dcb8c9d3cddad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2aefa9c1a9c60fb19b83a2f290166;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87eff7a92258e1bfa3858f929c33e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc2cd841afe6199ac8f76973931e1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175161275e0dee21eb01efd44a40c95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h119602d15d87be3231134e36d6a1d95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178252fba0ec867034ebed44746474;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189e2946db9c3e5d7d8275f915f5275;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f342bf23b19341360eb87d9f93b36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef6c6f3dbe3ffbefdc12b236ae3ceb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1201eb465b70f2650027f6a0ecad006;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47c6469c132c8e73b3c220dc3f0af0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h101e00465abc48bb39bd353890b6f81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159524a66ce94d86617ed309bd37974;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h776d8d76c8d15f443e9ee0cb36d187;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120898897a7f09bcac571dadc9c55da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1bdfccd240ccc414108c58c3b10c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa0d1d97200599587b3e66a0ed90ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef62159c11dd25e251def20abf8346;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9ec8e357dc785893b24aead34147a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b4fe8303c595b74d6b0a28975447f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27e5d503c0471acd83d2bf7a420c53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52d1d205de8eeea0103594caf1ec8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd8f2c16842a83066db7456a5b89f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa88d47d3c3884f799d45f50224c2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcece4588b77d34c6b0a302ae125f7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13dfe64a2be8a5651a62c321c98372d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9024eeb4cd9447a18dc146084f27f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec137f4e1baa22c3236be5ee17ec7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h185f00def36b09409432e025fcc8dac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79ff47807ecea25e5ab6e1d63dd71c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d30ae9b85ff9a8c6c85abc4d066f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h566fd6ad89b626060844fef071989c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b1859c121712680fcd9e1a764258;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd23c124237a4002bc38484b7bc6f89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda1b755594c3bf06930cf7eb8043fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h483e0c04beca3e2a528dc6da2e32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ff5b0f6833a3749d2528c3cc7ab54;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfaea2fc10627ab2422acf3c5e036c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92a4f311c0b6306aabb23d2131638f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ba38c49287334f0c85cf396fdfe70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f1e408b37ba3ee4effb0b25baec70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b61471dffe039f08bcc2bd5a3463c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27f8d582b93079ab9fa885a28723b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17edfe7a847f2648be2e0bd5148171d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e8c1004babf3213a739e451dcd355;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d66d93023696b92b11e96d24ea78f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ece747788b72de3b9feb7929d7662;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfefe4fcbd4407562003d914c254af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17014b0ce37a42d2b549a56692dbcfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23b19628025ed33522748af38832fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc7820ef6aa04dc0f1d3fd9c5b7f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e11ad8ac048440ae88321353e98cbd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7a4e0885b4588618910fc50fe8101;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41b4b191d36e68921da22d165fc74d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ce9b3e6d6e4bda8fde68825a85fd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb598b1d45fceb1b4b6bba8b3bce525;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he09303aae57bf2856d6d18d55f34e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a82510be90dd1ea69cb91a75ac66a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f45ae807dd2b2012fdb11b37bbd5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a7ed52c4db6b31e7502edc886e7b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a836caac976bd7c243a7e7e815460;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1764f4c094b134f94b47890c80f87af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18277f3bf553cadac7f90245523850d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae27142be423029205467dd9b85d27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be2fb8df0abb0c8b4b11d62334b098;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2e63f52c165a4a01fac233eef89fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87346e93a21db1b5f3ebf5f987d701;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd66a9142b3d40ba1ad8d593cd6778;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he29c016bc883ee6ceaf28102a2cb8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ea9239755fb0015ac21d2ca676f9a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197c7e8ebbd364f3c7275ec1b40ef5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6714974b6dd4df88b8b84d1c6d69ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a33e84f8616f03fd541f590a0e770;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ed24b83c2b2800b13ceaf15c8f222;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145e4a780a87fcfeac1fb3d4dd80d6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aafcfc9c18e352444a4f4073d2c037;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17343666c9a2472a9a143777e13d3e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd604df8d1f79f41ac4e991987e707;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdea776cd1738a1410eaeb22238a3ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cbe34a842c0bb8a3e0f710241c036;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e490cf9707ce24b437a7518f4169e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8a72481e1d20d1acae1c00e4f96a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2678422b4970094335baa0774683e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147f10c525638ee5a77cd8b4ee60cf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1999093fd7ab9687357698908fc11bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eed2c452ef4a950f1adedb1f458e35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h905518746b6872bc63a05a2e7d5253;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6599f996e8bc7509489ec95cbccbeb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102319918aea0c40069f02099e2e4ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6fad6685f05875cdc460bd5e8c71c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb91a9602463fdee3266dfdf51e6a6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7a0525b2c75c517f0708a1317da7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha48cac36314db785fb3ff08ec6aadd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f6dcc31b265d23b623efea0d83ccf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbf070ca64b908b68ba49ff0489723;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145f0f6e387fa7d65d464a20506094d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bbf3f73cb787756bfc8be3146ace8f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1755532f6bcc8b0438587169f01656d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d3f6845efb4c6bd3d26007322184a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b030d19ec7be5cb8506762475d0786;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109a6f51a4ca8f2cb77b654c417bfcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31b134b957931731efc896a460037c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4722410aa0c305bd8bb60d828a2322;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he640dec3fd085bc41984087d962a31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd284c205ef7fc19cfeb64be55edb1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32ffc475981ba6dba80065b5e07029;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1a364c97ca7696b406f2c239a3236;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9ddc2ac81171bfb4839ee4fe9b0c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90b47ee128da588da7430a168384c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ee2a4b7c4f4bb35700c1893081649;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3362d30736da5674398afbf6d35765;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168381f18e853e4ef083513b5d0b27d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h386c3a9d8665a3cf35172018fde1e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc198146b0370bef055a5456d30b2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd26c50d8ef0f3f07624b2ffd3ff11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd4f0d74b2d887a0c44ec6479242e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d300baedbaa8452955d0a29ac6af2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5dfc814504d1bc01cd8f7b0ba2e9aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a01d7707ac3e141c8fac9dfbbd9d7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h55f55d2081409ad1097ee4f97c908c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c17434dacd85fa321df70ed652a99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51a445dde95c98760e02c6c9868dc9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb0a2858b7c570c2b436fe01debd9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3231230fcdc4083f89431d3c915db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hafe20b364c58b78c0da7c3c72935e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b4095135d179e01ea0530f6f80620;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h873631d542ce5253bdd499f824c07e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h765d52873852c7742b652dff99e2ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hccd32b4ce1d0c4b4cdf85917e30621;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1a4528ce3045c5ba96f2a7550af1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ac8f0370d7236cf25f92e60812ea0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176d622bbb210ea5ec2dd611c01ac71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ebbe3019e6dd406ae40b11002f02c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadf169229bf00f44fdc32af89a91ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be0de1b9867b5cec05075f639657d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5f970779eab6f55e8a9ab278bc940;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12160928c598a7e5c518f7fcb8beaa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc92d5f00c93ca2b1ab8a958436952b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b459ff704d187eaf65a7bf25323eda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196dcc95d95f29a7e77d54005e910ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4e2292dc1983278788b38b4f5eba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15756f244a969cfd8477ee3d01aade6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h933c0b145e61fd965cb993e669e6eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11dea61f668cb195bae64bd5e5771e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0a839128ad58650e25ee54ac2372e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66bb87478f998483503f072de2d7b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123ec01fc3965cf8e9df29d6875115f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6d0999641bdef3a98206d334849e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c506240ce516680f30a96a69971951;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cec081e5ad424515a03791b070a068;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16645a1b5a59e9e98fac7cbf0535c26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce15db91b114e69b8882443702f21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce5c7ea8b14be97d7ffab1463c7b98;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1054440645848a84bfc51fc638992de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha249d504ec684e09a7d4040149f743;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53d46390875e476c080a5f3a028f03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1963f392e70b02d8d512adef3c583ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b71a1c31df5e1f24341b51e478aa4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187946ee043c852d22c760f18542abd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b038ac9638c90b442269beea28c238;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195f43adb3d4c516908ad6682361380;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h398f0e5c6d9edd7dafc104e43a588e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ac9097984760a21a9b67ddebcad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110635e4ab5daa1658a4ab3c6ca680;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5c713e84107bcfebd95755cf55468;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12542af42135bd6648df2e85ed5cf45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159c53fb76ef2df22312775e4f865d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc541e82a0367e76442fa32d8ab6f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144a76a4029de341b0543ec241f35e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b40eca00fe425f53fbac812ad7bd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66e4bfa9db14e174daa08d9c56c211;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ff938a7bca91df7dde324c9f8b937;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b728e6d8e7886eeff3520e5a6170b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15482f15f4e4018431be8a231fdb9b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1833b47c20e493d879f7c26eeef258b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4e30c264dfb05a261643fa3774d42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1406d6cf2505bdd18e3696d3f677c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h329bfb41773f95656906703809b3ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32a55c402590961b388cbd1a1c38e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b60e31741a27107cbab83576d3279;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a534044905d253462be86d3da55428;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b97386218378818215be865597853;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a679319f1345668b8693342d769c6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea8903cda2636f9836b33c4bb6523a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95c7f1906181a6d6cd3abbbb112ad2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17068152cbc47a4113f0d956cb8753e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e09b0e51e943dcc946ac970d5045d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a85632037b247edce6706c00794b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha1b74cb52c2a7db66dd80461a6dba1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1321cf4b8d807d03a3bbc559e38c773;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6e6cbd3a0f0395565febcccc45b5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75783e68db1f348b11b25898ad77ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h858745a5ec6e7cb759bb0d7e74947b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd88eadcda2d1a14c03c1fb3b8da33a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h542286e4e44dd20448ac8a8aba1fa0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b559f7999d473872a8b850d07bada7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5181195e0f52f6b6ee41cd96d2db5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfbc38824158a7a128fe4c0c9938e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h116d01f8b5d30d772b022e60ab86bd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41fca43ddd24e535466de05145130b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c6555d425221277f728af3235dcfe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f851a3dcd8e1b0ab7ef485f2b2a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb0e4d2b00be0ffae908ab378c10bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9fa859594e90aea0510c578e6892;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5000d27567a8519c820e2fc7a02de7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec45a19b0cc9246b120d41f060f04c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3bb27dcd380fbf59759be633881f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcce97ec48640990451192ff6370b5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f498d53e9a33d73206c932af78533e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34c3c003e310783284b4bbc02580dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1251b856200199a99a46d1110221678;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd85bfaafe60cbced985815eccc6b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1570c2c89894d2c5da9f21a49703139;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h798a742e950031735ced09f50b1286;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb09e1e97cb48bd4dbf74d478486b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c81ce2a0e1c845c11def4d899c6770;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd55596135e591c268800a6b58c630d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf83d5a60675ef37c2a1abc45eb1d8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5acd0d6bed4a42c49fa1358128da1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb9fb18c9273ef69fad40c13a56fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7f2cf066e67c3e77d73b89c05e9b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e383ca324573017831061c1bdfc825;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49e1dc35ed7af3cfc77c6760716342;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b7c6aa7420b00b0148a97f027de35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h29cef7cd586fd832a190045e6ee848;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h567ee861025561187e95176ee70b4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197022fa83921a07515cdd94aae24b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180b2207c1747e470dab961fbedcf9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ea4d551929bd24af5b98a1eeb320e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd88c0d9820c2280a2f6a09ff63f1a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cbf63323f2448d1b010082d355119;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f7ecae8fa038053b505597addc71e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd92f09c7769aa653a4c1798b1d2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h273f1305b4e30faeb9531e6d6f5bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79146bbda91b5da548a22f262bb7a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ba95f2118a215c90ff776d96fa8ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168d3fcd8ddeb8b8294e3a198b84289;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8226d6939e7d62512810b2c21a180;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128756fae36dd48c5f565541931fd2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1da8a9e4c90971e8947c2e455354506;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1d39cb5560e0284286be98f58237e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b1c28c446f015c8191b0ddd5c2764;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e6e2431408ff5425223cc777907b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1848f9b1be9a0a37f8c248786d49d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1890707dd605bf45c7082a5d1fc666b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb87a4edcae027608b16c75069e74bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158db5ed104f47dd651940ea175fb17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc4adb11c5864047d5bcbd66d3dcd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd7dc66eab0189acc08c11b212fb71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105cbefb1bf9c217fddc69bf40b09eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32e9486d96f8376c1cbf682f4f45ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d1d624d6a9fe200ce7e68cfcde19c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184530c0fbfc586066f8a19558d9d1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189cba4c6073d8a38dfee6743104b82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a10104b57331859f94503ccb63789;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9ee76c1cd455daf89b1b23fc4a0f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ed9b64f267d430fd32983a3f6f60a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d9aa62fad350c9a12802114ee722;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22365626ee317241ee56e57b949d97;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e081dcd386b6462c367f9b4790cf9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5189e98b74c6a4c92288b8f287fbe5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23e3ee39c6dcb42b7547007b32a585;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c643a9da5410795e293275625cf16b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1296f92045a9e08a58e240fa0d807;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb2bf77d381ddc6c57ddd2d2533a86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7f035c40efbd5ce83a618c74d78f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1529de20f41b0a4d70cadebc56200f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h846f692d759fb5737c96e2986cfea0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6cb59769870624f256599b28a60e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1497e8f6d0ede8316598da8fdf45a67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d6d4d6a6622a571b2cbc2092df875;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149419078aef4917d27d9302738e39f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79c373a0667aca5e4e565124936f6b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d14910a9a255ec76dfe410230dd64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h521de801e693829b07ad537e515212;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195176d6c4a362f469204f3fb195508;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3fdb7bc2fa77fdfbbc282218515e31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0e56b7989ec455341b6744e64117e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e27ce1b0aff2da009f08e1907d69e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb9e5b3af143b00095d58ce7f43c11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf18b1b566bb70ae2ff0914c345fca8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d375c90115a3f9a6692454178dd55a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4eb92c8c0ce7893db09b22425d20aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8acd76254fb0471947df0718bcb920;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45d1f0fba2706b6203bc4991f08d8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105da24b65335cd9134b8a776fd2aa2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb78fc83d08aaaef9e2fceff8cfe847;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191730bf1f49b11f95a96eee6d95e11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e402e28f3c714b378d0fe3bbd0e74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5a39df91cca3d8cfba4a7c9171fb0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8efb32b068e94f1e044af0944507a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd92fb9634fb8da86aa2ead636336a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1a311d2855eab81641cd821eeb358;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1409817e1f00469fb14f3941dd40f96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153bbae3870e0a275bbe51821379ea8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h232244b1703f74313b4527d0192f21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb006aa11758c1a3326456f5ee89e7e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb239b66edef4783961b7efd9efdc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19bc1654fd4d156997e95c6fe47a58b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179403dd1927d7aa01adfb58bd1d0f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1f0390787dce17249d5f2899f5c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8c32170d7f67e3e75faee707817a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h29885836f61a428b7396d7dcdddefc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfb838c5fe84d63289c97e8a6600a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135e4c541c4acfa4bd40083dc8c30b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e106a4b4b04786b155f91ebe8b947;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e917a49b31fb05db7fdf8827bb4c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1bb428a428674e65cfa409aa60944;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he5d8cc1e5f939146c7b1066724d847;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59c9b0287f280ce451cf254d9c583;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c517f7e378702c75168a2ce159401;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19936001af41501d85371272a65d855;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12fd8ed77f3df0afc41aa99e4ad0d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2a6d146375b1aa75e65288997cee3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c5124abc3de786d1125160258c1ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d69c6ad1cd30447a3abff21f6ac98;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b643d045abdfc0df20c3938136de2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a06a48e000f4010787990681fdba4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bd73d8aaf5b6bdd3197a06d9f8000;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ed03c5d06d4e877c56b46e802cf10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b288d1151c508ad98be90d26b52d1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170490e1207cd734ea22dfbde463d19;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148814b9518547a53b7a6e98ea50eac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a11f6f0380070993e913ad0f4b323;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5f2d08be62b0d1118feb6d4d72334;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f3344cfec027e4d09659db469fdb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h644d28243934a5dd6c1c01146019fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe754217d6acfd2e34c7130204c310;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h792e342a55512f2a3383df3defb180;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he67a9dd9309fa97598c7aca87cb68b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf43e741afa95904aae1c9a79c5a9a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e20837c1dc0912c98656d6616aa2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2dad86693c390134fd6f00c06d3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145ce41751ef1b24b3b135140700655;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21efdbdc085dcf02ad8a585621c5c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e835f5a44a7524faf579e5ff5c88c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f968f58a3a29fda9b32b7b80e0386;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c3504e99616278ccc2490f674d785;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134897340b807f194996cd6e1ce1865;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6277a9f4b70b6edbd526bc3c22f94d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89d8c23e2ab6d18a1aac4f47ae561a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1238566caf397f244b2b8812d4b7ab9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c66014e3d977d10ffcc5ba91300a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2f908c71e8aa8d8958ec63740fc38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109c859eed1357d257399ea68b83ab0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1583441aab9682f4ead596ff25ca783;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ea9160a8f633b2eb549f2b7ae5641;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1410d4255127f33c13caaa82989074;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb0305c79eba60ecd54c3a95d40172;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1498488a0de84cec0f2858c48541af5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f1823cfefa72b1aad24f6f64895b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34fffec691aafd2d14025a91f78884;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b30262251bd9c495bc9ae3d641ab8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h429249cedbb470a84fd6aff018c3aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b686866874ea3b155c31d7a3ed20ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2ab127217066c7758d9598e91a17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d534ffb4208224b0f883e36b627e24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd99f93e582b583b6c50a9e555989;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc8c00e40540e0f13c101984acc868;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78efbb1ec994fab6744c15411e86f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee48ba5b00116ba3e2a79695f9a150;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadc5160a0c0e8a9e89ed5b04405487;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0b2769989bbc15c4e44c7f226af87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9ffeac420566356e088a9b090863d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5d540759df2615aba5ce4cd397d91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90b7fc248de23cc5dc93a1bca03ea6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1660d56849bd4bd8fccba2da09b9273;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a47f0f53fc76ffc3415d663f686da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8f800cf127ab3f432da8d6d65767f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12fc05eab1d64ca0e3bad3fb91efa76;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176e5f0d95b93f2d72bf6f462752a59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c74dd35ac82b62d4c145421860cfd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bde7c3ee8ba0efe36b309e084f7484;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h611f23a5a6aa6221fa4eaa1b21ae4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18240843bc226506a492d6921c983eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed391f6067db3bf87a7bd14d81c57c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h933e8f9470abc7ad2a4c5051c7013d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdd4a3824001425d5cc5daa4fd1af42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1a179833b851180aca06e8690d3d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d49d3d0cf696f4b0f1ccec363b825;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a365a710cf882439142470576af89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2f3ba97494e1b1122bbda8774177c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc90d62c19488b79051c2e4c853199d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a385bbffe03d209bac027abd2dae9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7b6a5e1c74012417e2c6f266b95fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1a540523f369a23ba1565547dbfe3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190cc059b5e42620b542ee65cf34740;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7c9b7c9a58fae1e50f8611937e419;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb31c17c6b93a070542bcee044331f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4f5e7d50d2a9067fc38a51b651b4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aae0a0dd28309fefd0e16ea375f519;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c97b71254f0cc77bc7e18f1be38c7c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h825a9832c109497b2132926eb94eb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a51ca207403ef980d275cf72413e80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6d08783f660a9aeed3e7727adc1e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178eb759baa01941fe26ba503be8ce5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18330a8a3092849f03e16c5e3748dc9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111368e1bc3ea47b2c6d5cc50ab88a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109d2aaa1f27e5a395452cb1516a848;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1284c4b702cb5d81b2c4bb7a29eec3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1256e8b70b0f0f6b7d39b35561ac796;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71ce53b878bd8c317af695b5cf6959;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6eafa0d764d188f61a01c1de34e48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103e960e4b6011c5459562b6e5238ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h545ccda482d0136290aa7df96355ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88dcd188818e378719d96bb7d4fd56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3628a56a0ef16d60edde298b4682b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he298bed56d017996a9c2fb77c73519;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c33c7f17959c273c81d66c760b8c13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9b6fb601be0ef6309ffc074db0c0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af4829cb17e94282a874ace14737e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159381e0e8a031c6392085ea77df10b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181881d7f90b4806915b1ce02fb715;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d7cc1fb509e5fd57e9c8c60bf57b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143b860ef2720acdbf34245f19e5f31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41320e1794b548857e552de750aa7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc442c466a71f8973efe8001e48f41c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ef6c054d70e2147f17fd2c8ff1126;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eadcb7fcb1975c7789e8852b038108;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h844484e03e3cf2c4c244f797f573d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ad09c65053924078d33ab3ea53ab7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1955ad17c5e2b67cbefa2e81887efd4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h237fde945b99a3acee85c9065e236b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123c11d2a1503a2d76d875aaf593884;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf8a0874e296dceec808e99e30b384;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1787ec8c031f004aebdc91da8aee48f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9ec99e6f3a01658e640e8f7888576;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df75a86d90615cf11b6fe438f8478e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h841b66edb50c6f8d998f57b92ffe05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13941a537f512fd05ce03c9c3a12eff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e66a9a5b88d1bc66e586b6974a7c51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a79263cdc5a15ffa49e22d48bf06fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf38582fde6e892fdcef6a235cbf343;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h673e1e72a138ab0ae27bcd77dcdd66;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hebc8702c77094749b5cfe8e17ecd53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8eac724e44018db782ae0a5115962;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12aae6ec2fc1429a5e6ed9a57e657e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3df3bd213073e9369f39ff6423e016;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1522d7b0c7407d0eb01a775c293c83c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88d94c31b9b401bb71e25f4658f1f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ae1d216aaa114fc7b0236327f39d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e50c76d3bedc4366f60db6e5edecb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10efefc6ae510864fa23def3b4096bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe6888cb90f48ef788e57e0b1e3305;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcdd7adc438f7123b65d956265b088;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1196d2de67b497cac5035e40a08a0ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h275a2dc41ee7929a39baa308e49dde;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h286440c48bac93242c06d28d1f8f74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2982d49ee351bd7c77ad5370b969;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b3f4aaabed5c8e961997c1f7ca9a45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d16001972b0543e04e22896bc1b3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa482a18e3b2b58c18f552226aaf1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f70a753cb966ddaacc3ec0916cc9b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb04ca0815ac8d7e3a8b07c25d10c45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157a40a52e23d8ac6d9d1883dbaaf9b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2aec880fbb01c7576403932aa56db4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1a480a76be14ea9659609d3ee7027;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6aa323331d57c0098192b9834281f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fb6773ac8ec83d5e8cb0227367f30;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdeb35659aeb98b162b50a86c2916aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1080671a4d5d2428a63d83c748124d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f454dba1e2ddff35679309d6810282;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1818b967e6e8ad8f758bb8585f7fab4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8166b3e6291cf6cb45e2d1142e669;
        #1
        $finish();
    end
endmodule
