module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    compressor_CLA54_12 compressor_CLA54_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA54_12(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [17:0] stage1_0;
   wire [17:0] stage1_1;
   wire [17:0] stage1_2;
   wire [17:0] stage1_3;
   wire [25:0] stage1_4;
   wire [29:0] stage1_5;
   wire [18:0] stage1_6;
   wire [17:0] stage1_7;
   wire [26:0] stage1_8;
   wire [25:0] stage1_9;
   wire [19:0] stage1_10;
   wire [24:0] stage1_11;
   wire [16:0] stage1_12;
   wire [6:0] stage1_13;
   wire [7:0] stage2_0;
   wire [8:0] stage2_1;
   wire [5:0] stage2_2;
   wire [7:0] stage2_3;
   wire [11:0] stage2_4;
   wire [7:0] stage2_5;
   wire [12:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [10:0] stage2_10;
   wire [7:0] stage2_11;
   wire [12:0] stage2_12;
   wire [6:0] stage2_13;
   wire [2:0] stage2_14;
   wire [0:0] stage2_15;
   wire [3:0] stage3_0;
   wire [6:0] stage3_1;
   wire [5:0] stage3_2;
   wire [1:0] stage3_3;
   wire [5:0] stage3_4;
   wire [2:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [1:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc615_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[0]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_1[1]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_1[2]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[3]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc615_5 gpc16 (
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_3[48]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[7],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[8],stage1_5[16],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[6]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[9],stage1_5[17],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[12],stage1_5[20]}
   );
   gpc615_5 gpc29 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_6[48]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[13],stage1_5[21]}
   );
   gpc615_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34]},
      {stage0_6[49]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[14],stage1_5[22]}
   );
   gpc615_5 gpc31 (
      {stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_6[50]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[15],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage0_6[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_6[52]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[17],stage1_5[25]}
   );
   gpc606_5 gpc34 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[8],stage1_8[16],stage1_7[17]}
   );
   gpc2135_5 gpc35 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4]},
      {stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[1],stage1_9[9],stage1_8[17]}
   );
   gpc2135_5 gpc36 (
      {stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[1]},
      {stage0_11[2], stage0_11[3]},
      {stage1_12[1],stage1_11[2],stage1_10[2],stage1_9[10],stage1_8[18]}
   );
   gpc1406_5 gpc37 (
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage0_11[4]},
      {stage1_12[2],stage1_11[3],stage1_10[3],stage1_9[11],stage1_8[19]}
   );
   gpc606_5 gpc38 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[3],stage1_11[4],stage1_10[4],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[4],stage1_11[5],stage1_10[5],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[5],stage1_11[6],stage1_10[6],stage1_9[14],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[12]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[6],stage1_11[7],stage1_10[7],stage1_9[15],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[13]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[7],stage1_11[8],stage1_10[8],stage1_9[16],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[14]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[8],stage1_11[9],stage1_10[9],stage1_9[17],stage1_8[25]}
   );
   gpc615_5 gpc44 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[15]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[9],stage1_11[10],stage1_10[10],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc45 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10]},
      {stage1_13[0],stage1_12[10],stage1_11[11],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc46 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16]},
      {stage1_13[1],stage1_12[11],stage1_11[12],stage1_10[12],stage1_9[20]}
   );
   gpc606_5 gpc47 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage1_13[2],stage1_12[12],stage1_11[13],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc48 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_10[48]},
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28]},
      {stage1_13[3],stage1_12[13],stage1_11[14],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc49 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_10[49]},
      {stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34]},
      {stage1_13[4],stage1_12[14],stage1_11[15],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc50 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[50]},
      {stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage1_13[5],stage1_12[15],stage1_11[16],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc51 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[51]},
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage1_13[6],stage1_12[16],stage1_11[17],stage1_10[17],stage1_9[25]}
   );
   gpc1_1 gpc52 (
      {stage0_0[44]},
      {stage1_0[8]}
   );
   gpc1_1 gpc53 (
      {stage0_0[45]},
      {stage1_0[9]}
   );
   gpc1_1 gpc54 (
      {stage0_0[46]},
      {stage1_0[10]}
   );
   gpc1_1 gpc55 (
      {stage0_0[47]},
      {stage1_0[11]}
   );
   gpc1_1 gpc56 (
      {stage0_0[48]},
      {stage1_0[12]}
   );
   gpc1_1 gpc57 (
      {stage0_0[49]},
      {stage1_0[13]}
   );
   gpc1_1 gpc58 (
      {stage0_0[50]},
      {stage1_0[14]}
   );
   gpc1_1 gpc59 (
      {stage0_0[51]},
      {stage1_0[15]}
   );
   gpc1_1 gpc60 (
      {stage0_0[52]},
      {stage1_0[16]}
   );
   gpc1_1 gpc61 (
      {stage0_0[53]},
      {stage1_0[17]}
   );
   gpc1_1 gpc62 (
      {stage0_1[52]},
      {stage1_1[16]}
   );
   gpc1_1 gpc63 (
      {stage0_1[53]},
      {stage1_1[17]}
   );
   gpc1_1 gpc64 (
      {stage0_2[53]},
      {stage1_2[17]}
   );
   gpc1_1 gpc65 (
      {stage0_5[50]},
      {stage1_5[26]}
   );
   gpc1_1 gpc66 (
      {stage0_5[51]},
      {stage1_5[27]}
   );
   gpc1_1 gpc67 (
      {stage0_5[52]},
      {stage1_5[28]}
   );
   gpc1_1 gpc68 (
      {stage0_5[53]},
      {stage1_5[29]}
   );
   gpc1_1 gpc69 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc70 (
      {stage0_10[52]},
      {stage1_10[18]}
   );
   gpc1_1 gpc71 (
      {stage0_10[53]},
      {stage1_10[19]}
   );
   gpc1_1 gpc72 (
      {stage0_11[47]},
      {stage1_11[18]}
   );
   gpc1_1 gpc73 (
      {stage0_11[48]},
      {stage1_11[19]}
   );
   gpc1_1 gpc74 (
      {stage0_11[49]},
      {stage1_11[20]}
   );
   gpc1_1 gpc75 (
      {stage0_11[50]},
      {stage1_11[21]}
   );
   gpc1_1 gpc76 (
      {stage0_11[51]},
      {stage1_11[22]}
   );
   gpc1_1 gpc77 (
      {stage0_11[52]},
      {stage1_11[23]}
   );
   gpc1_1 gpc78 (
      {stage0_11[53]},
      {stage1_11[24]}
   );
   gpc2135_5 gpc79 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc80 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc81 (
      {stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[2]},
      {stage1_3[4]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc82 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7]},
      {stage1_3[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc83 (
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc84 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc85 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc86 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc1163_5 gpc87 (
      {stage1_4[20], stage1_4[21], stage1_4[22]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8]}
   );
   gpc606_5 gpc88 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[6],stage2_5[6]}
   );
   gpc606_5 gpc89 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[7],stage2_5[7]}
   );
   gpc606_5 gpc90 (
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[8]}
   );
   gpc615_5 gpc91 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc92 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[10]}
   );
   gpc1163_5 gpc93 (
      {stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc94 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc95 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[5],stage2_9[7]}
   );
   gpc606_5 gpc96 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[6],stage2_9[8]}
   );
   gpc606_5 gpc97 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[7],stage2_9[9]}
   );
   gpc606_5 gpc98 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc99 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc100 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[2],stage2_13[5],stage2_12[7],stage2_11[7]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc104 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc105 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc106 (
      {stage1_1[12]},
      {stage2_1[3]}
   );
   gpc1_1 gpc107 (
      {stage1_1[13]},
      {stage2_1[4]}
   );
   gpc1_1 gpc108 (
      {stage1_1[14]},
      {stage2_1[5]}
   );
   gpc1_1 gpc109 (
      {stage1_1[15]},
      {stage2_1[6]}
   );
   gpc1_1 gpc110 (
      {stage1_1[16]},
      {stage2_1[7]}
   );
   gpc1_1 gpc111 (
      {stage1_1[17]},
      {stage2_1[8]}
   );
   gpc1_1 gpc112 (
      {stage1_4[23]},
      {stage2_4[9]}
   );
   gpc1_1 gpc113 (
      {stage1_4[24]},
      {stage2_4[10]}
   );
   gpc1_1 gpc114 (
      {stage1_4[25]},
      {stage2_4[11]}
   );
   gpc1_1 gpc115 (
      {stage1_6[17]},
      {stage2_6[11]}
   );
   gpc1_1 gpc116 (
      {stage1_6[18]},
      {stage2_6[12]}
   );
   gpc1_1 gpc117 (
      {stage1_7[15]},
      {stage2_7[8]}
   );
   gpc1_1 gpc118 (
      {stage1_7[16]},
      {stage2_7[9]}
   );
   gpc1_1 gpc119 (
      {stage1_7[17]},
      {stage2_7[10]}
   );
   gpc1_1 gpc120 (
      {stage1_9[24]},
      {stage2_9[10]}
   );
   gpc1_1 gpc121 (
      {stage1_9[25]},
      {stage2_9[11]}
   );
   gpc1_1 gpc122 (
      {stage1_10[19]},
      {stage2_10[10]}
   );
   gpc1_1 gpc123 (
      {stage1_12[12]},
      {stage2_12[8]}
   );
   gpc1_1 gpc124 (
      {stage1_12[13]},
      {stage2_12[9]}
   );
   gpc1_1 gpc125 (
      {stage1_12[14]},
      {stage2_12[10]}
   );
   gpc1_1 gpc126 (
      {stage1_12[15]},
      {stage2_12[11]}
   );
   gpc1_1 gpc127 (
      {stage1_12[16]},
      {stage2_12[12]}
   );
   gpc1_1 gpc128 (
      {stage1_13[6]},
      {stage2_13[6]}
   );
   gpc2135_5 gpc129 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc130 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc131 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2]}
   );
   gpc615_5 gpc132 (
      {stage2_4[5], stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[3]}
   );
   gpc615_5 gpc133 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc134 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc135 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc615_5 gpc136 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc137 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[2],stage3_11[4]}
   );
   gpc1325_5 gpc138 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_13[6], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[3]}
   );
   gpc1_1 gpc139 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc140 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc141 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc142 (
      {stage2_1[3]},
      {stage3_1[1]}
   );
   gpc1_1 gpc143 (
      {stage2_1[4]},
      {stage3_1[2]}
   );
   gpc1_1 gpc144 (
      {stage2_1[5]},
      {stage3_1[3]}
   );
   gpc1_1 gpc145 (
      {stage2_1[6]},
      {stage3_1[4]}
   );
   gpc1_1 gpc146 (
      {stage2_1[7]},
      {stage3_1[5]}
   );
   gpc1_1 gpc147 (
      {stage2_1[8]},
      {stage3_1[6]}
   );
   gpc1_1 gpc148 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc149 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc150 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc151 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc152 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc153 (
      {stage2_4[10]},
      {stage3_4[4]}
   );
   gpc1_1 gpc154 (
      {stage2_4[11]},
      {stage3_4[5]}
   );
   gpc1_1 gpc155 (
      {stage2_6[12]},
      {stage3_6[3]}
   );
   gpc1_1 gpc156 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc157 (
      {stage2_11[7]},
      {stage3_11[5]}
   );
   gpc1_1 gpc158 (
      {stage2_12[11]},
      {stage3_12[4]}
   );
   gpc1_1 gpc159 (
      {stage2_12[12]},
      {stage3_12[5]}
   );
   gpc1163_5 gpc160 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc161 (
      {stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc162 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc163 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc164 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc165 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc166 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc167 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc168 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc169 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor_CLA54_12 compressor_CLA54_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he5ac046fdada0b714487f136e0ca08fe0d50bdb17b3c50eb2bed5f54f0579ecc1cb7165f88f4f6cdc32bf3de9e16a9b17716b4c083f572e3405376cbdbf4a1cff6ea932b58ae3baad3d146943931186f4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3bd6faa9dcda74603fa0f06d89ab5f187e005c442b826ebb1894236012ced596dbd0a28402d1061b8cfe5ffe6266217fab908c768128ec9a8f4df07290e4fbeaa9f0bbb3242bb8c18a931de04a5ed2df8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h2d07e69c23f2e6140ebe27501c3e0cf8cf20b81fdbf930ddf053e881084cb6b83bb8ff01f28175657b591627f18054c9c3f4cadf5ef7e9a67ff8c429e7c27ef74d3d62dfe7f5b87dc49716e326fdd1dfd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8bb48c58339ca79ac70d6dea20e94e5c992ac307dabf4a108e5622a1d4f0147d5d6477d18cababa5292d9f62d16a1281e6823a815e6938d56a2a76a7318042bc25cc33452e3e49a6c30b86008b8b2b7577;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h58e42790e717a07520538b6880762d9c769416eaa21869eb1c2ef4a954481a8caf0a8376d44e29a88d1518773fde63ff4339b3766893ff79eab2902a4aee4a39422a702663ed0668bdf75258898fea86c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h420d106cce2643b6a2f2a79c27ec2f7f6ff2f7693ab1bb5e8a80d5540512f191758fc9cc56d02bf0a54d0f3c3122d1620d41186adcc9ab49ac41cc81381ff7c308f349441910a9a0e9717060d49b30c990;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb6c4cf9708561017bc2b37d8b624219bc872a6f08ae6a9054460e85af52efec5248b61f59f0b7cf4bdb7edf5810bb0724c3d09bcf6d182901d64f9a33791fed0ccdd18e43e5cfc3065aab30e6b5084b58a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hca7dcb476a6c281923d4dbe5b0834889ac683f8c9a9bb318b508be151ad63c96c2b596dbc6041cb33f5529a1e4d20cf63442cbe63618594496ad2908d7319c6310b85864cbd5e0a962c55bba8f8a1829da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf6ed5bfc64230dbbec875515e9fdfb8c91f38bc19e8280aecd62b4a0b5dfb0c30e849d456950b64b5a28c6ef1fdb993baa121f68982c5707b59b4fb7ca490421c67a4be54d14750e586dd97cc1537f795b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7de66fbdc5f01bc5c3951d926e8f2e69a64bf4b37e8d19bc29fa64bd310527c9f938862539eaf67ab0cdf9b4411bb85932b4e2f20efe147fda2ecff86cf01c8264902eb886f51e445528cbe8ef78ef51fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hefb62e551de3e28aee6c5f09be643098d4db90c0e7b17446554c11b1a6d694580e6600538a7f3f6d3fb3148a7aa1a8339add7326fa6b088ab153c9ce65b4daf38408a582a7db951dd6a0c247ff646ed947;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6ba2e108610ebb8616bf223849425c93f6f89b0d5b7f8a9bf99b9fc7192f6c6841c21059de47ea7a25484488baadbc098f3663855f09cfe4d99fd75845c6f4aed50aab2338d01b28309872ae63a82e76ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7fc50badb8e83c2c199ad8bd41304f5ad78cdc1cf38de1f4d8c440945bdffda82519b068275e40035798e3b79b3485964639bfc87652d589d8e9587d95774661dbf643288ef4ce5e1d1041e367070f3b92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h50780953ca4396415a0ee78cdd49d11e21261f7a67d59c7c10dba41defbb2590e9279cd6b0ab328a0c099888e3eff90ec19e149a4d33563fe366552aa36030a3f5578db540902e5d9d67888a966e708423;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h97e535f0815b818d6d157d980954ef02765b09da8503f8757c879bf32d418f93403d49cbdb3361dc86275218e86f5012709454f9d3fa19651f1f5768f55d0c707b26fee645d6b2e03abce9914d11ea488b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf862dc23a71ed4d0a024259a2dec79b4b9b0ab6333dc5b35c474feab05c885d20ebb10f4a70aba7eadf29df0dd4b40f7d99fda01327dcef75095e8eac1ec3fa697c2758ccead5198b5a08f2b1da3565f8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb5f1cbd8cd2233ee58be0d5c39ff54c830c8c70bf17f2f8b634ac9a02bc7dab1bfa01b2dc40ce3cef32fcc5a23f2a60cc13619f6aa1581a39e8499ea265734cbb5d5ff98be5af79bdf927f613b5b28e2f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb3c825cba4833b5bbc7af32611c577dead3cfb7cb55bd3209584df1900c6ebfaadd150ac123d36756d55b43493722311f4f45cb07d135b453eaf025d26fca40377a0c631b96d6d26a010fdbb5c4e91e506;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9ac53936b3bf73abc19d8b080b060cfa694ccb343144740724dd0b34e204ae3e3ad3c032764ac21d04f1f0cfbb250cc3049294dec1b38cbaf5e65b431bca715499af241722a3c893b41233a3d18dd61b8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h62597a4aedee4bb78a7fdd139eb6418b7af86240d81b2bc413ba2efe58b8eec245b53b6035ad9c84402e6ae67e1f03c13c3dd74b4e635ff0c137e0d065cbceeca5f4f4a4601ae1890b1cfdd6bf6cbbe4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he9b8e5ec19e84ffabfaad58804aa8e703900b4ce9c4478f1f5a137fdc730d231bb23e942141ba2e45376459cc27e0ef4bc4542c50a88f4aa1738c50dd02566d180b7485175f0dc35786238f6a2950d16e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h53354b4d884a2e2cace0b1eca3854f371075b3fff85d7fadadd6b6afec2be6916e8afbe2b7c3f34e24df9b0654e8baa0df32f544afa0b8a8dd6c5a38d40922d38707bfdf342495f9e7594a2582f0126654;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb7e49afc8e93d34fc4793c9be72bde1cd7549ebde792cf5a798e2c5d28d43c9d08e50323e5c5b9dac67e1b6490ddeeca6ec9c181b913b0a05f3bd41c5efd32c41d71d2e27d6f5a001e1791d491eeb39e20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8501f3ada4de41bca9eafbd397516aabfc970ed2f12eac84377fa9674401c91522002124f8e0c4492a313ac7c8277a81f2ebb2fbf4d7cdb74307ed74248c839cf5dae4bccb54b0ab81a524bf793d321739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdf5ea704fd04298ba5f82445b7bcc38784ca6f3ca4e3e742b049863b497117d339e5e8ae0430a977ea37d9229a8635cbe15a7d063055b70e734de5ee320925de3bab10d678d6472d6cd6c98ec88f907197;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h67cd62142098c0cb06bd54cc8859051cf37877cbfce062db2e781875d31d76418d071cef18214e76446d290b0af0f8f4bfe04264ca1df950ef56023b5bdacb71630083919624d4436903cd412614522b62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb8a7fcec696e293b60294613a27699d1737cd2127602e8ecfcdde006a01bfcd07a0366f2d97275e6fedf5644eda7c30d0dfb397ec7c52e69d43b4f40d557570e0466e3e4324499627654ba6af9ef04c2b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdaf2393c549d0badf270e23b82625fba1b95c0fb0f21c277ff7397faa185d7c1f18130a397123cd7c44ac48a3a3d0f373f3fdd8c3da6d1fc2870ecc42f878928ce426943133ba460a3f9c121a1c7c1f8a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hede0003239cab6cc43b3d21787d7ce79221ac6cc0d5bc68494af397336840e5e115fdeab9fda7c57e918c79323475c009561db3f34be54e4f0a02ed1fd5cac67952b0c59ee0fd439794dc68be5e5fbe4eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7779c1504536a7fe4c363aec63f7365907f3419cea082fdcb7b65ce2525f8bc5f0c974b44e6ecabe42fd6391be753f7b4ebaa3cf415c5f53e12fc8489162783ab38d1b55b723bc9178a68ff6c56788df17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h72895d569b3fabc64b240b183a81914f404550f9c08adcf30a8d90ff200d7ed61721fb97c0d1f4e526e8291da27ac64e3ba336a3d4a25a1eee00837ecc54539b92a98451571f6a04d5cef06a1ecedbb475;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6d6c592249fbfd31e7caee7ce5ab6ae7afb610a2b59bbd7e42f9ac19c4f5335b4f379902593b3a44fcc52d5446859c3504094988c8f6e4afa6b84ddd8f01e3bd40a13f4d069f058d73b55106f44f3f32df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5b953cf3694c1699bdd0a30fcdbc3ce6e0240cdf352e2b1791c632cdccb22322934d7b5d125c2e946a714fe966e8fee800efd9fb546a63a345df79dc40c0adb894c23bd15b2c38866e7325f588da66c5a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'haab6714f2f36ec6a464716ef03e132eea83a42432b6377ed2dad7d86254e1fa836d3149e10bae0b2141cc4421452fea013a63f2478645b72cfdbd1617f43421a915049cf15c9b92ef9680f12e7d98469cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9e7d4dfdd0f1947679fcbed7abfb6b1a3b2e2af6e85ebaefd8f52080ddc382ae35b16e3b72473366122536e6c4fb04601448c32c179ef0abfbf846f99dca0743437fd0e1a326876854f40cfd481643a758;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h93e34efdfe2080b34703dd94590ce5687d5543fb21b64d2bdf34dde146e01e4f9a27024b972b8b1457bbab74c806a72fe2a47424e09f25dc3b795836c2328c9f5c77d4abe5872c10c5edcd0be950b3a0aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1815dc4b8ef10a086fe6ec34d858004033571a49c73789b2f1c5b3dfc77df57ed304f44de3870e5efd9ac7c3c86fc4f9bd4567b6c22f73bbe8fd84d85aa36084cd6cd0a25798f371d4605e0ea5d59efeaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h56dc319e9afbf17b4fbcbe4c199fb23b1f634616501c5fd914fd193e45102aa4f1b1b659e36e3ec1a0caead6edda27b0afed98f8ac459975630d10764941006b5dc7726c8587f9e3ac66d8d19ee0e089d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h44bccafc007ad728fd55e8fc99404838380825980a5342e65db0e48ac946f7cd8e8d2d486c07d9256c4b3dcc305a41a0677c53fb8b19a37dcc1acf36785a28892b91e0b7fbfe3b0826acde8ea738a47dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h908975caf742784a99b2de1660f5e884ad4f36c46ae6bf7dc3572ce89279b5e62646eaf506c9cf9a5a1c4196960ff5e2be3988416676e5e3ba1a9586db0a029f2331bdffa871175eb452f0ea4f1bc723ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h651df737f0e2eef505cf0336f6794bab9ef14ffd97c82688402af6bc131eaf326e793f2f45299c1fd9df28efe1254b54ea78ed714f5704e929e638f8fb86483c2cc800bfe8dda2609e552f10bfa9a76cd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4b0190e32f3d12f8e508a95021951569cf625e72db5899897cf210c566e0510c85bd015d07079b6e2986b6849477e1ab6154007361eb82dd7baa7045b23349ead8a01cfe579280a66d2eeef1c96979d7d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hef9f1773aef79eaddefad25426f11fcf9a5a71a2363b060fd0bde2bfe13b141d65665b3ba9368bd9854eca4ed41e44dda9c7b4ab7c8ab9f72806dbfab0ba35a968a3addca1d74bdfb8ab218201468220b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbd31841b95ac8b4a0a04f4a163810fd7fa709b492a1e05124cb074d65775b7f53cfbd83aa6f1ef05d5499ff3a47f977e5380bed5cbada501b8c8d46977a094ab3c1e95f60c584a92f0f1b623e6c26c7ceb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7e590f7ec25c7284d478255ec67744eb0ad7de6078e05302d998858ac3a231ad8c708400de82c16ea0bf576fe18da5dd598750b7d1a037bbc1ce9cd7675610e876c933f8a1a8a633ce3abaf4c73cc31193;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3ff0ba9d5effd555cad6c72607174117796fa5f1717026d135c956b3a01bf6cb2b426ac536bf6a0b3c7de9af2c6475625c2937f9fd01688b27029aaae3cc66725e77e52a3cd47943fc03327a9a1251ac1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9b1f45d6f4204a136e93253a8822d2893f5e13a8d18e08a17b136c68b248880a759da0ce8819f0ee20cb78225f0393b2ce25ff4ba112d109638ca91db5865c0dabd04c25ec511de8dcf0ae95b7366c990a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd101ac5919f645f1339dd3690ff63cd0b5ce9df87533012fe9c9c10ddcbccd3af5df9badd50d3186be72e31f04bf7c4f3e4747e3b854bf852e5e8226afb9d80fd30fd1e27806a1e270aebf48977d3a74c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h285f33b8845dcb0e7934b0502f8b2859385889ac87c00fd29a4cffda7dcc84a1fa568d5f5a08b77f8a1b54c725a4c429782636bf9cfcb7dbceec8f855a7ba99178cb107431c8cc9ed5c4b407dea5953f39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7cb5a22bea801461e3d1cf884b6c979c91a580f9c450f719768d9bc6a2810874503d502ccbcae1f381197918968513671949ed556d43ecc0af0f1a0f3b87223218fe997188f291539bb87c9c9e9a1ca5ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1f4ca13483bc1e35470f1b446f93c36eb55d38bdc8e1221f372b469abe9ce0b212870e1d93b9602a6efdae2d5f72c4927b2e1ba51bbfdbad31d650779a97b1f27cfd8e263e78afa320bc46308c03384b06;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3e1cd37310fb4e59ad124133ba8989e5fcc7fedcd212c3761c649693644a9f8cac8402cf78851b55689a0a0d5b4be6fde4f6b3a7ab2311cce91e49037748b7797ea4ac0d318d5cfb49e97aadc88177d3dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h731a191e1ed5ad88c8ae35355d74624bf8cc202eb5f7ca7947cddfb36b882014697ee7006640fa88408ad4fc3941862ecf425771cb0262eabdbf3010f90e5a1b03d5d4dde3c0f6598d49b85748cb4b100f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h78468066333464821b054bd2009ba55d3420ec3d9465a17dbb59eebcc11d77ad994407d94ae7f27e8b7aea4b3e8c82fc51e70bc1b77de7bb5ef8d0a3f1fcd71d458a4ffbb1fb1c15aa2f8fc85d50c42fdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hed7f063b9084866f030e4acbbc88a5a4941d723b38d4c3982b0ef6eeb025745e3052e3565a14c865465bf662d8eb0552dba5f0a790b38db2e8103c45917620ca832255824643d9f22e276832a87588b3ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb4c5d1857b03e4968732cc864dae4e03c426fd1e2272b779145fc4b5136bf401060b868598a96045bfcc0676d165eb17361c444b8fd925c6787ce0d7a9bc9743e4fab481f37246c110f1b5dab14add1865;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha0007f556587ccc4819ff66339deb0e830e14aaa2bb68f851ddebce01fc2ce539f92b90c44a243e913dfd0067834f216834889e460501507fccff37095094fdc3038341294c2d1830c895e5bcd2a2193ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h797afcb14b8bac3cf57a31059bb183df0128c98a77f7b5becd61440cfb109aabd716f503828a2a1ad5d20618feabcba41038b288037fb85ce8387110d9fedcbd6c7ca2d433689f559534bb9aaeba40d2d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc83ffe4159616f5ced743f221a3eaf47ffe7d7fb56965b07b454d4ec631493c04003f64d5d656877ac8acab4cf1bdabd11091f2351e8f440b4dfde608cd69df24058d28f1a20d7764cd618c74f494c03bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5c6366061615ffdd627cfe34f186c9226d0ff1eaa883a30894023e0c79b08014888320fd6e245f747a916aa1bc175fba953198610cc52053c8d2937d479d3c246ffcce01839e86750d34c8833e48f0a45c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha1228041292b202eb44f255ee746e22cc12fc04a341788869653365ea48f71bccf716d03767b610551d4d69c3249694573164f2aefa8a5e13475f9c10370e24e9fd44c668cb15a9ab739af922dbfaf1b8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5d0a4e61454fcfd5dc9b90724dfbb430344a253c60e06e1dded51eff6779fe837ce40bb0040da419031990c533b7a6e1715a528343165decfabcf73b7c7b26fc1bc333a7eff3e84a02840b2e78d05fafa5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd35698f61a3ae915e1c0a95da54e91ad2e69bcb2896d7d5fe28764e1e67ba35891d03661e4f55a9b01e670ac36f0856ec2fe425699f2f2143b98dff527018ee292cd7eba7e6a7f3a9c6c72245f7328a24e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h44e483507ad5736257b78212439b5bb6bf209df6d15e471426855b4a24db5ebf396ae011b89541b97dac8b24ee0329e844675ec1d24a36c2e45dbf5e0907e277daf788ddeec827481d8a943c9ed3051c9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcec19d09eb58ce1794aae2a9aada2105feacb409c21996522719ffaee4b0885df2e47d10f7b2a0610d0764f61ebd7e340250af3b84101ab2f8ad2fd937084f1a6e4166dbf55f81b54fc51036fd990405e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he8906f640424f774b0346aa673ec6c85f6778500e14b7c59a42347e43fb0d473d9fce7c33dfe6a50a6375b38858daec34159e10b2afe5c906956e03d42e78ba68a64d3a59204cba0c40cfb21b26ffa869c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd97fe7a2df9bd934f8b877d50d1f0656a0a1b9f9e678ac32f4311d94c89128a447115c40a792504d3716fdc3827db1f1f4824b2bd40d1b180eed619edc8d6067c499f7d652a782947c2b0467c090dcdd48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he885b8f6e685929945c24f4295de4644c76ddf190ef8380d09c02de185d96b51490c72b1e0a050829edfb46048f632c090d7e37c06e2fb6e2b414a858f3c89ac2716124492fa42654c6eb15cdac6abce6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h406ff3e4f215c60c4eaea5bb823cb6bf24888f99ff8bd07a078476bed7382e3fce1804718db808f5d41bb922374dfd19e70e14b95c18d86cb5248007cc2f10b3df24566b384116cd2b3d1fddac0768dde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h190c923fa98cada47651bb368b3090ab8d30d91be574eed11de9db8e4b0927b154fa903b220c1513d00e0c623f764fe101ae78d941618c56dfdfe295eb9a0762fab83883430ee7aa1665291033f3dea174;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h600e3e5eb6e5163c411d4dedae97801d1dcd5c7141cd7ad8b859c960debfd7e33090bad90705d9bd7f0f09ffe07edd9f057c8fbf5b027a6fee823809b82251bd16976523997cc68230cb8fea272d70acbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9787e0d773cae4aa06337894ab287a012fb06079958df2371614a4416143f6780fe934d706591e2f18f6a0c2ccebef4c8ea2749bbdcd472a73508e26f2066b476039c6855aa99fec3b43e2e01b3e2eddc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf68af0c0dfd5cdcef47867362001139886dc2031112a30e178f32f3fe519e7630e90d7b6eedff4864c5a109e092e7068a8119db4bb347f4b08c7abbf0b80685ba986a5e349e68ce023fcc613f88ac968d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h78cba4bebd26913ae2d78ccb8f8c5d0634114cb39f39486ae6944bfbe994dab7af1ddd8a059ebf94b83f3fb943a1b71b2d9e134024574086b55fa4b871d9528afad12d9cc1311e3baa71202d691d018fa7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h223603e212bbb56e4b455b89b10b142584689a7635dc8a295788a0e53f192d9b673babb0341b45434b69ecab669e5c9c9b4582f8c1a8852bac757dd44788b6ae028857f942979d92980752d8026d73140f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha537435af858d55671396d47992aea903c94ab14ae1332184fd0d62eb8baccb30a33683e63a79c961201dbf40d15d759a0435fa664b6aa3c402eb3f87d09f5d6796ef0aeb66ac6bf30972f3e9942ee4377;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hac237303a2dcdd588a5ac1af8de12a0c8f7471a6d5e929fe3eae2d71ce937c506626198fddcb6a639d73b4d002c7dd27083e04380699b34698341dfcf49e303723aacdee6179ff33848ee129a6d7214093;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h195ba3c786a2724cdd9b4c42c98b49a7a33b2a17029ac144718d517397b13fd3e4026412337428b71e8064f8fc5f31c344f618a5405a7fafe9adcb34b13acd8330a19164117a9dd0ef458f320715804b12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf79b129e3e3133e0dc562d2cc465d039845d50abb8f2295727cd39179428bd8dd019b0b39c5501cd3b3ae70ae8677edc700296cbae6b55e06e7ab7b0df04a7280d17b5d531e3bba450ce8f7f612959ad96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he88b554707a8cee679b392aa8060d32787ceed15c3c2b5a9943941f3844b88cfd5c8e5d605ce9e6aaf4455e2450a4efa498bfa6f6b0a865eb2ad0349a30b4417a0bfe9eab9fbb4a8d853804f7e56bcad13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h55b76d883d0c0cb1777508d57e8d0500aae0dba8b5e4487339e662efdb535fde776c12aed45d5adc90d6ce13c3cb8b7875de961c1d11b818d74d00c4e0461ea805e3a8ab17039a1017e91fbca178dcd3e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc0d6f76759573e2d4ad92cfe1261a31b6913c7f9d8119671116a8c77464aecba1c741aed9da77531d560e0162fd8ff95f2e7b654855f6371f7caaaa2ef3d8bd31b0c45d72b4f66b22fc579888b91bb5aed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h95fb876a617f63ced2633dded5e905825992bf71d83adf1d3b9bd7797de22190ef174d9e4be2b2fd6e527b4c419fa3195d0db0c1e09b81e9a9671b7c16ce6e2b0791f02ee6736f02f0ccd52240845ac145;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h73905a1dfc4878d5f448b45aebf7f93d24d17617b8e094c92e7c7ceff938dfc734c76816493423193ca178b620174779df750aa1b84e5b925cb343799e6e4e34d13af883e297cfba6debaa66bef11327b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4d227599c0cd2862157616fae96c120eb1166764b16e6569e95040cac18b59b1b3075e551518cba72c707305fa600b3c650062ea59ec2bcf3cfe00ba195b7c19c0de5a0ab8809ed98f2d415e7907b58e0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcd5aa2b5ff63c9fb1c826362d89fe45d14f8aff16f891f4eca60708a57ca2eea4e7a67c14c583854b0a000e6136d116eb3190bb18138a9fafc4b1fda80196227b4712e1904a6bb9acd8ee970a6a7527ddb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hef91a113a9b1a6d4a6d436d47ea68a094e6aca4b1af00ec007d76bd07d89a62c823870bc9e4b2331b4e3a35c1bb199f1d106f6c76c86b491a16e9a37de1dfb02312b5741345d7117a6dbba6c19184fb5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7d362dd79de7fdda92c100989a4b069ad500589bff109fb386d1c65ab407d35b64c4d6eba19207701a481f652de288fe0756ed5dd7af412e8621e73ebab3a2f8c51472fb9d2e7fd3f1565b4f6d86422682;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h90a933b84d4f2b779f2ccbd02047e779a63563dce00efdbfea1835a9a2904ed9752fa8ef39f6291a6b960b4aa3ff2c481746c0096a239a9f2ed2b7c594ce271d6038738528df5b49fdf031056b2f9fbe53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf41cf0fcf718d1f1d45b42036ef1d83f258b6f7404c689e24a24e7f31d38f53b8d1f1fca67f0acec17ef6672f57a285bfa0fb8fb3b69f3c58adb01d710e0b62d154aeebb04ce9070a4e15f46068a55c933;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h732de344cee618d6fab1bf250ef0c69def9da28def503e708aab35c33a2c5f47cc48a46fea923a0f024767b7f103092fe39cd3248c4e34a6c37cbb9479d600828319b8f4bd5fbb94531f1d0e6c2ed1cdf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h187f7deb5fb190e6b0563b6274f5e95ae35be49aeb4f9fada813bf03ee4168525c427c70f87d25067c9b0c025225bb31af2e81f50903e6869be20851de21b062b6514b83a5ac3a891c4f71aa4b96a5c6d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbbdb33423c91e9f5309026edc347fd867d1867938fc4f776b018614c0f58fc25232e1a78c1d22d3513bf23416299bd0caf4a70c5b3856eabf2493e1327532969d923627ecaff3d5b56caa5533d392e1780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfe369e8678ab537782496af5f39c7a87d8da45c50587ff066f6acb1cbc914438460b6e75bcc0d92079ec7704be13cdf2338a1194233d80bccc6fa6cebc7a161f9331c9cec3353eb1d62a43fce5d8f28961;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfe3bc49732b84a1126db4d7dbd6d113eae2bf759c58fac2ff3010992ee530f95603a7bd0185add5a1d50084ad4f494e7aa1f75010f242580b0e0e3da8988a0c79144c3eb56280b6f32a864ff90d38c634a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h850258c84f3a0f7858f2f3125a40c3a14dccfa68741591e68699c521a235335ca743faf3cd939f395807e698f7d3195dafac7ef884451d4e7c6b8877130b6d024ca23a466c7ce7ed71a548b59e236b1643;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3fc002b97a95c6fa57f04e47d993901d1e5ac700582aba70ab26c01b95c3c0954446538e49de2374a523857533524e125b331488a15fd44cbdbe6ae973bfa6ce613d5b7d2a8deff561c6b25d6569a0e1de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc39a3dcde1519792f0bc55481945bc9f4c65fff7e27dd97d0d78d903b2b2fce4a940a4e7a75ef3fbba66270f72e933f9db782da5894c2f5c000489e651cf0e348b02232e29826ca2a6cc4fd59c35c67b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd6bc750974ad948875a272d422c95cd91b08312f6667608b4cb1653d680614ae564bff12db2c93433bda002bf376c431409ad3ab7216c261f1d61f201555bcf23c697f2a475adf0c1d7212b1a1582bda51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h32cacd036da84aa5929730db6279fccb99b03ce5e87cdc13faf4a34f3120e89f13ec3d8a56b74aa6747ec236cc3f214e552ee95b227ba94177b9e297ee4df167673f6d9757ac9b1e20cc3e879e3d4a920b;
        #1
        $finish();
    end
endmodule
