module testbench();
    reg [23:0] src0;
    reg [23:0] src1;
    reg [23:0] src2;
    reg [23:0] src3;
    reg [23:0] src4;
    reg [23:0] src5;
    reg [23:0] src6;
    reg [23:0] src7;
    reg [23:0] src8;
    reg [23:0] src9;
    reg [23:0] src10;
    reg [23:0] src11;
    reg [23:0] src12;
    reg [23:0] src13;
    reg [23:0] src14;
    reg [23:0] src15;
    reg [23:0] src16;
    reg [23:0] src17;
    reg [23:0] src18;
    reg [23:0] src19;
    reg [23:0] src20;
    reg [23:0] src21;
    reg [23:0] src22;
    reg [23:0] src23;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [28:0] srcsum;
    wire [28:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14fb11b1536bef609eee2e748d7f88324bcb8f8f6d5d31eed1027aae7d68b67d4202fad76317844062e786ea807e86ee06f93b4de848511b0bc5802ca75279596be0086a00b72fe4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4117548f24649f1a7bcfcbc91fcaed2e38efb91789d92aa5ee67ae2a499864d6e77d6dd90667f24a5770d422612a6ae4ca7f8029f663da505ea8d37f4bfaf122fa116f7d88ab3fa4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0b09cd3fa8ce3dc3e9279383c3c213bd7fac77d79799db9f6b2baeefec772ccc0ff92a51f4df228e625bf5db6cd58135d86d2a6f224cb6543f278fabe56b635342193bf8b3f861b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h238badfa8ea244b112442b5dbbf3775125404365faf433d1e461b0b3ce8a458238df9afc5c54d6faaa77a7d57eb71d28904f0ebb2a6b0c4449b6717493b2c69f9a35c7111ed37fd6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefb2d963ee9adba1f040192831957a00dc11b059391bc7676caf1d75b05f05001e0835e7b443f2a3af791b3f98dcff8803af5b87025e859005e670c97b0cf71360f6d9d81bb91077;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebc27c5cb3aa1f27962f8f747186f84f7d4c92d89724696d031cd70a8f0a7c3b724f1a3a50b4721366e3889f297dcd92e91152af512f81a8296c86b0d37ee7d29f33b5d59a1ac355;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdde0e346110bfbe03d5c5eda664fda6e80efa828cd739dc84ee45a119f79540028a883c5a44fe8ceafcb1756a9249fa7b17af449d8d21d275bfaf382190dc670f764cd391fb361a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haede6fcf9c3738500ce98d282892f2098aa481199a0e7df09714d6a52db32bf16e1fdab8fccbd2b8a4d8755b94377f467b582385bc098373da813c6fb83220a2b2ce3c68b54c63c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf64bb60dfb3e9c1faee936a6d067f52175c9fced3377e82ca6290e5e04dcc196647bc50c8e7e8701bbeba83d61072cb4572051b6bf697e3d07d36aa6a6f5eb607c3628402101fe34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf0378b5debf00eff51fb4844aa32881364046eff84cae5d277a743e2ef36ed17978aaa112a98244bca5b23f3b970a7d9039e69adf8a81dd2c2018756cdf6abea6edb9b8bdb05d42;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24b127b923decc19bd7118fab116fc978a279da1390b0c78330e69b4fa8210925d365f1106a5f5bdd1e837821f1897c14f7e3a004bf622f77766e6f578baddf208d564876c7e849f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ac36481ac77463495e6cd8b6e64013f0b86c786bfb602510ce589add6e96ed32df9ef4420decaa78f266b69f8632eb203355311d07e0e8f66bc94777844f4d7b20a55a3b41f441e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43a9702f6769fe3171611efb066366775b2afea27577563971f1ddc66ea1d3969de26165a1d7bb0dcf76395f90d70c29fb357e3453d18449833cca849cdad8610f463da0db8bb7af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d98c5a3552db1cb6371a9db112e5bbc24beaa26a14639352c782320d680a8bd9031c9e962fc3c46ba039bdfc58e235bd976ec523fbc6059ac559f7e738981715b3f9dd116b4f0c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa874083e4d2db0557015ccb080a3f5031c2eda87622db1a22cdc5043de425462e34626d9e51419732e00d8deb6e0f4711f5057ecb276118ebdc476da7b46a02b6aacd8c1bc08641;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha90d65ea1bb5ddb11f075adc5d83c2b3b0f16d9fc6b5486de31ce7f9633f550207ec0a2a947f0db4a2a417a429b970345b5e336f1e64d8520ea7567abe94023a2d5d248f99b1ba71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf201cb5edd7422fcf3e42be9047a1fa0c58c43c53d24bf19c47e386a2825817697aea83fb70564477d20afc576db98ee0cbc1a508631533483e2476191f4070c5dddfd454a340b07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha00b0ce85cdddf073837f16c60ddd232fb44034217e7a6d6fee34f94076a9ad5d2b20f1697017fcb39555d24760d175d3c517f7f4321bb7f86e688aaa5befa0aa10b9d8b45a1e084;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52639775a1cd27eaa0bde3bccd29d63691aa25eee86a27fd5c352c77f59ad1eb2d4ac406ccbf7b967fb94e2c95aae803d5d0af04e66eb3fa40de8b182bb207fe47bcfc9e1749a15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ef2a37c702d12641d5954972af5f6b39c0fef60d705483d835807dedb5a9f04f3601a1a3428ee5b468c081777907945bd52c860459b425e83c15e4b7530577076568437d3d1dfc6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7e4b31a192ebfa7689e5a10acfba764b90fe7f40e23756a51e2b5dbb91f54d207f8f80aef38e6132143f8a65c18db07faa99a35c05fc90f21e984e82404fc3867fae59dc804e3de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac66570e78bb80b01074096b4d63b37439096ddede269245d6bea61aaf5e9fdfde297b0217b4f5113c3b77fa0bb0ebc35d886215c86229509c355a7c16f0e25761a6da3f5613752f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc378c9c95acd4ec8b528c43581bed0d78b7fb0a071b3360ee53933da82e16aa13b7e04cd0a6699e1be17547ef4d3c02861c91ce2d32e69130899c0928b44b29c527ecddba3ec84c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54c044d96c815887160dfe9fbac70e53b4ea557c9640359c4dff85c232fd68b6dd7b5306181e05ceee350811a5ad08eb500418aa19b332e31446194def2a7e3ac52190367433f45c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdabd0a5047740af8c38caa4ebefe47abbc13a73683ced0d02fa208176d34f7ae451d472b15d7d717a77fec4cc0f5b3a098ebac8e2250fd956ea0ffb46d18fcddaafe61d345154d98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26bfd68e703c2f465df3153e38861ce3af7de4cebec208dfee43ceeda5bb02c2bb54f428eb60bbc0c9def7a223cdc3fd44673b9c632f537172c297eb73edb952bae69ca2e4a5ec1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7745c73f0870c1f7d7273a47598bb999d13cc33efae3586b399d69bacc02e9e80db82fae0ed51218a0ce00d78e2f9bebe1019adc2a1e787c0f2a79917f35eba79501aca3899209ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5bf1fff7560fe96d48951350aab1be3491015f81c8343ebe5456e70b80bbfab683b75d4662eaff1c8145fa05a2a673d56bba489a04a984965d94f4a5097ed4cc1228998a00f08c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h314a86da8b1859e3c437c529b7fd9454edf1610321245d83a5ec4c17d5a7442253e1ee88e3ee5c0e0f88dcebd86114b0fd527219a5fada10d9fe70fcf055e0d9ad9f577fe9e99b9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha878df8254509f7334d0e8c63f3069e772267e3f94ae0bb681365de80cdfea22b4491180cb7f798e3f0e08b40fc4871f4a01c2da19bb5fa9cd0711adc104d9afda9721290fe3b6fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ce8fbf416b469fe9b9480db8cb9ba9f130a31f5428020d2304287de5ae00fbfcdcaa5a14e36d6350eda6d9241edf954da6cc0dac128d7888109fe5c4528855187df5b2734e4a27e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2d6ac14e93f96106a5fe8e0d7a2e3f7ed8c85fc37ab72531ac6930965dead77749514364086d7d2bf02c75dfad3a41272237db59f8620a60a3fd5c4b2de4d0f99766a7abd365be2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac0cc3402bcdc518d2df96be09e6fa00e8f29336fe08600865429eb8ec35eaf32821a7ea44e3ea6dde07ab9111bfc48c123bf2f0501b1143a32a4c16fbc5c10b03d1a851b87fea14;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbeef413fb21543817b4691d76849e46300e0c22fbe010ea149b8f549ed932c662a9b991450c1124f38d16e2dd715c10e7cb75cdc9b412821e38748f0789f669335eb4c9856af376c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h813e7662eaba9f4025bd3f477b27436ab6f321600539c7aff025445abc46c5c4fb12993147fe8cf7c2f50cb0a8c253b420a46d11f9f28dbd11470f475791eaea1b7e46694858920e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdeecce51d7ed8572073a9dc2cdb095568802bba4d2254080dbbf5618fad8ce3c818a7418d2f4961b3d1aafd97a94fde83a870b72d1535f85fd78bc9342169a4651d2726150eaa43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf3a757fb7ce85967245c8570e06459d183c21bd4d3914ff581cc403b09bcced399d1731b66d142f3d6e8969895ff9b3bb9174e52658a3ca6f2e2bfbd8e2ce500917c86ac97c2e0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e2d2d1c849f1b8cf09b8b73881bc7b1d26e00e2020f2d6f5b84e7f3e2a69660abffd3c5827a083590289ed0d87403e6b4ca6e04cc5f57b0b9db9e5138c00c46b036bbaad82c7f84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf99b662216f874deb09f9ac41f172be636a8b85d2b80481a9bee380cd4419e40670d6800729cb6b785e066e483baadf1679137dec0b2d049500d6bf76e821ebd14f213fd302b99f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f0dbac038e8f8149b4976ee5f2d51f1ef4fa898e5e50d87004488b02ca0b3de42a6b1cbb7f3b40bd2312023f6058d49626bccfcc0abbf97472eea5b3c3e26c3e63561fd973bed83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc800baeeef3bb60ff087433116f79f97de69653c147c3a5f44f3c297d02f040fc68827da53c2dadd9b949a38e4e82a249e6759550e6729c31a60b4d7d33a7d6acf203f6c496a3f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5955a8b0c1fa5f3d7a6fbaba50a2cb959dff27536833a371fba63246a3c876593203ed32e8378eb5ee0676a6dbd9f6240f9b7abfdc0a704155c04e9c97c299a2ac50c82415b0ce9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd989cb64e852acf080ec80ae9233c6a4e7faadce389c4af327af5560f67cd4a9476ba47a3f93846416cb5c24d50814c2cce972d0528502a10c743d4c664a551b0d2cc872db61b5cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56a9618603b2f8a9edf2e3f4a7a8b2744c24daacbe34aa1ebcf8edd3457e5845bb0d280b134c53e9966348f7cbd7b4b1a1cd428a4e15119a969d4d02d2f6434f50328372839a1bbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e95dd6531b22b90f8e1c1d1f0f8a84d426a41427ddbee5f926a44d156a778e9b8981b10c8ff398bd27dd09aaad96600bb8fdf00529ba04ad29843673ab6c1283086e70e1369ce6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc41dc682c93a1e69416184c68b54b5a908d3a060e03eef4d0b8ffddef64844dd0846fca7ad000e023202cb2942981d77b56c4a3d3e2e0cb934b7e03e869c51e350ceab1ca5a91728;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8db0c716e3569d47129348af097161ae5b3ec11b97fdc95984ce9a253a5b1134b67550eb1966dfb25ac324532e593e25f4572ee5c4154816424ead4fe8c15534d6bb9bf0c9eed63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3c823e357830c1a2f39f10e4a1331d4e52349973d440db529ac83b6f66fccb3b53554694ab032e2aa1415840a261cc679f1f348c54b9d6fe62f09cb98653ef137ebadd344e31eb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc65ab5728ccbf9741682af757c7ecd275b13832962296905ae124d3728df8ac77d46f17ebf8ac2ed959a5b9d5b523a3f86e4c7a3cb18c5086e1918a638e8e59a01dd9933aa91ff4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6736d7b26191bd38b17ad40e902218c7185818cb5b7e45eefc7c90a95baf23718960ed0a5b9c2768469afb3c36c151bf3c67c94f86870bd7186d8ce5e59a06b952a0904d0ccd3e34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49233a3a41f418975886e397444b63a860017c8ba601e63197738d273f961bb74f006bffca3622f4ba5eda00d17ebee75f7a90a58dfb33ba9d4ef3266aacba21a4fd385100b633ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbea997e48702b4a69d6e7695f91820e0fa0a79e3aa7b5c9cd6e380cc6eb9e69bfbc131c630b2c4d61075cfce0442f0a20746cd738b73fbffe4996aaf283438b742e3f38f99581838;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70a34ef0362287a06d769237d187e2ade4bb452ccf6358d30d4be8e975d5e68093c7c5c961300df23e13f79d7eb9ccafe49136be7ad77e68169c0b1c8c2d72350608ef3d462a7a6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13ce95b6fbf0c22bf9875cca7d9ae92560dc72e0875186b0537e622c6afab891fb4a42280c06d2732dfe44c9844d069036d2dbb6fa765907a8747d254ea1f2721e0353f69ef15c9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e8381c0caecfed7546b00089b278900749ed5b96993bc82fd15b797a9eaa3c2565a8a1c5dd017bea2ab7127dd0f3d7c7edf4fdaf5f9dfbb754badf49cd6ec702b50b84b51a3d0a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd299dd2fa128f5d52251265b7f30a2b5bcaf6764e542d03a337bcc3a4e7871dbd1dfadcb46297256fa73ec1ca35b285e31e57926697007f1a3598f1546d799c5afb8d330577c550c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb41162f07955b0242058f59ea8ab6c3b5230606042b225bfdd97c124c44a7d72777773b9503dd91a1808b534413ce287cd67703b2d156227896ee77a0ab2f4ac7320f6076ca9731d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22c21178f106ca7ced18ac9a0242ed7d7b84fbeebd3ceef7980b06254c8ac3a0dbbcbd0bfd3def97d77190f44c7c307bfb523a0326b9f3d57b3ec0b7e42b4dede0cc0f51bafbf5ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44721d7d9bcb09eacf30e65856bf1ae1c85e9b2e64285fe8d22cd422259aae5083fcd5e90233ad2d3034a0bab2c52ef3cc9f0af2aeaf710180bc67f535bb2da9d8927aa7bc7bb443;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heda2d95e2e5c7fbcd97059771930843d4355112da998925473d438ff34fe08737d14d0af4444b0df5167b3625563a205ff451f8211fc7087126866f7ed99a2425710262eed35ed84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ca8b78d4504573473a37e318a216fad8940f81e63fb0df633cdac3248212dced75561a5bb99c58f88138a0ce3d0b392002bbe02b00c1475221c23e6b67871e722c4ad824b9e5646;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bc454e3c18db0d9efeed46a75ac4c433f6a68adf5a40b1dbfd4c98aeed965a5ac3edbf17c9f8f8d484fd22fd2fb881d9236d04f35275a41915e0810b5736822b357d4f81885da67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95fe60a9a5e4b30a4318a3b2c66eecad1a087c8af218b498f55b062994ad35c24207e7d9a696c29fac2cc38cb3507afad0ed419885d9a1d9695884316af00c54e4ec4eb0d7541ded;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc4c6f4ce5fe9ed25b9dbaa6b1832bf7d04374b01d4ea787f5bfa33036a811149fede17c105fee032548cea7e66b9fa270abb93600fcecfc4219370367bde47dc0ded7fc86ff1bbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dc31b12a04ca0e3b98413656776a996fa5fa89e10a0fd7dcea2152e941da1f7b2dfe67321cecfd5123e881e49ca1f5de63a36ebbc6b43d6f08bf5d8871e2bbfa4554c3a42218aa7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67db0dd39b01a11a351464513a904a42edae6247a6fa22850ef3ceff4d96719b7a98cbfe2a5988ba9a554ffe96031901071760b29081d21133c994a1c655c8e9d339ce56ad7cea8c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd51b2ad14c00f6c4bdfc16bf800bceb6dc0a7be4496c066764d101732dc3305ee3f60ff9ff69329fa58f64c6e878851a157a04cd21c6fd7c961f90a1103be8acb97dd776b9f0cf8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a8809947af2f1464212e7c7dff7250c00a0324aade8ada7064a996590d2e4e9213d973e15800400cd701cf10b97a944bcb8d54e405fceef4b84c4f89b2f49e4b3cd5cff12c6df66;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0a76cae6f97e2693fbdeb24c4ab2811ebfd629760b75cd81e35f8ad30c30b995813477228cee52e4f227e873039033ba2557315e9c0965d3d29178e69e5019fba9fbfdb4ce0f8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78f1bac1df56f719786c8c27d13bc3003d1ea28e4dff2950f607e4445147b16ff0388a60a70e788b7e77f5fa4d492e3677ab12179d1d8eb18da24317d0650f9788bbc5206d9a7534;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h112e2f871c4ca1928d2dc4fd63a7bb920036fd24dfd3c46bfd284693737c15fad7f8fe6d0b0646990576f2d692a6fe05d3cbdd6f727653f6b8ddd68b6d9639175657177097131d63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32a8b37e911f4f2090ed318c2d8db9bd1e414e6e13981a91f8a4c0f20256a5567515946712f94adcc7dc88a4462811082c757c5fbf316fd86ae3812fa749a3e701e40e1094941024;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ce3c891d318788527043ee15fcb686ec837a3c2c29e2bd1d07e6fcbfc0723222c15e2868ac26347318ba09d8f8f6d6d6c190eea836788fb72b25c92beb9869edf1253ba70705906;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd64de37bd2f9faa990113a714dc09b48626ec59343d1d3a70e66e1ca7fd8c8351e92ff2236bc9968f9b11f51ba9bb69da6c3ba363c5657ca4edbb22948de19554a60dfcf6373dbb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h131291c8a2174c8ecbc37e5da9ace619ccb34cb8f80658fb739a83e5001c16109b9cff7ecada9b15c77f75fe691c1e43d3686acfda45b498ab218273c7214d8462452952ae6d1867;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5088955694cb04f7326228d2a2da0a36a8d902c17a242bf6873f3e0397be5d209386d08febe947bf3a277a4821f534b61e30e6aeb833d7b4e1bd308710dcb3d79720aba0a2205028;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he949d7638ff0ae2d76b0dbf0b792042c3cb2254282628567f9a2a788fdd8d1d557ddd4b4fca7e5510eeb116d32b95024e2b4e91ade0969ee7e73a1f8c8f7a73a5fd5bff6ae021b16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33c17056d747f48a44530ab2b65dbf6e70ba43612212f98fe88caf5513939dd84e9c3b5fc260a1e12a7254c5e88736dabeda33cd1f5ebb76e8ff08a5458c65a5bd60ebaa682b3beb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5637cef95a75b9328eee2c024c634737189b65077ef0eefdfff84ea9f4a51dcad714265faa82872e0b499c7afd9582d670c7c35d5f3c2193dab4e0480ba597010ee3533d16890fdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7412bdab8944513de74188671f50b27c26219543f98c77af40232284f1cdb5431c6f316137996792e3de88eaf5cd76e2e5f5ee7908933ff3e59f2887e96f59b6dae9e11c62fdca5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29aff2d52832d7211ae231e3ce37fac855cab15385182de99ee3955af3230dcbeb0077281445790895035e5bc2250f8aa2b2914d0a7a711e1b3619a148d4339675929fdec9bac19c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fc28a0a95299c977ae3d2f56fd39ce7778232e6e1f2e30288baa87af1b767ba2da301965a18e3be5669809b23f32bbc43d2b0c00ad473d7a23940de2ad68520588d886f5bbd8e39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32bb3ee8f0807060736a99b15d2d7b9ea4b3fa99c609817ad734842dc0e92b8801b9e2095c58aa7690215121e8577dfbd591e5d1baad29cc84f60b374a88eb16996d6b540eee3800;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5a03412d87a6a03930c026b8f4f60a176f48af09132b4796786162ae5c24b3a4edb4045e6559cbf64d39660734310129ee5f14d596d026976117a2131ab9825ec0d28f4436eddc6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h374b3bf6cb0146995185192e474d91bae8d8ec8443f2ad341af6c637130e6472eedfb878c0aa5567c731ae5c6d6861b37b29f7d1ffe3a539d40c4c68ad497fad0e69220e6276386f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6859292ef1adc2d2f35c794b997c93748c91599079a809d0b6c2df83644d89613839c6daffa8061088ac2e08719dff8542faa089e12634f17cde7c46d296109f675f9223a56cc52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2fa195e2119813034216af25e339a9fcf52819bdfbca9cf07dfe662a92bdb249ef1295a3bda371a76aad4815237e4893288b4e42948f1716c561df83b28307d6cbafe6608b76054;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5fa539c08cf42f442e5119ee9a3a83a8ae2189d6071431b74c2b8da705defdba1c4fd4bb5a19ef5ba1952c2c41c9fa7a5c75ae2f7a785d509c2d084fb4720c15f5ba4e7e9ddd230;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd76285f4a459e100c4fafb7ec66bb05fb39464fec44ff7c52bac1209308f876b2ca9c23f06e5dc87c6e8637f2afd8b9b97a35f67b92e4d061fed90530d327d5ad6090f02721edda7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he52dfea277baa82b40c78dc6823568fa49d5c147e2e0cdffd39ca91f4787092464b9fbc068bb36583b421a22fbd20fb9bd5052e08dade22e493578770a99da78f739139a8d430891;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf36f5c94abd69688aec34ef18c0794f10f7e7c84c3bba4172b68cc1670aeba2c80e7f00050062f8b82566d4e15b15ccbd512d1d98cdb02b48288f246ae136beffa401f274eb094a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6805f6c861f6f9a9748d8c4eb3f5c948ec53211c967de0cbbc8bcc4a78e1a05f9e33a51972a67bbcf45f0dd4aaf0f94428902c82969a5d618a303b1dc0d29cf9fd22e043c634a013;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f9f4687cf010d613f85a0f25c9b2530577b43662ffb591ac2aa60251954837d2f199484cb35a03443dea7a0330a26b217b6921ffb4fb1cf3f3a060ad007270684e93cde8499588d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9607b18f5e46ec52496e229bd38260713011777a15066006b546fc093afe0cbd92dec1e6cea79619baf576150adf292d453eb8712a83a1660cc5e0d66e967955ab7d7d443072a58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6f2c4cb250ac40314950c73e0c168f8319cf4683e000163a0133abce75eebffebe20d24ffe30f5b088a9bd180ece816b7ca9dbd02f83cb34831c0eb59a0815c35ba99b24fb55c3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f82930d1dbf93d2fc9a904416b3ea4d08d20a8bc0b0cbf11536474f96bd1bf2c22da5daabe9ea9f808ecda91db434cb4e2299bdc10256b7feb958a4c919e25baeeaf2336e97f76f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ea866de4bd32a1a3954b5f6afb9f99526142adce0cfec8f627d9d9899ad4d90745036d3ab07d46ae61bde014e917315d302e502566f4d7bff9adb2c02ddf7bf988ad0f5a8e7b19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h975e5eaaace2d6eccf6ab0562939301a8057655da99fdac9040dc43c672c2dd21c1acb6e19aebdc8c840dee149d10fa2c417f1648d6c72f0957e3a92dda23091af29ab44e0d245b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa0e800821d2bf0fb5b32745f77889bc71ab2ee81c0be689e4cf0026184e110bff359189a930981990306dd8790e981947ec3ab6707d2b71e1b24287c90cfe2d7f32d3a463c2273d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d0e1a59589c1be485734e72c93a64c0949dc85b59fc8c8eadf732f506c32b33cbfb72f29325bbf217c30a52741d3562d892661ff8799dc7c1475b8c55da02355fb469dc1f7f50b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e9e58bb6615d99b578e47ef8cfeba3d6e1e02e7791098fbf02bcc6d9f3292f98bebb2b3bb5f3e64c2de5c5a41d100e743126a697bf8350cbf41fb966699b16debfcc636d02ae30e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc93374261c12b8babff034b44227c1b7a114dfb879dcb7b99e7625f85fd2d4776842cd21ef8f6e65049f24ab9b745e3d5b5b6de891142507683d868bfedfcd852316d01c9498e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dc45ef61e7abda527d238a3f43b63d78f86c22566a38c28bdc2f2d02d554e863a6891e5d45ecefe3a9f5a12a7adb2a0f0f3275288dae96470da5769e88396d557e2c6051659dc5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9befcead2b31a4b2e8072be80ac091a18154ec0f0da678f1e88171bb981eab794846b870b6430a27c14e7536e5d951633faf73138401c13bda809ccbd0b49adeae5c3c82bd2cce2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc99fce4e5afb2771ecaf200f3169237b9136c39a57150f82cfe7e4867ec059a97dca812a902eb4eefe552fbcc905050e6e7d622e58f19f9f6ad1eb6f0d5b7818229d7f3d78d94d43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h357090efbe321706139fbfc46a013182ea16e4c5379721a2cf8ec84de3e03dd83760dfef61f3635a55d49742d04b6d7dd76b96bdcd765f3b6d1531b77edcc704c4733376cac23a89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cffd73ae26826dda0aeede9c3fea10df8014678677de9d49930e26be4bcfd37e527987f8bf3d68d6f0b414c1140fa09d68dc68e50e5657033c39b20500c67c715fe7b87a6465d59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbfea5dbaad61d14ca3d1e1095ed54b64924b0e577f1e2a09d0f9301e1521e82a8dcdc07d44433427c7ca1389f33d2b0e9023becd10ad444b2bb84ac3689ab1cea822c224cd54270;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha24bbf5e4a89aa205c60cbe70a1faed3d618c1cc79bc7add930774b703c191172d39c865d301529ede244c05644cc7279317fc2ba1c07933be2d3dffa3e9eefa53db96016b0271d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a86f2ec8a1466469cb4a5457148b71eea9bb47ed0ca382921b5b21b2a066edcc66431558f3b5f4297c34841e47b2b589ce471d28443df32a3e837f55be2cf42c6f4bcdb7f8ed4cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17f6784f191415854163c158a17b92733fc9ae902e703063dee9053c56849379cd226676a0f85413fb09d3da4647bbfbf7d73e3f0e8a874105ff89f5a2d17aba70e5b6cb2232c745;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bcb5299acd41e63a02979cfed77adbea44d16a0a906b67e84b8be1eeb68b4ce60af030d280c808b8264b10e53bb233bea2a40fd7c1d34c7f13f91885a6a8ab7d5163fe1b6dca43e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b3ab336cf946d69542873c1944e785a8396afa502eb1a58991c80d690aa13c5ff161880a36ff4df7f844983aa1e9333bece016e2b72f5a5266241daa90956768b42256f958c913e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1071b7a04ea7243d8d083caafc9e3f388321b1696a8566dbfeb5d42b936468e4aedc13858d19b086abef4b643444ce18344c8d37d31b056a654ecbd8d74f87f5a44b4d67b6052fa4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57f0c1febb18f24750e1cc9ab6dc5e762df74cbdd1265ad179e7ea10f27060df2111919b1fda6c38b2d9a8d2e08bd6f1010490f61f0bb13713f9b0c748011dcf9e183da5320e9874;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb610a07ae5bf54d2ec888130afc97cde29a52292d776506fd2c111948b53ec6fa5d4063c960c2e544b073513b43d39462b86943cb0d7f4ebbe8fd9e0bf8f22fbd42ffbef0efe3b86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee35f28465c32a90f645ec5dca2e68ed9a17ed1a173515c03e856307928bdf87acf43c80715dc9197bae9e9d533c19dc67d36b9e95b069be134b57e4e50982f39fe16d3f443459f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6ccb86f353a4e7e995e2c324331a21461ff2684f3f26c8750e638e44cb9f43bfc2a7cba66fd1ded41c736eb10de82834853ab2f906eb2a8757d894550e025155cd6c3b64cad2b11;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacbc9b5c78997aea6dc00ea6cb87f1b29a122d3de29e8fa12d6b4c6c04435932222f0d08ca5e22589d2f5a07d2c60f3cccd49ebe6f3dbf8a81b7a535beae2a67b21d644a179c307c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e4b16e3841411589a13c3cd0ca3e4b4a034ec142709466bbd6089d4fdb92392417aa9ab0b771fda1aa2ce29eeea59f97d63a98a3594a07e85ae75331df842d7a57c2dd8737a3814;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h198c2d3141ccdc334afb299dfb9d191718d9b1eee25e4cb9d1d360080c20e48f347ec0db8319566b1d728026745c9e1b6801216dd698e452e3c7266bfb55b59e84ea7243c05ee852;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf336be9421e5bc298621880b6acbce52d539ff82f6af1f8a11886a8a7414bd02ea95f6f61f0946bdbd486d0d610f76e5b2225adbefbc640c9abfad58e7e4b6403ec06287190af2fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a0ad41681a8e5ebfbe71ede977c7ea9f543b162e814edf4f9763f8b65bc5f503dc5d27fcd2d98157c435c2107ca86c8377f5be0744d3e4b3a82e226eb0756d96e0950ab94dbe3e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a9cfb25bbcfd65479e249dea1ce0cabc7f195aa712fa3826af7b8db38c0b9db26b082fcacccf3964a6753e6f3f4c371e50fc0cda434ba97782db4ade1761794b706710ba32b55b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf932b448afd2d77bb7f9b427b7f719b49be586b875bd8fe19cebb51f441226d5e17d96ee4cec0c53c02ce3156635951e50ae6585c6352d2b0a91c881119bd33ef7550372bde3a716;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70ca0dea8b85f9a541972a5c5a38e0d4b555c8d0a5d7d1a9403ceaf7dbb59029a89f9cb25e62098e8773288ca7cd7eabb33f0a5760415ad18e03e2403ddf5b11c2b4dd7741143b71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a6d4ec6a16b78b572f81cc860f4d189d5c08dbeae59be0bedc3719eead1e2aec2e3e4b8cc83d096d48989fe5ae5d5db12ca6500079bfbf44af03ca645da73a925d050dbde6febb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he67854cb403332ac4bcb8f7a838227985bd34ce78be062e6a864f9a5d88cc6ef7c6f6c6813e508e14aa9d635d38c3cef5dc2e041d319763f06ea01d404955f6e2d6c64e4de35a235;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e7b4939da84b7403ec6a33ece6fe0c8cdfa3b51ebe9b160706b59353fc114f690877eb2ee9b3635a46c9c6a9c23957e017b1c4028fe81b2b69cbbaee0fc182ac3addb1085ae15ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ca7775b692a1d5555f7c16501a665bf72aa37becf4a0d6415773ac4325cbe5e363b465878df49dd9df55e16990c8c8830752da4c2f3e4e2ae6d76d3e729b94804697e52c5148df7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h412cceff16469dcf8c44286048f141e920f301f34a47629e37d9182d020814f1a0d21e2e1e2d8462bbc17d9eb6bab8c71174cb762921690cf726759424092f39f67717847e46fc57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f5f8f3e2d9a0e18495e93c336828a0bf161fba47b04b0c6d8d9871d41d909fe57e4e0c1116dca52dd667f393b989fcfc6b00a9405a29fc4a0af073ca709d23d4b5bc7a0fad5d6a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfeb6260f8940a2c8f47af2e32fb1d33b9156cc15124da4f5d619870c0313a726e253ddd301ccd664d7b990bb551fa1328e54df8773c57fe33dc6e70f401fd040c4fcb2eaa17e3c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd68d51bdd6255b94ed2d325d1043cf383a3d223f23faa9629ec1326e7a944db11f2819214b48f74a57dc43245f6463c4782602fdb34d21d2f73c3ee666958adb709c07a9aeb73b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93531ab5df8be858f8ad7ce00c32dd900c3ecae74a063103f06bdef81f49b97defc5d9871f4d6b736551fda9990dcb3700f5ad2a3d4ce3d58e5e180fef588232071b7f4120f98a23;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b1beb0add16f5aad7033e21133d0d677c4ceac9e611d98600d4416a29ba0c256c2b23419e2e597abf3bfc1332d2a651480bd3760ca62111e3809ec5f81c2959e87548144f940afc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82cb42237bfb67db265b068b72660ec2cc8024329bc070c3aea7a747ec63c6de4c11f539d7f8144f8d5fc2ce2c74da2099ad3f48ac48f6d03d602a2eb40fdcef250f4fcdb154e8e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdabbe66f36658c48c978dc1b454853a0aab113ecb0a0eb9861e4056e438fd80104ba85f584fae884740608a62ee2a3adbec1f6ec488f927f0b20dd5b630dd9bb01c08a49fcaa171;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha63cb9a5bf5030fd4381b376e32f538f5b4a73071486c466aa8eddea1a101fcfe70190037fe35b6062d6eab9807b13e93785856d937c0b834abcf6c2068f665cfe1d792cf4cd6f8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40011304be8b9dab204c1716c94c02ea49f1cb6280c8df63d36dabe99635bd7989afa7ce3d9ecce375c612764ba0734efb6b20988ddb2b9238f6f2cbc22d499bf798af5762e305a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha83df3ffa9f81a75fb956045271e608aa720d07e4dad0c26c2954235d59a6f43fb4e6f4d37b618a497bd60a3b2f31f2bcc1521ff586aa81065913ce2aac5aa10509a1d2c6aaa864;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2a6bc062b3e22cd65aab7758dc8b1f3b0a812dc88fbfd86812f7713ae29e4b6bf918facc67acaabf4d3c1500f0aea4de632ec26b10bda90083f4b50c39168fa2841c188d128f10b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38ecb2c4f6bb9aa934a7576a4fee6b3bbf13d2482d90ccb83444a286fb6a4d61880a57c7408980ca6f2fae5b38a3a90616c77a11fd695caa715eb6a79ea6dc030b8237d09677d08b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h383e5043b7c1c6394b353ee36261bc2ee9601ef6178c32c3f1dff247f56d6120152d184f3fc08cad1fc813371e2b07c7bbc76e5f8d51d0f74ce3a843d07d8bf54bcdccf214bf27ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a9b33c6758b84ba56766d50b92005814f17235e32da35aa659adfc5220e88343e22bbde5e532673d02de371d5036b8d950ea1ca7f94e966f053985c3f0f45212acd1ea2e3b77d09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc63ae7c2db810c0238f3dc7cb8a498295590f481315b6fff7f9611f2ba5782ae0cd495f7e5dd0a74884b0d1d6373242c36d57c5824914f74af3fcb34f157bb68e8b5a894c9614e44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ca6597a2168cdf3406de020c36a06f0d5393203bda63b5d08cbc03011f4a2eff858bea39857866f2bf519f6e0dc5c8798e4417926d3a7780936a68d330aaf96df867b2f3a7e3ece;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h727bfb8f5cf269f8a731e29c4c564eed04a2d8bec33c5c890cf85970ae74a0f3797a546e4baac2571c64649c5190b62f4b862d0b407766ab0f8561e3cff9e0d7937e4b46745b70a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8f7a4e611388b529b99bea4b2f4bb1eb6ce400e738963383155b52451cc4fadd19616517641329a65aa670a196692ba62d675b2eb4b7cd122998cdb935c4d5d8062982f29e2f72d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd15e685edba2b72d24a9daf482024925743d809286365218c59d724008bb1d6c89f04de5371f15d1fb3a8c070f1051a147dc03353c42e461b6f9d2d9194218c82faa037bc1a8c666;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae8a7c3f719d48c08086e159fe9b7cbf7fcbb5239b4216c70f1a29df3163192055587d58442431b5483612691f0bc588f83749b93b2c4cc25d98d0a3981a1b51841d27b0c43fbd0e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d78c309fd8fc88f2803171409da4f723f1497c909d1fc23ad2e66cd328b034771858ee5f4fc9369e0a61cb293462e9843d3a6f0582d16605cd4a5d4060a261bea75f681522730ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6c2db9ee34af25fe5da40c11ddd6a8f51a0c340e149bf801c85fa089b0eba58d28a86bcbef86d5e0a4f05bb15f9b18c4bf2830d435ca431c59ef6b8f339758a192144b3459573a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16d2c7d3630a4cab29acef73e8b49896e5e5227e61c84627ebb61fbe0005f4c076e097b7f894dae1c35dc6c354268778d77a8ae75e15e6e4cbd7c8ccc175d5b70b4f5fd250ff8ff2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h303335bafcd0d5f7cbf47e509c22e3291fead1bb7971ff22ac767f335e712466785bfd24037891c5ad5de7a3f72e48eee2c90f554d92eb58603d3f9a5f20f2eddbd35598bd4c76c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7245d6adacb1b92dc17c362786f2e9c5cbf00187394d23d17e487cd773eef1fe30b8a2fdc295fc76919ae5397a6d0e271918c00e867dd7e3814c1d78dc58d3ace28b1292219225d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4b5745e33fa8d4f657febcab9ae9df6f3a702239e3f791c86b26db1d48fd25956f3de158ed086d30a8d8464b776dfb8cbd3f9aaa1fc04e428d852e776258e4f5c756caea1422389;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87b8ab8de25a856bb3d7aaa8f8c584efb5d996ec8dc2180a1dd43cd25495e8de0bbd7dbb20331113cf69cfac08d5ef0d5d22de08465dbd63f12caf4a300c26a9b3f06d2200976d4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h117f7f599af591201d007d680e657f61f9b3a7d42bde3fb1c2ea31bc1444902df9a5d380566ee9df4a1b3fba8e2ad9eb3b62ce9f0b9c4c237ce2a9c756e6d606d2f824e3afe2e512;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf0ed5f39b7d4c7ce4bd44a02791c92296d316f61466d7dc71f2ef179c1bb6ca32c981138ef86d8936ea6c38e45aaddc77b20769fa64a27e4ab230a4e8d57b088ebe062813b12e49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf4c9bfbb736acb5a065a98aa29ee72db66baf93a4bc1c34dbdafe08f0d30e5ad342ed57d20a41249507fb14be177ddf7c3e11ba3f8cea2cef007a6b5c2f274908eca813ae193ac4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfca66b864b71d3f4aa4c04584bb452d5d88569febcfee3b1e584da3dd9e9da7759fc71f31a5da1add6c62cacb583411621ef7859d68e97e9a483572f2c98f613fca48dd49a97eade;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e1d3587a95d5f64fbd89e975611ce76fc25189c2d583b1d676ffe71af41f9ac4f9558d9166b95b92f4f7b070b4cf191f2c758a31ef972ec327acdfd81b8dd541518e777c34936ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1619488bb3f8103eaf684d12159de07d99cb7961ab2f7b33287f3c2d00e4fec784d12cf29d534bc30da215366ce7a883191a41ec35cb91737cd690fcf20e813948ff53c784c5643;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha92050e218ddb0666235dc5fd56560409a9d878071821f16714a0a0e8ff988b42ffa6a88ec571dcf1226760749aba3875321b65b2875d72796373e44ab81d28e2c0363aec36a0a85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc8efdfb7729a3d0f65a310538fd8b7bdaee4739144a8d409c60f74f104c47d8a9ddba150fe614826cda1217ed4b7f5690fb76cd29ad9056ded332556af903491d7dadc41d0277b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc94bd8dccd26da9ed5de73bcd902398c1d3dbdaf2a619c2b3830f0a0e68891c910cabc4c294bab2ef7ec510748a85c3c6d68f471780cfdc7ba0d916a462a44b379116b8646e28317;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he881571d3b45d575882bade14c555bd33d96024fad585682cceed2fddf3839ec4bc107310e1cdd1aee007aee16a1ac34bea1e5a11a6e11da98262a83444a4ee10fd2855fa589b065;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48628e7b9cb6bf344b30d0aad8663bd3fcb80f6fc1b37f32646a0a38f2818402c52554471ee4c4f291ec5be3e270133b0d285c60e69561e780d8b66cafb8439623f4081d586d2a61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf587e80c1acaaa8908c16cc7709f53846c39bbcb95187320aea6693df55da142ed404a49b72f50ad175590e146acc607622771ac0d41db88c51ab6a77700a1c36901e4e136dc86bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b994008b29ef4e042998790a7cd94b0e58fb43bdbb98866cb0ed2a8996e330c44e0ec3ca62dca5612c11504b9446dbb3eae8dbbd966eb9a105ff9b5894b97019263e7e8b9aa4f86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ddc03f4c869cd3d1fb1d17e6d26fd6db97df3e8ce748522bca891f4f07eb1d56e7a615f2ca9546b2776ad86abc8c9f338dffbbd1727c11139a1bf1685e384a84765eebb79c8e150;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3d4a48b9f077f05370ebbab78ec9a72baecd02c7607c2c09ca09e8d9a1e473221ddfb7c7798ddee413e47ed7ba0976924ee2f7ddba8f58cce32de7b408429532bb848adfff0ee69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70af8475d8fac76552ab5e53e26616e3203f1ed32110f76681b0ab6bf1e6f840e6fa2e571fde0985a7c812cf9f4a77c40944b3349ba23f3f4d64115d9044837898dbc2a8752ce71e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf67f1127241767c2abd90dab280b26669e7af22d795ef7c71606639c02300f201ca0106fb253375a0b32c2c9895ff2f2bb93a8d7f8314a55789294c51ac2d09860a6c07eba643cf4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a8d1ccec7eed9f86d6e3ddc8881b4ddbe311dde7d93bc1fd6469599ad0c54717b78eecf1967367d55ae3c1e20deea770bf2eab316e185d2ab8211832846376c1eb45a4736afcd39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6afbd7a76cd1a494dd21312b5134460d2632f8a70432cd93e0b9b446a18fe475a501fabebd56a9a3f34ed65dfc24aeb8522ec3200025d82fcf3b2be2ba28dafdfa65bf123129c07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e5d88c6e2551b2e5b50154ad4f532a4d7a55313837e84fcd539da60af7bfe0d0e99c513633fa23588d9069093c5e0ff5908ab63e9978bed9cbb98af8f659e314294150b58a0d3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc75207a82b1f519314e2eb5887ec355865731fdefc68565eba0468c8714adfbab9068e15f63d11acf4cd9c357a1a2c817842567d294620a3228fa81849a23f83080905eb88f2698;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ca5503b4e3080966f80300e249519f98210c8c3d903aeeeedd9ee95fa26a1b932f392423abb7a0209bb0d8318f768b27289049262c24167a1169d7083aef379d8a869ca1380539;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39d944fa184cb883965eca9177a7b2ea82c383815dc262b7e3e980233b9ede28eb8bc5df38c84595a2f40e4a4638035874b65cd68d97f5980146f6be92ccec92dae4fdb232c49b17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c3ff2103d7dccbfcbdaffcfd2eca1029473a634256bd460b95a8e8d5cf079f837a41ec16f7cb7f544d0ea77e430955c6b6140ea3b2d41696f845605bcd695e09b9ace12e9f0c58b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5044ea39af125c2cdad9159949172f9cd561dd72ebb6a4440a4d408794a23ce2dbf6ff877859458080f72fc228f6351937aad74eaedabec12257d84b915f3d6bcd53d42e259c3ad7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c17fc7aea03e5e3b82b711bb0442ff29abc091db52da85b2c8f941248ff8d39bbb7923c87f20ea049ca7c3bb695ab586a2b3caef4f396c5203c774145d9b1bac3aa00013dbba3b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50ebbb94ef13a5b70ddba197d2f652930430e0fd229c8665006d3a821bbe4e8553c32ade5ae1a82834414498b6502d9e4996b7dd6b4279d007ea877817e1bbbdbecce40cb0d34a0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47a808af5fff45d1aee3df497b1ad18f413f9bfb4d611d682203884834d11bcb91e76bb3a54a65e3ffa246fd7863eca6f16361e7999ae7d2dc5ba13376827661c432f0a1f1e251bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf12508a887e05cad9d4cabba8c9199e0f0db3eb1da60a5e76d4c13b1af2e40a5ca6658868c12b7b831e1c57743d94ae00735a4cf5835f73c355f3de3ba1fae9b546fc5b678c4431;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7fe2b862d580ff263465d42926ad96b50eba816b0cad9fab19f8023188da2622d1093eff33da29efe77e4a95d7c6cfcb4843a392bb4564de55d3ac264014b7c4c46bebb1a4673f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60b0552471d50cc04a3fd905db5bb6879696fb647389b8a97e389c2106b3f271cc265b0f8697d959f14c00063b6f0b5219e3392c9cea7325f9581203dfe894bed0272aa3e774271a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20b4b983f3b1445ff2db29d76d014a6bde722f70fce08582b954625f0523aefa437a6885c904be82ab1e2fb6f80c95e0d99c908156da161d2ed65752527ecf11733b090ac8aa2918;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2a520bec1ec199c47ab2e68a6076761558ffb1ecb39a9dc70d33c91f6ef1c2c5f7764fe77c1ffeb1703b6fa92417cd0ec7bfd5da76e7b1f2cd326e9ae7921f77c63ba995c869465;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab561ed774b5b1f7590cf770130e5aecd189724ead414fe54a4f406382e6649537b8a4d802aec2117ea92559621f31cb367b8398d7bcb88b72032dd738e6fe76f343d7cd09d84d64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f54fa64ff48a8d25244b25a29106d10227ec495234d39cbe943a49afb36a291118028787d71abca6418bf62922a18c6b5c89c99042f6c02db3993263272e0ed0bd1927cd948ddf5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha616a9f5a08a03ff224a813b505c4e91a2e72d9a9e843d05b1b52dae72fff9a9f3bd4eca9f5b7c115e9c8fd1ba6c587b137d92f75a35bc28228a4c4fd5653c360bfc9e89c4017446;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h650f705d825425c4c4e32371f534794e5d8471bd493ebc75f6e47f6333c245ff93a336479e15e3600ee6a9a85d85df78050ddbf6818e421cfcb3fd2f0974c97a7e5c2ff5ed25065e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a629c04725a074e298272bc22b6aaf699398f6e60a72b2223242edc29d5eb1ee32a0b9b4f1db72b9333cbd6a19370502342cb49b9953e4f69c7812fc48a9b74625a0ec721cb6a0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb50d92f444beb9fbb2192c0e607a6722535518c6665ec7052976fa9dee3ea8b0318a502620c4ae11b7a5db563798b176195fa65e37a0efd5c60b921f3530b0e3c3814a2bdd7cd1ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadb53f02c800f9fe40eb5d5b079edf4f6e99d76430ca5b2e0a4516865386c27be9c7d35bc1c5bbd65b77d0917f175d37b9f612486f23968b3ec4880bdb43f1ecafe3729cf07fdd39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95c6cd2f6d53ef915f174138e0a427b67a62bdc03d37b03be1beaa26a50c9025e41fd3c8c291e7fcd7584b6ed76cae7c03527e3c6ae56fbeb9425cf36d26d43efa5a01929e0010d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h134485512c54c21fe725302fa26d78cd34ba7c5fd93ce14f2179297193afde2b0dd832f9c1dae9db7b458c37786bbf0098c95071be985e944b2aff9f138e8193ec00b838eb334316;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5abe9b689be9a8165d01d0d95e06935ebf5121d17e3ae0a274e26c970109914d74c408e3a5e099caf9eb6b7bcf224af2a65fa01a6fd99fd63e1bb5d1f31269a6bb92445a03a0ffdb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c6ba260fce964bcb10ec4c8533b70fde2d192ed1686b75e36a6a2e73e8e8fb66f223c838af0ab4ab7d3e285dd47c328306a4fb0016802aa8858e0de3361162aba60286ab19c2ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaecb723775f05a2c7422eda18d440922ef017212e6fadefe197b57540f24272c778fc305fbe6d1dded0404071c55815e9598ea49b3446abccf3c3bb572bd85beb5273456f365e6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8c3d57fee28530b6477c034ce90f8d6bdc5e8f3525928fcde29948449eccc34ce538dcc98b52efdbd46549fa2c65132fd62aed0d6975f397685f62eeef9c1b7fdb88a99713b585f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26af056ee416ee43933ee3cb09aecbd2c16a38721fe39d5672633a5dc2c4df948efc4c152b4cc4ca9e68f0f9430e9a19779599486883a72b9a3c1e8d6af3efb3ed6ec2a6a81967b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bb5a7a0bb6e7a313cfcb54e4cdacdb9ed7992ada5c695ac07559a3d08fba43832ee7d6d61ca12e6c7fcf93dd4957439594e50bfce09525287960c66664b7411cb5ef67377f962cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ff6a3a96c39b81ed1a6d3ac1ad8ce892a641a3bfb0a0007837b37a5c111c287b809f8b034bddb3613e8649ff0883a348f78a717dea9e772ff625f9aeeffdd2f9735e68112941a4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc667baef1ed9b03867401aff7ce989d8557be4df2ab06a5dcff4403e900271b9cd70e13a8775cfb5a66b37bebae24343bd39c169f824e7ca12b2e0d5069a6bf90fa0a0ffa509e2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8474e0e851a4d146b3e5a351a27a0f5b87cdbd059fb0bdc9614017c56fb5dc6ba803ab62f5babf523535aa659fe150d16ce69d6e9c74d2dbfbf67ba8e2267d02c0a3f12e449dee83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97193f5f5c7a67958641f515a76c569c10c9fd0fe8e841e10140cc0db3cd4ab817013c15837abe1457ee80641271126b00a47b3fa7448a44e987e78b19ef68f3395cb82a2b45b8fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h608f35e0515fa764485b9e33e69b0c082201fdea6fa857246cba381fd0864d593bb4f6ca4353ea9655e3679d781cc55db59289ca69956fe90f1a9d838d73c416ea553dae26e24fe6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65234a0f54e5a9bfedc24353a65cbb03dc04186df5f49f2f91aceaf12776bfcf10f93a4e00ea1af6054d2f06c209f0157f22bbeffb3d2caf9613e4a9805e13e029f94fcd0da22ac3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61d9e0f80b364b8f41aca42420d76fcd1aab6ed841ff5564c5cc549cebca83473ba42bb2f2990f4ca713ab86b265fbb845754ad6831171a40cee2b2d580e9221522632672778e841;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a9d84d95624c37fa13f8f86dbdbcd761f6ee3cc5c6a6020323b26bf61c0e5329e3ee70c63db60e5e5261971495f54f2e8ccbc6a2ba3b3cfbc2404eb7497eac9a57091a3f6cb2fd2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9519f63617df6e28628c32a74322bb87060980aabb61c7280b4a81b9cdba97da7b78d0a24d39b4bc4d69705119db339a739682adffc056207cd8d2abdccff1382c678cef7c6fe89c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a5bb087c76fe1bf7b79b1c70acb6a413ad6453e2ec93be18fd6b0bec8788d2fb094a27acc1f9e6995aa445547b73eb03677c21521e6b011d184a7e3023f31897e84aaefd8297799;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7e8b2185fc25ec3cd70eb028eba2902bc2a629ab328aec0fe3291b7248d52b82f331cbe6b85e2df8141cb22e5edb5320c03c06ba563dfb4300910dd5e065fa3e7bd8f31179615ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d2c34ab4bac1a6f1d1480d45880d149d60876ba28512d18a6fd646e92cd2937f87f4808a22952aac4a867ea2483c79a41b34bda2178497e3091477d1c6395215110bb54f6b97aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a91daf2cce2d6de1b2009e58c4a6d6e690bbfa22563471f6b8c33811658d808c4d5239d9f1b52cc49b68b37133a9821653d651cc30e466c4b1c7800f14b5be23f9d91a1ced5685d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4df44ee64296a4b80942936b42a0670068f52b3ae4ec68698c06147a8f74e58ec8894bb7adb5d56d32c6142067be9ffe70d5e8c33332471f6006f6383e2f60db5882c3b7436ac57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79c4f7865b511b19d73d6ba98c71714a12dc7bdd2c0de66840d604299bd2fda05b589c8f0b602a4be4b584055614dfba75ebc3820d71c2a684854115214a043105594181689ac2bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2579ab8e5cb79eaae93ccc0752f579ab911d23db07329dd2f7be647a83ad9a926b343d2751702929f43ee6d86df8251839c5720eda9aee8569dcf171ab91e7b11ab621e15712e6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha803116639b98d8c475b0f4d9668cabcc5b8a53f521f05ebc3d79a007e9fa08ede3ce5207a1a4fc0b95c6440d6f1418180979742f8a76dc9c4001afa14eec4b1a8f67b514c02ec4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3920090ea5edb3e47315ac3aba3506c2e8c0fe41ddad5a3c49436d473d20b2abc5d2c51e04fc1c7e210fb157e4760262a34107b7fecd77b443a2ea72e1b23ac483505f4fc2e13968;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h972e6d26c34865c450ba34031139ab973f2103dfa4f9b6fd1b456a147252c823e26fe911f5681e6c5c1c35663c605dd9d7b9231d8f2ac99ca6524c4a334d17f91888aa84252e2948;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b3a2fb8d0b033ca11aa8073b438607b48b8da1b08e4e8dbe547f698b142a4da4f98e863c9e1634af301e32ec26d641274cbc59d4306d43c4484d9a9b88c489cd361bfd65b965f17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80bf97f7a6ff3e91e98eec29b77218380676b99ecd5495d9d49af9379aea155d9b375ee6973dd376cd6a0d5a0395b335b2775268024ef5a72742b623823235da4b80fbc4b4c51a8b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf04550675c73314a626f1ee24983485d933a3c47e773bd3552d780e93f97dab360588845bb9c90757451b690ef88bbabd633366ab93dcf66d89f06f0da7fd67dd992f3efea5bb8d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6f8633d8aa2d151603c707fcc89bb6767966163f8c3664dc54d7c66bfe5149ea42e7ada78be302f81d0cafca2fc483a82cc2c8685f34f4ca8f389735ed9403a646e835814887956;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5082caf63fcef0bf43cc187fd5abfac1b99a11442cd0527b47a0dbe9e983905551e8e41b7712523fd9e4fde274ff8d14674809e2a7b3cc9ea3aa5a74228f0d9be03e993e0f7bbb01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4db8eb2a4bd9161f4ae75f20e91681d46213c1fa182c50a18fcedde8c5cd62184b9bbbd4c7ccc5c2a7dc7174039a557038c41b60a57b1a2a0ff56ac486b5272115e2e928c54ad407;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cf1ff8d7ac7030ba94ce281f50da5ebb6434486c71ae90f97ce3c30f071bf73e31749da640f63915f1dcda43fc62677f3f7a7cacd8afd0fb8e4cec969bdeb3a795eb2f9fda0e203;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2aa4d09199cba98ae97d882023625c285c2a12cf86e6637088e65e411f8ec083cceb440cd1e16ddab60e514cfb5a7fef01ef5e9dc2033cd4bba369f881e7e02cac4ad8a7dd163f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he735930fdec41473dc4b11bac4e0ef9f1277a0bc7e57f341c9f05b283c3725e6953b3db4d8bd74012a1805d41c9fb9ae2e93503d16dd1a55bb3f873784ce9380203f736f8e8fc71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha417d356d9cd4900e539ca2f9ff7ae79110bef0b69222e19835b174f8b1ad2f91709d04e340dbec85809c081de18221b16ad34d4911dce7290110c124e6be3fa8657ae448f40b076;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc876e82df8bf867c3683ad5f63269e789a2b97298e85950524dee57be5af2ca94cb5851fb80c63162b74b6303c2c5dcf199ed41339bb34111e078adce69c0f808ebcd6062b13eb6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d765147cf7439732d4d920d2c31b4298e122461d78a9e749a12e5bd40b731c55deb22de639286157b778179a3b4690a73a3aee41f54102a2e11b2de0328ca79bb4396570e5838ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb13870b49bce925c2dd48e0dd751334d21b684ea930565c9dc09f1a8103aa337d5ad51f19c17cf93b89cba43755b075d2779a73bf381519bcf8d8687885b4fa67b3faa1ef47611ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19eb4d780af674741e41501034c76cd4a34c492868654b12f679e5d0c55e502b17dd5603ac3761a0ed9c2f8ecd6a570b9be7bb2128cbb21f049c172b6e8edfdc7ddb78afaeaa1199;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6874c58e95ad7b5cf992de4e68bc0561ab168cfacc968f1732e9f65f8eefc806d892c039a4e0eb24a2c8aff5ab3cb3971dc16006772f585af5591b7f5ee4fff85563abdd65377259;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcbf59dea82294a7cddd51489e930e1c1bf3f04c59b3a7f219d0d3568a9da5bf21ddf90ee6577ae136c2cdcbc0441bb4d4999ef1129c1e4f7469887a5ccb2f8579d2e5ce82cf9f58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fd406098086e77d94699a6558f6ba03daa15e420cf55f426cd880f60f7e1544f7a8af2f5e25218d38885288ecee63245e857160ea4d3fe7853e3615a6e214b22e1d23b176bc778b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b6342863d2cfdf92ab0f67101eb07755444018fc879661978290ae0a8546972a317d0601b4d3c0ae8c3aea61d4927ddcde40e773433c4c936f87bca287a16696857fd9c216afd40;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40a03d51b87710cf5dcea4366b30fb2472df40c51feaa5db0b4fb3d46891a6d299a203099319c8722ee5a66f85ea4d441b875c9a0e910335e82d767d670a4c73d56489b8d8122cec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc70a763533a1444256904b900193009e519deb7dfe58069d65c59bd401f048bda90a7963bcdad374e48d29613b5b5c7bbea4d706e6fb00659b4c7b62bfda18fbb31f3c71d2f37d07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf021550588faf37d1282e076dbf20d015418a89c01625e86734b98a5f8ebf646d834245320ca25f0824283cb4172ec20ca25a6f2bf3b3d7cdc5d919e5ad090cc3eb4b729bdbf4811;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a953c63cf2ddb6c7893de04463c761ff9f5aff327b5b312a2fe6dfe54a484955b327e9fea1231d633371fc56925382386fb4217757e135b5d1d4f8e645fc5c63108bf4b25cfada5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb222411cb1e19a79c88c02e2373cd69893e7be6b8ed4e7d498ee6e7c68552ad29460d2e5a79c2f145e1302fb9418790d042eb85307504ce05b0d82bac5085f44d0f36834fe3fb60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7eeabd857bb0be4eda8214f76513eb21f7d54034c2bc6e876e7289be731ef7598365693ec4287c1e44f30d6af4eb7e9530904c8a639ab081fe8284b3d873774c8498d0888b1da5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddb3375eac7e4b49c1ed8b1d9f79b0dd2ce65d2967ad3f6b43f1034e0efe7d208917d2835dde59f444a7affa3cc31b710523b4c0bbd9f969a56e3fa4988908eb7f28c92172a4745f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48d14eb67b22d3e073a7d3f8b4c1184ea9d5027444e05b7ae1c1cee81eb8c62292be1dbd1730db8c8387c6900c1a2e4695f017cd71c9cf2ce2c5d3a174041ef9b29e492043c5744a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32a265bbae4c5ef009f0f2c35394e43471e7c103ed731016314b057cc71dfa7619875b374a1f768dd5aaca990f1ace3ae989fa37494f442d0761fda60ccf6b3adf89bd86b41a06e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha74cd1d9b96975a9f602ab656a08d696a5a6045c271bc67f40907f0460176605e5449e6c2a3ecd45154f0f52c375452186650e76166c9597f847ae3525786e15d4cf10b16e5c9e45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccaf9b49e4651e1301616e898d50baeff12cd8de24f20482a04460cde6981a5e8997af26e81ed0e24ab4b761d5803963aa928cb6d57c91e7a7dd90e75298202dbdab59fb6fb413b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37987d9549848bc11721ec890963a45aa09493a04b454719b3dc1729e24c026f6f04c988accb86738ec9df39ea931fc631eaf79dd8b30f7fa2d547c61e9199b97b78abce89c1eb5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf8cd33150bf5d557153d473a055c9d9577e2b8f9f7565ad1ec5f57da083e46aec22e32cf10801996e54c25fd84b66aa0825b6a715f94e150837607e572f040baf74275c83cf57c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36ffd923fe05dd6be382be2cdfa151d24fbc7f0d344b1d5b54286b1b1cd6f5c3fbd7f59417a85ebcf02e7e4c00200300246c6aac0c6ef2ca3e675a95c2d58ae59219d7e182e84c62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f7133526b3c9ac45ce23aeeeabbfbd65be6c686c081e64c7de89ef87684d7c203fd780784ccd06460773bfa792240ce3ed9f60c3ec7445f9d2fe621c0f4dd452afe66e202df452f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbdd2631cba6a5793c7783b944592d891bb57027dc966c7566217fb5daaab7dfbeafe5815dc9115a5c7e3d83fea5c316972176be86bb3d8e893bd1aec6501ae0b427afa5804d6ac3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68a15df2cb05c5895f423d8ab42974b85bc5c2131fab387280804c349e51dce9c9433fee3664761f0ac62490955b1218d946118042edea192a9d40fae1f8379effe09a829b83d7b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h716f4f1511609a9f38bfbe9852e0183c45d7b09f1f501c4fa7c7917ef10408fe8b2dd03e16e6e4328bd70d966a8bca67a4a804f46676ac70c842a4c9376841780f0ac7a9e473166d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h738b6180a9ec227bc53fa21aa130bf965376f27b19536afc38b8107ea60832ac5cf27aa59f5895aba6af792363204c410e123f35f785eedf7026aa26ac9014a226a2f6db973d33c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc3342c9261fe7d514de1749d1e320db9d23a1ed177ece2c359dfd4d1c0ef08b98c526e30524cffc276af82bb3107c71032d7f3f6889643a865e4a570838ee3bb589594d7e5d1172;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ea4b98541195b27ee57091cc35f6abda92db5bc88cc90b699b5934e7d6f8423cda4916791cb555abe740f1d7396f10f84d9e51717b2dfe32af7d97738b41901ffb98ef0faeffa17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf51d71c37b6a433520f1856290af18ad9c50808b4d43cc1574e6593cc5a12b1e5d7f3a59d09e9297ca04a472de9c2626202a0e7e91ab272a48959463876454ce74ff2f885e461ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a360963b3169ef793b40e12695bbf359be4435af3e058ea1a1e194ee77cce52979a880c1c58d2cea498fac0642fdf5fbc8514e2dc92871ad1ca919e5228a3bf05401430a27359f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0a51945e362f48ec28e40fee69da8460f25188afa0328c4cbc6da6a4774a4cc0b70e3b38a8b293218d45111fa2f548c9af56e9e720f07b37f87d23f70df10786b0e4ac8768c9996;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1be27048a8d3c65a516acc322e93d5151efc91f3101e166128c44dff235a15eb19c169b8216464ec33a0ef18da002a925533eb7f659ccb2afad8d6280f8e99f2583134f05ffc728;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h892576e6fe7a46db9504bcdebadcacc6aa8cd04ff89909058dbb6583c3a95fb629b48d077cd7a2d1d5a5413c8657e11874d08f04907014ae9d911de84819ce9ed0b4a09061927ee2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30576c59f52fad76b9df320b15b0e1ca773a793bb6ee92b5d58b66957bea6019d72adc13b0bc549a5511c63a8a247bb5ef8b9b1ae125fc1b940e2bd42236b842e6c791b4322aeb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha07920ecd71d49fb096140d61e46fa5139f1ab5b06894b30496d52ba0f57206d343c3e1137f84825df4c560f865adb14813a5f0f05ba11caf0ca87e62d87d4259cb5cb79284b1a6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd30347e5b5a54ae2883024ba56eca23e788f3badf45a21c481422f7c724c2a14127c427d6ca9dd1f44ef1076a5a75c5ae6b371fd592f7885cd847da793b8fdb91d670df4e04fdf52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f40ff8244c010981207062e5b4f6dda2e50b6fd1464cbc68254582131d3563b1a807f58081e151e1e124dcb5bf9ba5e36df0e78c45465dbd06566c0dee12716dfeeb4a9d1cd95bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda94f30a57346f4fae8e557de4ee7363321d2531e7fd769fcf88b2e38752db8564b7238e10cd716f207395b9748d3487ac10bebcd5dbaa2d3935238566eb2df551a48de5cea3ae2b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h545a97d8f110775f79c58753f784ced917e2c237e37f65985b93da35acde69a2b0f5fcf01856f21f07eba7699ebc20ba9a9c16ca66ff3206545e86a0e5aa1dd8ee503afa996e4469;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbd84fe6142869f2164289c584a72696de0f5c6eb3aa227040547f3816af6254de7d7a22a12d078a7f07f08d320becb2fe512e4f142c3546265ef943a1329e45f2df0a851e1e30fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b18c26e107ad7982e69da0cd9839ae64d76fa4b36e7e2f727342a557ece2bfd186f07bf76e87c3da9302a6c256494150ceb35d1ab70b694cf12e7a49287db0d0d5024126d72f765;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7144a3c56155e4ff19feb61efafd2147a167dd99b45c4d5178ffa0dedccf620b9ecfecb6945c31c442692b6d000257ecf69873480cbd7128206fa45a9029dde983aad96e56282f6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5080a69c2c113ebf06a8f813ce9d58c3626c9c667e7b3e1007ef748ad211d18c00366c59fee832454564190dcf3fa3dcb5682ae5b82a0225b44f1ed0bf244b0bb588336410d0aa86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a403809f38940a840ed0318d0534dfd87538961c317eb0fd905b1fa53c9531f2163818c60d6feeda6815651c75fc00e886e5cfef6908b2916c1190f19d292763e4f8d6d1e99fb06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5c62f0bb80dc49b54c68688d53408961a1e4fb74c443e64dc05b70779a1f8cafa5298a3f34cd22696670b34e15e1035d8b94c45df5af9cb17e30eff02e83ca20ac53cb80a1d2e69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3111eb5286f06739ae3add4a5ee71438ff26a3e9b85e710a5b7979c27396ce70a609f4015b27349e159d87795ef7b30cb688be15fb5bbb67dd2f27296f571a264cbc3313c4af1ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf591f9e6723ed9c4557257ca2614066c83f7166d7b2e3d1b80f0255b1826a59a7bc9c9f5089b38ab326e4d5ed0638e34ba18863f2c4c2814f162eac4273fa9c68d38b044cc1eeea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fff48cc40fe75469529f7f1acd020553f743824e514dcadc082172eba0a4e93a88e69d0b85a5a1300920ebf48b0a5262cc8e9d3ab6cd5c10d590f088f268bef7cec97dfccf377f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9771ce9a4d6ce69b96ac28160bece9e24ec0d05b958f56de2a15a125e8ffe968e6145dc68350b6f8f107e7c68118aa89cf69820d09ae0cc29a65674fd7f98e01164a321e85587d83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b87d9bdb4aa30aac673d242edd0e5315f7f68e4d9df2526b2812826f1e57e47757e1071c70868e986be6079993302dd94dadf12e914807d039bbb6bbfbef59fddbfa6e987c5b4e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha78755aee51d81912cedf612485132abee3afa5ef870d10dcb4fd668ed66b9adec0b159844226cd03335858173f116e22e22b1a52c6ef2aa01d42ecc66e796c23f6d7a4c8c24e781;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2339715211257259e333b57fc21ed4e92f383b5f8aa203be4467587f1f0db1bffabca83b1b05e9b6b0289e3c49ecbbf43e811117576c1665cc778ba1e3a3fef799ec770a1888c7c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97723fae937cdf634d935021247f674a5d34c2607723c5f8b6a72b86286cac93bb86b2edde864c5a9935379d6ebf7a6a856531d0a22130e3b226d6850b969375643a1369bb39dcbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c572c47cfa725f97912e89598e691f6297a49b769cf44db8712fd1607e61c83d6f38adef85074d42bea58db0bbe56d2f9287d309b4586bd0376797fcd63f3e35df80eebc257cf81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce945ba37901f90d3d0282e911fb1885c4a9b77fb7b350a1e9f1b9c4b66be155c4aef81de38e7688367522f32023130aa0a36b5b29cc30c1cf07599011e6123837134cc4b04c32c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha892148a8d458ac75c60506dde746dcb6a10817a400692a79907d1edabe3b4c460402c2901ff6e169f9096a94c4239d4fde499d9332512d27808126bceb1c1f96631564c0a9becb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4cf190b0e596dda55c877761e91788cc01c8207b10842f68e357b1ce41f334958d39695cf2aca4ae72988c0ed136c6f22c33d14bc32d1072c0ac6331a8a65ac1b849e827343525a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb427d7d0f7d1ff6af20bf17bf7cf35b8f1cb772a638b6f9af8a6a033079bf2a3f9a94d5f0ff6a8f49039dda0138f9bdbb0b5e16e6f4845bcfb8c8ccb6e02bfab04bc8da3962dea29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8c5da9b084e2557ef05df047e278963a273e7a0fd4dfd1f273f86ae6198da688e5d2b83cfe3e9887ed7a55dc7518b4d20a253bd11ff75b22835338712e3adbe91c8b5fe1ae53ea4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ab721709b773a4b550ef3f9f233d0e9f6e05031176476a8655add1ae49ea108bac7a05faf804cbfbc29a582abf368dae6500fe959256f0658537fbe118671e63c4292b6d25b77d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedaabc8bf6748e3d45fefe0c52c775868cde96a61e3829d630fc433f16685bb254b3116fa77b208536686472993466233af51c670eb569d98451d8ec1c5d29a546a7c640ee283ad9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f5f9c5c6e7b1995ed7c73e53942f6e7d1831eac2413d10277336deac148ba6f4c41f195cb3a89987d2cd82b6d3bd25ead7464ae8308296f2bfd2dabcea87767fb7b2478cc7135ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6e858d74cb37335248cbd089219ad439c2045ff92d39858a2a4f7285134b8152ec54b1b2b7aee8844323d086bc1b1c5f90eedc482aaccd6a9168181dc2f533d86459bdd4b68c1ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0d48b7fa50a43f6689d23bd952c957fb300fe4fbcf0b68180b222e6d8336b396fcf4acbf5ea9b7ad251d445abebee13f3d6d93d9d5a3766561206692789ae7ce901b2c24b8ebc25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4e9809adc732f8a2e9a203e9c2c192409ab3fd4f10fdcced3f671d60e3a26d194402d34e5c89ed257eafccd9eb2aa67ecc4e3f5102d3a88635456f91d30938810b1dc4a91ff82b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2b88276da55b42ff8963f31362ca2697804db151f68b8ab5cdea7b826bb822b74c7af6532c9fc6f0863b69329f2ffff41e987bc50eb91bfaa7239a2e0094014e33b4e1ee94537e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a34afa37503a08956fe80b91b0143eab7a9bababe6c6b97f0ef6052b46fd616b9a6a240db3a29a3bc9ce2fb3f1cb171e64fbf947cba1488d32dbd447dc8ae2e8f7613027e488161;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9de284abe9d236bf3842068878d23fe08bf9e4964156a4c38d3071b25a413cc5962bf31476cf4b78d0e821d91b2f7fcbd6423412f2915399c73ab69180a068047c7657f5a0651b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1be18cd248a4f07d90a387ea656de4a6024796e0c7edd8110ed0dd0dd5a8bfba89ce232a6e0d60fd90e890f680e6ce1c32028bafccc2f958c38953673415d2fd52bbf82fcedda0f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha941c514ee45ddb02b2d5c11a52477fe737070ce372ff1021b82813eaa7e679e19855e761cfc39f14b89add7ebd4a6d987604af1d2b8610fec4ff49ba8fdb67d390dedd38b383ae5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85e05b92cd2e6ad58513a4656c3c92eca9aa7a6149a6cf96ec13d8b8d75281e29c849771c15925f763920181cb91d8de3f151ff344eb48c612dbbc5162a3a66baa9f19438f8ef5f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f6fb3e61907f081ac9efb19ee6ec21ec67c46f93951ff058894b79cae55725100154fa3530ff3dac097bb22863d5bb21a9385d2c31cbb357a577d2d0fbc177e6b2aefd89c7ba858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h519dd97ccb8e5e50826b2857cfd5bc1896e7199dc5d335f023f5349ce3111c66fb539b7cc308af252e59bd31458243f9927d16c364a4cf408468236d678f02df41566d88777dd3d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8efa7566d7c9ad1adff9e6306179bec87a1367cb9f04745e93600f212a453754601412a439f765e8581897aff16fac2c4152af7166997f2c9ee5b948c1dbef2cd9f8114376811bc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23596c64d84070403ebf0d300716ec638baff023458e1aeed686a5ca658736f2102ab431576a99dcfc49658e6eb3da75869b733c9523d868af47051f33dd598ed373899d851e6926;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h685270a89d1111dc0e4931ee6af28b801b251d441eacadd391039894728232dbf2ec5e3ab75fab043c7a40fb6b3e6d977cd32ea20f40e387e2bac30c84db5bb9c1e1f65bf1fc8e86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82f83e83a5057546a9f1d73144b0090c6ca93ba26137c8840cdf6198affc15603e49f230aede7ef8db91f5f904216c302550611cf7d1f54597b81976672fb7b7fffdee9089ffa1ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fcaacc66909f6f08b7b358fa0ca32535b87c54d5005b26e1fc9fff6ee903117b99005774fae333663210b8a75ae0f232bfac214137c6db635043837226a1739bdfca342500b770d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f518078bcf9e4bc0294c4fcc819c48f8225f128f602a0615e94ceb5248344dadf63b71c40368d6f2448276622550325052c7699ee90d49aa30ac51bfdd448c38d4343558e6ec699;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha60d57181047d521534364b747e0583ad2dbf9a7abc203d1b57dc7604946457150b5820a1d9a24328dc0da0a5102c87c0419661f35082beef72d095a505f2d99c10adc32b2ce2035;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8571499be5cc431a94c41206c149201b70d27c1c8754c1b8285f9e81ab5f65954d75bd469c687f26967ad92a42f1232b0869079258c4053f1f38c2b88f3ff93bbdd26a9469e4912;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5f8bcecaa1a57dfd77273f6a679a6b81798514be53738a6d706cb74e2c4df8a0bae2a30d66ff38d9a94112f46bb658a6169a24d5363626827bc4768a94a06a308fc1069a2128b5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e47029c62037b525f63a8d3a067801ef9f3a632789a178083bbb78e35d6053126e6f7f8da4f0f563724fabfb91a1d393566278fc75c2238144ae6383689f81898a33b01ad73b44f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h780591a82e559724b898137c92ad1804942cbd2e98c1965153f701282c5d0b890d67d88cc9d9192b8da2938d36919c8dd84aaf955409faa5de65559371d708f63bea95edc95086c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4114df774fd257dcb027406063ba48ef801179bcb27d6fd252db152932461ca0213725356144b0c6c8dde623e6bc0cb6eb414dc1c89d99a6bdde13b5b2dab035903c7c3b5b981a0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he92ec37363ca92c378b54a130c1eb6dd390ba3b406e902b04b56765de30583b6c4845a650dfde23fcd55ab607f76b29c18d720fa9662e51e6a92a3654f2545435e4459d9260658a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd45baaa20dea4009162e47c5bfa6e94c19c70c250747c7c40f0b512e6f19a88e13a97de10bcede866cb89e9f45fd442eaccfc4518a69e4f4dc78ff8bf9d720b73e547297b99d2cea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6feb9f7b8b715de2f8d7309db4869a4576702dc84704f5ef9f8d40dc60cde98536b35103140a37a5751142c6d4816041c1d2261bad6eda2f110c7ded2a6233d07061da0e971b544;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebe3d6f51871612ffc5e3f0cd6f56414c4be0a7e8603e723660c0aa82ee2bed8ef8ec5813e8cb1fe514d2b643a551f6871fca3dd1b7893b05f2e1e7bfc9b360d035e7c4e1fb9d417;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8db2dc18a561496c85ba7ba9f74659d69cd5c1d8c831039c56dd13e7b14525cf74d598a85572ae6284a1a085d79db99aac6d41e3c51de916ed71f3cea251ea4474e37fb3435657c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7f40aaf216c310b571f7d5b8337a78640e8b68726d72c417fb9e4abf6267f7a31cd718a1dd0cc116250652f327a981275f2220e5d313bbb73f540fdc8e4e2fdba77e4a9b9354b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1c4e6a754834b65aeb1ca4c383825f678fbca1175974f95561f9d71ac55db4d84c3803b851b00afe08f0a6942c8351e251967a09c0a378d9e00048206ff0524ce9459b68b2c8855;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d1c61d64cb29823a4c08310977989ec82432220b0d393f464c08e7a6d7fd614ad0ed5a50249ef8c4dc5397dc872a74df61e5af3dfdafbb737cef444098c162d5f4c566c29c62b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1ce24f5579cc01350ca48c105bf7eb42daf2ac975ec0126fc4762adc59bc98abb11b2716a572e6fb1798d17dc20fd303a7a6eadbc58562274f3b104d9a59417eb058f0abd66c377;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha77f5ae471fc2964621e9d95cc377bb3210789d4ab0e569f920304c059aa8fa3b12595cebc4bdd517333427d1ed2328966f325b412fb854021a0beed7f3e6ea27482e781cab163a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cd2e854ed938a74ecadb272195316369a6a10f3c1088d9367158cabf4649b851aa682c9d0483cef77a70110f6920bc4e58f49a993526eaa2c2395c4c4d7b94a05cd4845232e1ae7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb28f8ba6b2d995da715b59b83ca670474122269d5be7fef2f634c884209828158bef4ce7b62492355caa6b9eee9b254ade10d1f5fbcece77feeaaa81b87b906bd0424efba74bd1b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c4adb176cd3912350d2ef8ed58b4e203aa1f09af9fc650efe12cdeb7b4d55ac98313eebcd7d72035bbdaebde6ed2a5383f60a85317e29a94d3f67ec48b69a317ffcf99641e0e50a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6979f988f2824f172a7611534a024b53b5d15ca42300115c2885cef0a8fc2034c3c149ab3bcc3a98278c3fd86ca858bdfe2f8367e44d4de15539d0ce2564256a59ea6e108afae18e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h832f14944826369325101261e64ad4fba51964873aa2d3ce657ec1f5a0e467f09e8ff124a04988ccf7a95b78d2eca74de4cbba965b96ccd600511b42240bdab6f46bc6da64c763af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h711eafb8e0fc17608cfca194b4dacacf5dd72fa77585ef0d5bb06c133c84f5593958672f7892ce64e98e3052e4161aa4cfb3f4958c1b488640628ab1115886c89f44982981b224e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ccd1591b727cbe860143781e960a0598b7659d8a23f2a433db3375602a52567938b2f1c7b1052ddf14f20a2aff05f59b92d6dc4a8e5b7f5f5c688fae1a5110d2dc039d4e6c98860;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd78ed6fb2885d4cccd9361613477059f002000577acf5cad612586d26ce9f9d830e3e29bd5fda8a502aadd451842df9bc0fad2e6a17826a10b0af450cf31a5803c8133e50a99feff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a95f762f7eab3c3dd087c904405f23313819dbda478178c65eaa5035f0953d1fb7f92ae29c0b2118c604b7de4abcf432c23624439b2516543d379546e05c4fbd0d62b7810eaa458;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf19369af25776cbc6c9952e05b315f2b44a263be7472e8118a5072e1a3b58caa9f4e252d3837b3636030e7a8f51ea140f78473b8c1340aa261bf4fd6f92559198dc4db50ac72e3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e219e11932caea0f98b1eeaf8d5e2cd89a0c9eafbd1495b04fca81f176ff88246c9bf0e008ae7326fac056d37cf60c9698a3552ea69b19bc6123306b8ad17b8315d0d3d38c80a4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2801ffa0183eb07cbd1fd5d4662efbb940035ede9e8b1e7c4e7e79c222fa47274d249a87e7206ab87b204e7840480e26934369d949d5336720c3c02334994f868f0b4898f4e0196;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70970aec5def90bd427f0bf85db5195314137f2287cf848fc3ec298e0311954b4ddf607b3eaf9bc3560b04010964d8d9a9b26c3c972514d83a959ee5523985669d84040bfb333f17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98667b07d234f47eb1516e53e5a894751a664dfe34885119fbb8dab7908876a5f345da865dff650f031c7f5825b1077f998e9d470e3dc0d9917b10305b77e52460a39fbb6f573458;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5863edb995188c1322bde2cf42111e8f90e6767dfe79d91101a184323e9e5fab21af61c25d6945f129059681d0aafc561f0fd81348d6eef8a485d11a2fd058361ceed36e078405e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ca1ee982e584dbca62249003005e7c6b9f3f29179895c89fee264370b2e1ea6db720149b8aa43816ae8bbfe07842ac5b864a8c230e58c624b9e805fc7c179fbfb925bf7c9208801;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6830a73f4b73aeab16998ff2876876541bb5ebaf3d1fa72f0bb76b91116f0bbd9a4ee918e20809e91960aa27d0dd2d73b3616b2e3f7852ff1f5f2d1c5e8d014d57de6d532c4a543a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5184c15d9eb015d0c0b14f3bed552c504b3155b08f1a6c62abf74b95e26c1986fba08db7a7b8de536ad81b60be753328228092da998e40d4c20a1c73e3db59420244984562c654a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf56e7c5ee0991079dffe6f9db631a5711875d1a49a1e8e64871b192fd6a80a4e93a955842d700f710615e269ee5433ae2b27ee594cff4df4c71ab010d55835434d83484b1b8ec0a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e48ab7db72d0fadd38bc12aa4aa903cfc729de2cbe96f914c41652ed1f082e2285f434c7f8d2b18a3e28d4628f7810c77e131aab93d36d5373e1ea9a82809eff265c7aa0ae651e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cf650ad2b57293d0c6101e435658fd3bc6b07c502b0eeae67462f65837cc66f37639d7818e93c96b0e644e5a57bc0e7993f137dc301ad1dc2d47a2147eb37e9821f470e8c69039f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a5552bbf383ef99f747f2fb3e4926e2971b65d08757f32135b0394567f7fa7b1a899344ae4b792892220cf765548e3fb4befe7493e2a06f00ec12587ec86b517926b6453a640125;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf1b2344018d22eef770099dbf5826f26d7bf7f30c69504d3ef5f6bc10c1d0557490ab2cfd9b1e6d3ad488eb9837d9f2814306254824e4c640d4952fc03d0cf9869007a539853901;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b35e1a3c65a67034da96690dfa7b43e352e118e034185def323557954fe52e44d00a8827e85d654a62c3eec9959fec772fcdf9d148b1db0bf3a9eaf02ea20c5b44c794771890212;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9dba8c5dacc726a0e9bbdf8c474b4c5544f2c0eb8725fcef0ba219b943b87749916efc92b3f83f9b97267028bd30e5b8ce1b126db7e3979ac5f18a5a3313cc5b3d6c81be12f6bd1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4debc6e20e0f950c0de8b75c3ec89305acd47eb6e584f6bf8f4674bc63dbd2443f890442a7d9be6e8ae806ff4223c61c383ddc1360476f00a8b9f70782a70baef58e5b4909f3fee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4b05aa9533290a825dd3439013920e860b2a02d10d46b07bceaf4ade9acf1bb7567ef04d5527f7c1faf7b944b775d38130e956765a1c7525f74c82e36faba83fa68292925a4a5cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4846cc25665768c2e808c8fc3189b2d8a0be17b57c9ec02cd2030ce615b27467bc6a8cc512516a9105d1291ff56cc7403f13abe20b10191e5e9821ff8307c9ba0df4ae498af4a907;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab1151d8bf6224a3fe82cbb6103a0234ee517433b5a586b1b643813bc134b9f6e9e1430bee7cb6c40fa44611fdc8cd28181c85533acb1d1ee3e1c61b856c4dbebc0d3829a803911e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e45d886f2d7d30239779300dec62de013e15b47ce1229b31f198a71b753847ae6c4eb39a18b760b34f4c1460c1c4b9c5340ccc6374a85d189d6830218a8fac24a02cb6cc28427e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1583ded81ec4ea7e3c3f4acf40fa6c1a257a07a32b60015d4701525c5ead4778b8718622eae77b94f94ea80f8550999b31fc0d40f027477804f973ca8f9b82c8e0086c54364e544;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d7af7370cb857ab448431530635ef2196be5ec8d453949b0aafa0b032a1226f6ec2aee9b33412016a9b0d2e74e01a69178f06a70d6238a194c3c72043cbefd6efc6796af64c2710;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb02f92f4119b73ea0aa81c165f5d315fe94f4bbec6f3b16aba5f21cae29fa9f16b015bb0e23bb0619957ff445b213b9c15e2346a712c2bf76d3a9f08678cd752f23ec967c667595;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1273454fe4ca8235cbdd5e188b61acb1a0e0ed5b05f7e79b52d7bc61653182a22058332e729d42c7b60a283e8d2aca9daca7c4303abc6c8cf65f862ee64c4e3ca8138a30e41e0463;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b523dc7198dff02550140f1faa65e2a0c3177fd767ba4a31f554248abe4cee743acbb2c542df8eb416826f8b6f26e29a9eef508abf47b6490563f5ed8918f0581110682e9b4f23e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd7779446d6a734236e6f20eadf1e0036ab3b15a9112fe6ec6865e7d671cb3a21783d56ed9cc98fcf28fa773bc54d73a4a388584a80c25b05a6ad9b0ff6f90c2bd602ba3c074ecb2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h702e94b645d70456821de09149eb8ca542dc8cee9e1b54addfae2ebb4b31ca85a6e63155780082692242db8a24756db35e1664754f44ff0549ebd2953e892601fb8d03f99f54371b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3076d508fe45afb7e7c0675b06b5c0f3b3bcefcb7dae616d61b45bc1e8f70231d6e72241f20a44656fe193fdbe5ce6f80bd9bea6c8bcb53eba52a432cad9ad116c18e1ca31875d1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bfc391fe6633e9e28f3ee231eb41dece9ca26938e99e8081812fb60b99c4cac9e1a527da404a7ad8db2ae4ca3ca97eab1c877efdfa10d1b75868f77615bb8d9ad8552cd40709325;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h230e7b3e3056649a9a2da0201cec383d868aec3191b94c27d2b4e7478b6d3aac986a14ac5a90a564f63f7d5757f9d8deaacefe555ae45eebc9697265e51aa389d6f292ae6895816d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h201f526b3813c2b972ba47d77e0e64be209f67379fbd8698b6f8332eb66a92c14ac13d5ff2fcf9f1b8d968e8f9fba962fc0f8c0e57ab25125aa6101039461525c9472948337ea802;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefaa860bb9f4e29e4f882d698616820be6ed370d97a265dc87545745979900eb95d1f6fa1a4ead7fac4ddc872219d5447440a19a6a36b99f75bce113138a9d639c7ec57c79bbf945;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h752e976973c646f79782a2a3f2aa6bce91f8208b5e4522ef74d1e9beeeacaad19f99eb08569d62116052a382bc36256cc195acbe21cf832c682b7bce5f7a0a655387833747f53057;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h624ab9eac6b838d7e072ee5299cbfc0502f8ecc5432a9954b2d9239418246d2a4e4e122a4267668f6dfe6919e89cc9bb027edc1d5fe9813760535bcaa8c9066cf98b46131255f96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbf7da2b7aa09bfe13668691ca6d9061c463110526291ca33e0ff7a1cadf5f72dc02f4f9659cd8ad9f019cdfa56c2d896c9090f5f7d47b454bff77c514982af8220780b9471327e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf39372d2e9979bf4a5719de4894d4297e55690523635c1d1735ed614523abd3f8509d40c2851d6478ef17369496d2aa6b5382e25a323a90b5137d5f4e1c810f623bd96b3dbb7fc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b250e4e3c19d989d3f466d59a6ed2f9ee4b5951efe12cdbefdb316a0e9282844c7debc71158c338b8c3e053872008dd701d2c4f5c33b771e1185c75890388afb37bac59a729d58e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba7a85d3c097e293a15857d325344628203fd338b2c6a2f9642146bf34a7b7176ddcbf2b259655139f00818f617b8c6bea995a5252f9171395a7f0c487b4ff3b39d9c08840630420;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e8e94e28a710f5a16af99ffb547e67ef3546688d596b37f6f28150a57e52154487ab734dff3d2e0e397c988321afe2fd1d1f2f421ccd9078184aa0e837bd20510b38c94b3cefb72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafc1349b580ebd2f0bf390ec000f1a5878c7e4b4f4892be337e8ac4349ca5125112527bf0a95dfdf4ad3e3891d5227dd8f641bbcd8ebc00f59e0f4a844e94ebe06cfe177d7cd5348;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4e5a4e910d90a1ccf839d958d20613aaeeec41264bfd8452c3447ad83037cc7c4cca8809eb2d0b532121deb28b8cb9449f52a6a9334c01e11e3c809cfaac8e681abac0c747b5b7d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ce1c3c13d226fa91e0724318a360759174568d0dd3a7f37b6fa868b48b93986418190b023ba4c1663a7fc4ad96c90e009fbbfcda4274110689402f00e00f4965672f70607cb1330;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd64373f61020ceb5490a94b22f9bdfe4b7ad33fddd932610e2c335f9a89ffd96a6494d2d9300bdc4bec94e26fc6e3ea8ef3556c042abfa1962a284e965eba80bec1db9c2bc015a72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e0fe0fd0398c492dccca85bee3fa4eb32fa0c8bc1daa5666fc35af686d8be1f8167e4c1b3885d8bb621306e72562ab7eee298846b8b44a320307507eddc68065797458238238548;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8bc32000597dfc7a5cb13dab3388542659104376f1f9264ba5e9a13229890661bcf6afe923a774b8ebbc8dba95e2e42dad6b8678ffac64b073343861b7ca0ecf3edecdc3d7df0bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h442b4bb737437b763a01643c35c229c478233d058ceff2c5256c99cdeebc27d1114d7e9552f8f53f3c670601254ee618efbb3463246dd762d63d47b364248ebf27839f63055dfc04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb24cfa7e8f3d9f300c98cf4161f94afbd3caa215ac543916518f73b3e5f406cc0f0ffdec0278d184585e9d00018c85b8c5b6518c762f7577f65541e11a2ba5f261c1e787c4b03902;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e831208df2854167e8b6ded442d666dfcacaf64fbadff8eacf93bb105730918f1a5f4fb99a18230d70a85ff7f9df0bcf447d1918350c7217174fe63ed409cbfcfb9d006dae776d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h586f2adc825ba356b5497dfe03bf3573fb1e25c42ba6120bd3a8ae39180c79734d05062dac80585f284f41ec0b2d48185ac9586b60ada8f366b5fbd75a33c5f039637cd8ea8dbf77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10b8567e777d222f0032f6d56c0d8d44de4274a411738c076588fd32a01ad269666da80ca0b090a8691d2a7dd8cce7e0c0c85cd42f9f9d24d9678291835c175a801612c21a1ec48b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf239732490cdbfecf84622632fc958ce8baae2f722f7199a3780d27da6bbe0262086d978396233133a56d874652b560d820c0094156868101b908c22c0a833029ccc73c564c76f41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fcb6a9f441db3c1ee720dca96e7d7593cca8052fdfe08b374ab3ca502cf2917e43914727adb4b6613400605c143eca8ab91915bee9b2a967816ab159865fbaac5e9199a371c81a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6133052328f878f5f7936cae16e4c8214f96ea71c6b3afb34f832ab920e7fadaabbb9003237e87570c15a0d1bad9ee01d66a43e7f869da7f798fa3efd17ec86558fab6ea27507c9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2573eec204d0f8e3c68890b33f691872f6b2175026ccc3a37056fe03f4cd63a0effc644a8c223927480abf47b5fa12e9eecf6718ca2854b65d02b8950e079e485667a56ced867d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8087a49803e44fac74b2bec515be3cd645239a26429f1b280a3293f6c570fee0124ce865a3e3354ebc79b43bfa28fe6d1e2684abeacf52b2eba3461e883adf3d49b88bbc5a5b4614;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5807b4107384b1f5741de828a327791822e65f898818c3a9cb2ed55258367459403e1d15dca48627c5e7982abfda3bcc41d272a5ee03cf06edb41ca41f368d04ea500955c34c5a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dc9219975f0738e9eb2cdf3f864dc32c913df24fa1285c39017caafa641595dc71eebdef161ba56ef9dd3ff96f50e246e3c8012f7cc5cd35fb41473090ffb6f68e723e3e03969f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5c77bed095ad0ee58caa5be3dee213ecc92b80c1211482fdee3177bd39f83b951156d014b5677f36e14ad03281d9aed87bbd00d808376f75ccd9b141d6ca7b6357f37075b14df84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc32af64502ae4d645f26cc6bc56f3562c07c03194d972d20a47bd71c680c169cbf7127565661f62d33c0f83a844bfea60222823033ce022c0c936fbbb8bdb4e98c5c798d9f0d6dc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd999eab8bbae04883225251475941924efcbd3df2823b2741343502fa551742f9453d972744d4d9739216a21300e7c215d05f112f31f08c4251f6fa8ae02cb51eb0944d1a4e17402;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68024acdf8435ad507fd528e13f386075868eba161c6939d15756899232ae87c2e2d477f60b3478b1781ef87956300bd7af76d27ab5a65bc9deab10c7558cf81fa313afcae44a89a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a558aa11a233cc0ee463565cd0dc715dcc68240f933540378687cf22a7a04f27f61d6c5fed2e5ebae27dbe377a6fecdfd496258f3843d834d06f5a32dd910a022f1cd188849bf5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd686b3d573ab0d03687af112e9bbe936fa60884698da7fa579c36605b0b19abe2b436203dcd5393eda6386768f2e84d8ef1fb140cf88f9fbc49ed58b160491fd6f44feafb70df25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc353b2d4b73237576b95beeb5006bc087b0105a7e8db860891d52709b4cb53f60d8308a311a0a26002c7588fc4e97679210852493ba34f89fc98acc33349da978cf446d9a20f08d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83518015c6555c0168ddb1de09b0c7df19cfc474002e8c505c034a5927077cd4e85eb115c4de58364beae499bf3ecba7bcad5cd1f1ce0331981642b099f043f3ae3f79b9983d234b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff4011c5063d640552f8e4f623647e9ed2b9fdb8d4c237bd755194fde036fe9ebe7f795763691a9ca98b13565a1f71c4b005f3384e3dcb2c6acd0f454e8bc1d4c604ebce2bcecdcf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3b347c856a3e9436d2080f2575e4cd7e0b9e12ea13228e6e385e230b5891cd8845db2e9b3984c7b47d0010d491a25fc6fce82f6c3f5514dd832018e206049ee46566cb768cadedd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd53b63dfc2968619250375c0028e7292c07dacb394444346fe6ca106c522ea64454d13668f835460c9398acbb37a344c8204269946de15532a4087217eda1a77b477ea3349ae35f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a13bcee25cccc37fa5483ee49260bb161b09af41045deb2e242f3b10cf1129442c46c0070441ee309b5fdbc799eeff4a927ebb1e6e2ca6f7231ce6773383f55b3f92046d8fd8be1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd97ae239ef3a2defe9cfd2711d60b0cbf5ef2cd129fa2c1880f81d4c9200e35e234bf6f710e78bff162135f5c6a05999bfab3daaf1de2405e8cbe6338d0526dc4770034c354d1ac1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf3d251a3646c8694798e3faabc50ea4755246fc9124689aa9242b122cd240b668478d3c7974b03073cce711e5064f07e277a94168c278d240534c53f5a92a13e8c790d35530adcc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ffd61ee2f28630c60ba0910a2e7002da738f31baa04497590d08edf02b5bd31b8338323ef106a161cd2defd08975e206def3b9c38d3e3e2a3b65a8f64b003e9675d6b7266c44792;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h200aa5606d13da14d24315c4f282d32c31d58e9af9b4ca9c79901a09eec8064af05005b12c7c8c965f5315bf41a107a586c8f1bb84c93175b2f212311fed00e827115a920c9e118d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h912a2870ec337a86e7cd030033a75b57d738c4504ca63fa2247ef025069e330859366a6ac561ab59caa59c7a0e204cfcd25b730fff2c06af7d2959a7c4375b921f464dde0ff02cd4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed0c473f608b1eccfeb28b2e363e357554931e675e0497756ae78842a61189c5ab7c1858b297f541dedca6bd52e345d043820b1f0c4966f14789a335e6e936924f8fc12d1a59e542;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf7214a6bc1e55e9e8d0c17cb69161543d3e4458967acf597eb6ac0244c687585548fc63e0a2d3a24b8577caacfe1b286a4b997aa9391f0c5e7ddf8878cf8d793f45d75d4900aa5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52229bbc61452ffb2e752adc70852e181e23df9dfe5fe2efa222860b1025656adbfbb29bdf2b7274888ff8935de1dab8ccc8d22a1bb185c1e558acb0ae7245b08a5b99637de9f953;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef94fab4ec5c78d72f65426277c9835f1a7e4c87c39573e1143d8795a526aa95ce2b61c21b56067961f106550a47ff1359d9f3bc098e603324bd84a5230df0b9c10d05e416d46521;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h295cba1f2c45d5af4a86e56c831ac0759b87d6cfe548f488524c5f7611bfcc17676001fbcd64d1b3fbbf3f3e99cd004e52719bd617b466332ac9a76311633342495d198fa02b14bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec51b541ac7873bb449f6272102c48ea8bc254d9c974b7a5a8e72c6e4b40d197c53f9ba0d8e00409166a8f130ed32b8b171afe9c296ae1c4e0d3d1704b11198a20e0ff7bf290eee5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4c99ec5a04f5484521c50f0bf28f3d549093fd1770910024b681f9a8a6b9e78a9174ac7a69569cfe4103a0c0e4d981ad026606071f88608ef541dc78caefbc8664c068f03aa9d05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h780684ebd81ee977bdcee88be5302e918b0a56d868a9590886675f552a0d76aa87d8642d1b801a1660a5b435c766fd4aeacbb7f547009a4ab26382e1446a19fd09a11fd2468c031e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee4e937ad3fda9496591a173335ce1dcdcc1b67572db14599c0fff92c07899093e17e244f817d952d5821f57d73aed9e5a7a7f9b719e42b49c20a4cdf4423d9c9f2c4a3e5ba5e0f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61523fe0fe50e14a7dbc66e6dd0ae7c1ed2a5e8c37d1a4a6e75df9c95310b29cc154f050fc98df7e7311502b6888e8bd998bcae76c09b9ea6669396adee858de0dec74b72dda422a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bd3757c062f1f6dfdbbb73a924929bb13cfcf9b8a9be174e58ed5e459713139ea4e8b221a96e31a8e2fed006698396333be9ead0280bae405efa3d08d2f2c8e28a0c5b9d58be262;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h827cae63e06ffe3b16042352018b341b7599612b3651e4ec71ccdc9343eeb5c2cc280ec8c43559c4c59125edd7c361b37bd36f943e8908694b7329068eca7f4bd0b2f13e3690bf79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5012b840d0cf2035dce31f0a7896c507c0dfcea0e8bd69c94573ead0eb3c5ea92fad5e68c508f1024d1710bfad745e3bf68abbf00ecf5e86e62f84d000714c548171e470e3ecfbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbcec11ca21181fd7b4cbb05e5ef5a96ebf864197608d3a93ea313e14e4331e2ee25a5f4ea142fbf069055a6c5fe130132720c2c4ed0318e7ae71a28554c4c527a450d110bdade02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h678186aaae0ed43251a91982bbfa20991c1e55b96cad71cd54502a380490d8825e99fb12fbab9cd1dbd18b2639b9327a43fc7eba3bd5388d7233473e173181169dc49278ef202f83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90baf3a8f28b63d09d95bed19e0728c8cac16c56e41d749c532de5720e7edf480490b9787a24dfa3daf75f41e14a6bf2ec4f6d5f44ff21faa632ed49574741996aad6aba1db99104;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb69d9eb5b4afe57859a57667d3bc651e449d0fa81c3c4b6603e3706968f62b755587e89400da60f4a2a83df8bd24edff766cb7eda5ced1f174e279dea535aa99ca56089ac4a72e7f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he60b7dee104b0a73b1fc1cbd1d60542fa4a58d3b107ada12e4570a8274f3226b5ba2f0e402bfbc9a73699326813ec3bbc24f499961c6a9b5d0647147861480cc8aa69e864ea07743;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11d4fb484bda5ca792fcb526daad5928c7e476d5b3fc65b4f2dda8d2bb1b53dcd5d14a2e792cbf4fe80f7175ceb90277f7b864199bc45bc2f577979a481b03247ba91c6dc5bcd13c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce53d2328c680aaf480d3b2c616eb452edcc3a90837d726874f47cf693acd1a62afe3591a79dd283ba44d952f4acb3f1b72990803217140ec8b2d2079d39816f14423aa95191b8c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h229569adcba51dee9493744476da0bc2d888f79527dcf61790f9d74ae2255ee6a292981ee74db8420d81c332018b8068783ce041580730206b8d777975c6ff7fb14f64435526d04c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5673385d9ac29261c05449beb5356c40d8f2b094bce69074b4846ea299e10a78617ee06c836b4adf5824aa1d33e4d506889507cde23549c09407791c313989794ab8d06b8409b07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59e414be6f612c285a5f059494ece3d959417517aeb9ad717aab3a05b74bd9408ece03ef666e0cb828e0799c260de7827eea42d0514c7c2ddc35384973bbb849c5f3f68aa1cc66ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2276b7b4853694eb8b40c37ae6d39f2c3aece473bdd4da9f29f12f8d128196dea0694e9cd0158c2c232033e27083ead65948b252425427cd1d434710d211648c2655ad231ad160e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52ec3ac0b62ebfb9a446d000a2b62d6b891f9958c81a09b5ff4cd342f0eabe8895004586c75b8de6128f83dd7b87c707407b87f54ab5ea7e580a007f9cdb268a987088aa877af5a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had972774cfe0a99c90ab6df9a28ad29647889dba9041f1947a5e0e574190f6d966961da7d69ee5955c12721cfea7e83569ee7d5f1e2691ce1706b71dbd4c7db48e4721919d54a1ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc708638d3b1a2bf395967099c39558a490e1f462f28dfed1449f56ce477e3084f826a830104fe61fd8d788fb465296648273b82227285cc234a7c69cfdb8a56be8bd62e8cd0e4927;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a0cad5590f258fef6e3676e8952e4b3334820ed445227c1a708a30f7eee283897fa7b78db601d675ff9390f3888fd0897496c6668619b8543827a25f02a97b293c01e94acd337d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85c557682025acbe40b09013b785dd4b2107bb9511279d003a54d9b5457360318860b49ff915734078597991bddfad7d660f41a4a2e60ac7ac97b24ec5441e2327a0df2716804434;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77cb768bfdd7eb52b6f73db5743369e7124fe074df4c1955280b8ab6acf2c144e485604d3d8f7b832ff4c6399dc005965348d3b55af1e7787282989648c232661b937bf2bff4ee5f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bb22469d8090bd41010d65306489bdd979bf2309b134e539ccf77859d3a6fb63085bdbc15428c34aaa3a3fc9cb922c6f4c2c7ec908117fcd0475c71d78eba7666a3b9b4d930ccbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h982fd02f6d5423c0d8c3fd09bbf43e6ec98fb28ed559db0e063ab978a54598f135da757c41ef1bddc21c7b7e8e1e155fbad42afdf1b10c9178d9faacad9b26a28417af9182170d79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec0551a4069f1297e813645b80b84c3d1f4ba748c568288ae37ee58f5ec70eb071318f5a6d4e5e076efaaa94e5838cf5e5942153025ed1125df13bc6829c9c0d7834eb43f5678ba6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47e74778aab5882d563bc99f1ba019adbdd4a9ee99d63cd176ff16d05982cb4b466142682966476a03467a7df5110d34277b2bb235277070992bf7660b296640c66017c6cb66ea3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14263a916b6e86e4524adc746eb4d5ea2348abf78b207a15b36011bde4648eb7256661d6cb9fd875a50d187ca34db006ffad20962cc78f2b406cda81638108d3ad04c63e5da5648f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2492b1168eef2b57b36e1dcfc0af4d09646854dc8393328c91d6681f6345ead05ddf263041c983d94f993228ea0cb794850783ca0f546394419b89dd0a6a87336591baf54ee37f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb6800398e1b26145d228f23cc373d856f37aacc03c303ef87bbe629bf3df48a601b321d6e949466593bf939aa9539a8b4bddfaed3a791dff2a89dbc7fa64c9fdd6d6138b46a79b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e7f90f512727192116fb706f67d4a24aa609380520600db1bf69590652c8ff279a0caac88ad10e83c739e42656965aaaa4cea760ce28329fcd51f55109f25a209ccb7fc2903025;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d91d75da1485cbd2f769979ce8e9892d9408baf867518893fe189fe86cf01617837c39de73e5b6863d097d28ade45b2c1f28470d1f5f67f361e8f957a4a3479baee4882d4e0b80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40d9550babdb283e680bc7fe003a8e639b1fc736a72feac999c4f154a4ca847772fa79da251ddee74ad62d8efde7280c8567c583d978c62a5285f7a70c234757fa431c669df33cc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc0afbdc1846404e291cab94803c4a693a282c7b40ebaf2e2d17e9a9a857649f9d5dad87b79894a1c3146cb53bcb64ef6537ee9898b364da66d5f5105bd54d346dd6ad3cdedcb923;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19545de8642b9ba3fce3ce45eb10580330c0284535797fe8e5ffbd6b73454b8a4e22a1f78fa167a1e3974f133e165893fed7ea6c133f439f7a911b5a2123657970de1dbc9720ff33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1669f2d749711b4cb7fdc580a2b10e05ee4207d4b4f62a7563170d55ef7cfcae9153ad758dd8487312465112903b3e6ce8bc9b0fcb996f834e1d11c8e37782a6dcac5b83da9ca333;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfe30997190cfa0730225de2ddcf6b4bef3d391a832991c81bd1e5064477d04bfdc9dffd81a8d89f827d3807d4ac4853e66e144152a5d5e875e116d710704de22c78d9900610a858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99bb75c9cb5851f24de630b4d82b54c80bb1e6348c98fb51a4660b2af319af5cd50811d94f98b15c2963591daa3d8c35c82c07f169c8612d25cdde6bd455d021d5b09f51b20cbe27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc83e97fd817972cd6e5810d4519e2352b49a17fe03176de30f1d03cf38fe8a51e17512b99e85b93db7ae94eb6a0175330e1b9feaa212735bc1e8ceec1d3a186121471273c8f08de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf62a6776404a80daf208ea9efc302be211d1c4efeda766d3a058cf2c6cdbf8cdc4515194953f04e943c014e5050c6b6b072361bc2a65521bef572564589e72f687502ea04277781;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b97a9ba7510a16ccba64a993c0dadab89e5e42c880856ef8b38da0a02f009be20716b6eaa35f0fc0ed833853fef65702e000ec9dd3016c431a2784614f5f72af22d8dc08dd6084d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7105724e915578a5341563b3d1e5099c553f13d2004f75c28a7f7c194471d90eeb7292948d5642f0561cd882e398ba814db909bafc8ce15da4af1a2fcb3c043756d1bdd41b118a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3542f556f77f6fb37f1df06b7342e00da4a11524337f021e810c4242f6db6725a227aa8c993530fe1646c9df4dc0c8e2887ddc5e3c2e535ae71000d9636949d8aed8ec0dc9ebbc43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8b58930bccdd75a6ea8359a58ed4ee5481e0ce6e21ba407ee82be14483bd2e2da2131f051b5f437c1620c780838d947fd54ca2def7b120226a7208512dde027069f4ce53a6606e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf659fb7fd359b49736301b1be9101e809a8d2d3a2d7a2a1e20564a8d7d742fa7b1684b0d661590bfd099ac348a05484d36c82703e989ad7bdfca89f1af8163729a4717779b997010;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cbe543e887a4f15128b07cc77f1c7ccfe031ed3bbb99ea2bc31647396d189fc66714b6eb3f00e058b60137500f8f4cc0d23b51284f6472044a9ece306c06ca9d38bb2a48a8fe59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h454bdcc46633dd3658ae8d4ca835d4f7269a16a391330f4a70631318f12bd4d0fbf024fdf8d7ab52b989ef20d7eb89d53a30074330d25706658631449060a1e43c8dc1d577605eab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9f7b296690bd1757dbe04fcbdc9011f8184b288834ba72b1fd877b5512e0b9bbc365fbe334d955a3b8d8f9eb8c51364d5648ec8a8517d3172883e9ccff2518cd5e8fdf149d16b78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7f031475d38dae4061753e92829c9e1414b20f28e91522a595ba637606ce5134717516ace9d64089fd6bf7474619a326ecfc77baed681665c645d95c90660a9c2e406b484fc4125;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1461543256153e20dd190ecf1aebb2da1ce1be5d8101f30933aa51f8ca40f910a35974fbd227a75afebf30ee523ee193347c85f0a0a0e5c6a0983d791a47319adbfea1e8ef604eda;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20e0ecf50b8d68f101c8b525e3ad12ddd3dec11c36168947effa7d5230e59fd149bca5a0405acb13cca65c346ca6bc290f83bb47aeeec432432d6d86937e41a00a69a5fc3f0cf017;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h504327a4781920d499df3740bc0a8177f4e9065967ddf15f7b8e668dedd4bfe9b7ea58fc05abd321cf2fa911a2ad334a1d3c9f56c943e84f505c13835c31aeaf24a06df665e99344;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2b9d0da1e83851f09c733c5b05867825c6c850ff76c129edfa8f886a227c11232d006fe7b519659a803804844b5717b75d56a16ca13a636e43dcdd18fc9bc28ea1e8a9c6bd03c6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8ee8af0485495d6827f64d82a098edc63c788216f5f595689f771f572b3ebf04c6f31bdb7bf09cb03540238344a7a875ede3c879b7432eee9a2e3d2124023dd4787f665c23f6f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he966b71c200cd5802527702a74b13d442828b1c3429a80518e5c33ae5595ff51336760eb91c5d26ac355f81db16d4b505d8747f398a7a6acc2a67988f500adb7d21b4f164770de81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0b2bd6f8f2dfc33a0806c74364aace638a332683b93433592416ceb5d655fb40e0fa57fa6dde1e3a809af21221a70923fc2f64da0ab57525c2f0ef8396933526561d44a217afcf9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h383d8087db13d947e9f5c62488ae5c417511fa57e2e4b32eddbe65d84477eddbfd6fc7135ad19110862020d53b970b835aed39c800fc40f35ece07a0f68fcda816f7f53d39c8576e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbaed31fd91104f3ca61d98416b7320f0002843dd6048cc994eb672c38e8fee4f0c79806075fbd31ca181dbdee3a82f9d111dca170041f36c83639d7a8b02c39261f9f09d340d5db8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f1988a6d8c92aa66f1a2be6352197ad279fce648ecef279234fef4db044cb800de4739341db0e91058fe50e3a1a71cb562cdefe36fddf6200d23a1ff99eaf55775f0a467d64396a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ca2dff120db380d0b1086bb507550b6180eebd2b4a3940703410ba7a34758b0957b95563d13e335e61e962d57c867f208a5bb0e12be45c55c3fd42104c7391f3b4b592a23291ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h432b241e70624c6af03e839be26f412cb83a05bf278ed44020cae618cc1cfc4cbcad8c3b9da6e5b4dee235ee7db637ab06c69b750da7cf94cfa36068f854cdf1a91ffafe371fefe4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74f0f8eda4c34872047746855a332c9844a0cbe92ee263c70dd78b6cd87d53d0d949bf7eacd2ba35b23a25c703ed2cb39606d95751683881b5f4004f53b47c5189e691150353b060;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfb69b575ce4b1d3a715f226b0e6fe82a0a915ad6b61b9feab6df3fa77659826a883832d92bc147eb0ca9ddce1f1e66f628bd1feb63f649a37c80b9aef706c7cdce593c1f6efb310;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2aa314f5973216197b7ecf02331fffd86fd0ca928f5ca43b38762527994dd2297b8d55e826b627ff0895a758f4f906885a3cfeee202b000974c7100ac19d73692519b36e2e29e07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef0adeacf6df33d3dc75be5898f92adb2162b891e58ca6f42577aa9ae6f1e0c2938d9e04662507db9b8b49bd6f89b4f520ed3ee7342f22aa5cc81fb9ef3f57a081b02c556777b620;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h488b136c2b98064e45ac404a9b87e0eba7d5a3273379ac0930206b2bafeae6ea8fc3f73dc67e9cd01a436946d7b174219dcc2ec1cb38a15e124478be0db962f7beca9bfbb8ad0892;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h682e4953100c96bb0aef574baaef7152defc58dab52c2ea1d7a368e93042fd5393ef39b58029c63617026c09176b0ad2e13b2b970b7ded13c000591d28089fb82a2a9b6fb28cbaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he25c8571be7d117ba215035d75ad2a4e66dce73636f1e41ca9d581e1240ef297f7d2d6d71a4d4bb54bf82033d435ace48c18f6ae0ea0d59a591a897720748f19a3ded0ef7aa47555;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7174dc8a45ca4789d965478b72b79a956b76c3633da8bd309dc39de784f82ba4e82c25c74c51489214ef669d86eb0f7e05c7a3eab386ea8e8157144b6e377a8c9b8ad7079a4b455a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2f610cf4c2fcdfc3da26eeab1de1fa2e58557066ceffd45fbae9b5071bfb663a270977caef7c6424141308975862f77e353d4ec7bdfa6360deef76ab9a3eb3a12db8bc2321b273d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd186b077ca3df65583586a9a82ac1d63c6848ed3b217eda0888bf9ea89f4750b8c030a12e2951499182cb909cf88e5a54a6b2a853aadee4b4d34ce1f71169109863fde58788b267d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8060b5e88334722ebe6ed6bd47dc9570f3c2dca5533e3abc6054d636992dca50aa2b0b71f0578abe6788e3802ca5a2e08af40f8057ba71bf55dc6932e1f83f26b85bdbbc363f21;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d3478bfd895d36750e78a4a4f1b471fe9101ee5ad1e5add952041ee0d70ec4b716b09a776439ce6514c9d405629570f06d4fae1194ad02dc90fa0fea4b2864618013e19e3184d8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99c477b04bd9c613934ea8067dd8e5a13f07106a697269c4fd6f29d927d82d1d3bed11948681f67add684ecfc62056b4433f22dfc90aa6a50a2adbd7541da7b604ba9380f8ee0dac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec3abc9bdd0e312268e4d67e8c124b481f6d5473b65a17d343173a4a2be9249d21d94aa236380fc1d83740c683fb31ca26a565f1fd043de8d15306a85fa76eeb07db3903ea50d0b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d22784f7c07afaaf5a2d1c3a5748e0b6ea81871f5b4d8e8dc1781bc61b7a78d4a8f5b281218dc3e47f029750a773149984d9c5a5f216d352aec9e87f017e3420dcee1df7ab83c47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cfc0f3a1d3b44a0ac2d82ed4332dd7cee15a0f2fa9d44a80d1dd2b5bc6ea0b327da4a969034428450b7033496911f59aabbfb0ea67c812c67043d16a699c7a6828db8c606df673e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8575ce39b82409e98abdcc8e59d7e22f79d366cce7be1a8da59238b8083efbd71266249f2ac46c42f6b226111b705a38e4a008934d30107f9e64cc12f2bca4d764c190c1eee15d6a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae20d9af2d1c73d30f653252149b6db01c7a2af9f2f25ea979937520515afb8e9ef873f90f49833fe0721add90ab1ca683eaec25d38d077f8545fa23984b769c5ccec5d53b3a2d4c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a3a37a62b2bfe6dfb26ffc15ba9fbba091aa8993d8aabb73bf54bdad3fda525f00f09751496c0c1e4a91bf0caa47ccf89f8c139c45820f9df722abc94e48112a72b2d1e5139bfdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb5c759c9d2fa8a56065f1c3872df16d2048c32433f14655c215eefce6e624f37cad9e120e326b38a0a1778caa9a02ffa828f50f09c2aecedaabf66126065fe5ac8c1c4945f417a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h698a0fd9c6c4b8fa32541bdbc5b77d9cb46fadef737de284ebf273ae74affab27ef4b787706ff02c9a1e8ec8040c6ff3f15acee2437156e2c621648d640ae5bc277212467561a181;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf95fc5cff7794e5dccc41db57d639220ea750b033b572710ca90f796fad8e6d7eb9202580b4c224e4bd76359ba624224fbc832988cfcff9b701846c63e45749d97a9b90478fb165d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9301222612ea2d42d64f74878c014b8ef55e1143eccb294cce259b35d36b4ebfb2a8ebe6590beb67bb6a7e4fe696863326ac0fccc3b0392eea3ec61c47778ce6257e519d9ce69b27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32717a524fa096e87e56a7692479c687502f6885c4a4f5da50bb8472727ac620a95c6810cae764d3c3ba1e4290beba61381862d71962206bcb3da582922b90c912c534348a837e73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9178b057b079a63571692c30b8606bf291e8867f0d0df1b891425f2a81034a5b63f5f89707ae2c33a348c4d77168ab582ab339ca6411a82a559dc9fcc26a9d9065f5f82d928fff72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92f5011f1d5a6fc9ff8b61dc226aa357aaa313de33f9a65248dce07fe7f8edd11c67707ed28cc87dd38a92991def183338594a2ac429fb199c1c1ce200be7c45cb5a0c249de9ee73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf511434dbc978bcc0b5c0bd22eaa9b676b52c6e959ef9d8fe04bd441854fb1c0f42bd84196bcb3bbfae735a3f33383b9a3d4ee6330a16afada3e9dead0f1f8f28da58f6ead5874f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb799226a7267d21bf5fb275236796d5f9038f97b7608753ca6027b2b793beb65c401661c0a690786c70c72f0335081ca7caffaac0cef65a9103c28e6da40bc8443b667495a4e0730;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb810c3b4ceffffc9499d37f078754611537de42f803f78801318eaec4b004b4fa3ed27d9358e886bd96aaf9dd7a651ab9dc2e9ebd2878910a6cd31ebc69ab3d11de193f4b053d26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4827bc4753046f543756705cfd4dfd14850fd64abc3dba3e806614f73b3a9ba293ba92688a035d9a81517246accc16e10e0aa42ceea506a0e6ea46a51fdc82ccc2e18f3a7d55357;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ca4461d6f49a19aa30d991ee4a120d03d30f0c20c60eafbfd6d3e2bd39415cf29c88b700bac460ea20b034097cb2479a5cd0777f15b383669f3cc6b3c92d82ba73d6d88186a4d9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11d3700b05fc8b68cfcb1b192651f1e67e187f40a934d67195dcf304302b1edfd9ea68c458e38161e563e830b75e16070a780fc7317d4d654a1def8f629ddbe87c60670b5ff7b493;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6997fe56ab13c10726fab3d995d61c60b40f1287dd4f56736fc05142c85a841ebd7b69b70ed903f3702b437a8588d128f48cef022f9983c9df49939a070ca66db0992f22e561d990;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5152e8317389816fb3d5d126913937991eddf3b6cdfdce86b71b48fc971e8c353d9c56441b44f671585b88c95b15d1e70bebb3a87f74304509cbc9501f37fdc23f3cd19394ad2e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h184483307974d5c246e057de926920c10e4346c8f7c0d397f2357f2047f2455d7e655340a4912a4b0d2e27b00aeff75ee9a718363fa33c2d150226251a2d37b7cd595427464eec3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfa347be771002e55898127f43a400c666525bade463eabdbd2c53df5a7f21a1860b8561c48b8fcf75f392749b49dddd04716bc3f1e476bd780fb50edc6bf1f3aa37e88cca02295;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he499104c0c9ec6d9caedeefabd6943eadf144dcb844fade0ee2cae9f5fb662299fb5a96a835f583dfe5c6b831af744c7b5b48652311b4780a3a9bbd97538a527619f43be9676f793;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ef27bde6c668385fcdddef0bafc452262e25cbd1186af8294ea7493d7912599aed74ced90b06ba5ee007d803ca156fea7e9d38d79d828c5c8267d5d8dc3c376330f93eea5fd9f68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd9cfa0c7a935fca06a89b12004b01494f378405ab4cf7a0d919fab95fbf545bd603345f0cdd1c7f26e667beb1c2ac2311330d3ad956acde40eaa9434189d721020d2c76e4ca3540;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5882c288e1a324d7c9694e6f6fbfe2391f87b413b7f710f99b6cf3ccc9e2db4669a633a6527d2ccf2d21d623274ec3351a67e630a7b09d3116f7b3c4a06207be20a158e7e0f404e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2154a8d636704951940749db342126c08720876cfa0b398b913dcaa509e8129a398da998fa556d6698991c1ec32bc549ca41b9aad1446d79ef965714cd549424cdf8a9b9e0feb97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65a75f8c87ef0c6fc5f6b2002bd9cf99be17db27ebf9ac41a22e3332e68100c7111fdcbaf79b49e2ae35d7b9c2e585b83df055e3e8c8694bce5643ee9fdfdbccdd3215d5674cdefe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21bade187370e280fda4d3030c5beef4675aa6d93cf9603128efca6550b25fb0ed30a2e6ef8b7c6c3b34824ccc38de856fc15c62c4cf89beb10186175eef37af989810743204602;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29b88655b46274e4a5414ff15ace034b3803476a2bd8f43f2c292cfad94c62e1c7720a2d564a95f24fd9b6c07ff3704b1e5127f85bc717e46393fb8452ad1d032432c5a59c72e53e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44b41d1b69ef907788d525f064eb9576c6402e800ce9a2409f819ef2a8f78a43b8d1d4f01ccd3723048c18e694cbbf45745b397e54c9e75cc9ed1eb6f9308b3a35ec91de7b32d9ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde3c9b9065f5f420796359c24ec7358b19a6cfeeb6bca7c9b0585bf7c59ec3eb9f6dc9681962c7266904b27706e2fcd8312e3cd44907e53312c63e8481b24fba10177e48963a2091;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49cf9706d1345cc015701bd5097d25f1bbe91bdb2e6305eab4c8137786d8390ad6f9d1adbbe18135ed7ac0dfc50bd5a0ca465bdf0731be590dda95032c969521b65364303dfc894e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde041902d76645340512f026cbbf8cd3b4274eb24bdbcb5335926cde449d4c20eb596ae3838c9e38267ef82858e6dfbf869e914ec8297a9a469d8349858ac7e381def9783bacee00;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28b400b5249859229e8101c3bff8c253c0e85996faa25eed821d9e4eefa1e79835908070818b211c8d156e818aec2c12d1165a5ddbad42517edc6e7780daf39d5bfeafdbba9eea9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bb0c8e367024ef5ad92b239f77767fb258c408b9bcf7f30052c73ef44549241a7c32c316bd2e68c5fa7a143e1907d7af7e5d701def6066e5fd339df6bb6e40396e87cea2848d93c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81b85b4174df8177585c80961962b602cd65206e6f7326dc52eefc30293eafdf437b1f3ae656ca4b94d68f66ad056ee21c0b45a7b906fcbb01f91faf6f7446d5f6a42ae161c42178;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9fa7b18d89e731815f3d1e053cb4ff6f67ff73ebe30c5aac8d7e46abd697bf7f4f7772b6562e264708eba408a1ca1905a2d268b446fa5aeca2e4e582d08eaf79765583e2d435150;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h197fab0868fd2b487093e67aec6cd826899c24be61aa66b6fa259589a7860f51106964e5a94f6c42af82a7267bac3f01e9e2f4b01a5b2fc0ad6935d6f917bfe3ebc957399a2ef327;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2390b51fd2549781bb9fc0fa47c590faabd12cd40f1846380ac8fb4fbcda8a8edc9d31d34a99131464b4bcb960209884f4a277c081c980fc3ec33363d5efaa5b6e1ddd3c176856c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26e0437a10511fc057d52d1c3c2170ca7e1a78224b171e0f3d90d55bbb9fc3e967d4d064c8a63ea31d42e55144b94c8aba0f8fddbcbcc309e7c5df8c401047f24cfed0e6fb99cf3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e5236d81fd2c6fed6568384a95ec906b76ae64219c260354b7a1af98f5aa900ff0f9893ef801bffdb08e9f8320deb139eb3c3ca3763cb1a32f39cb2fec0b90d9688e74bb4d3fe37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0bffd1603c139b74c45a6363c1cef140ecd52540e1aeffea9bc823122e8c7e6fab9482aed0191f2c9edf11995402c77f1aa06ec365e0284241ffce2707348e4f4e8e38388e3bd02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f4eaf76086fab18513dfb1bed4b7dfc1bdd0c6e24bb593ff18670bfac454f34c2e019e938800d8bbb23f669950412918c818160c1183357a8ce058ca6e7f3d5d8a7422deaf5cacc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0fbc79c06f7208cb8aaad5bcfb09fe8fef8c2e3639d153bb7550239cd6e68e6940d1ca135eddfa8b554f870956621638de779f591c485538a1c64801f3b3515dc5446a972b7073a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heab0b388095724268c67b6ea4cc1e6e94b6df0c8dd3f66bc093c8c2f23671e2967d2b516cf40bb2928cd439d7de190531090a4fb9528d844d0b56aa6f457f2d2c3f2c370f308a903;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4671ea54318da9031f96cba90085117f6d115796c280fc9c3815857d684b49e5bf8fab18c2b8606a14487ee668061046a4a400bf6c133fabb7db7ab2cb7973646cdf19cc7e475302;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f150d60bd73bd908dd75014666f565fa37be8e625248ea2c38d332d115f243f987339c2ed2369603946f9f0e48e2f3563a1938543fc3707339bdd403b17f700c0e002e948fe9e25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4013a9047d50639e8c4952d55767478650d5f87626f037cc8bb815d9b572e9c8a00abc336d35d593fbc611fade10e27e1ceddc1bd68fd1c9301ac2df03c98938db736c2ac39237e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d7eaaba67e3cd5332f5ae6effd8b5bb26d21b771869e61b8888ccbec5d18c1dbc046f3930ef356964eaab225d32e91bada71089a7d0ad32c865869703ed4bb4a0061c28fc64d78e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8f30a9db0d121b4f4dd64f5be2b145c46be69cf2c3db94310838fa3e1ec48b8aff50b55c5b068d7475ea98d90c03bf36d70cc0a1ca1a6d3f230193a3dff0162c951f6d8db37847a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29ed6b72f0439f926241f6bba17046644502b16d290873588fa47946137a9e3cd823024389a35e7fce31240dac179d61d9dd7bd8fb7c411b668b456182484be211087fb7216e4839;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h493909841d4c1b75eb24c56f10f68942bf51fab03a30e283a9f6568aa67877d9b5b5c441523531ecbe11a5e7c7c972475bdd4ffd8f46563c6806b3ffd673ad36b3bf9cf005816190;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaa76d447eace591a31b72bfc4f070fbbe126a8d4bd48007953177391fd71569f9ac89c733bc5694f41d194683d4b880de971659634a3d2b4a11828b4221addd81cdc9db4407934e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ce9bfc3011e175fa0c5f06cadf68c047f6b31ed46c79964871d0e8844f61323ee746be402f0e95ed869d1a797f0e1bb219656b9b1a9271420f032425289512ea7f3fab3b5231b32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5af3db903976bf646b4aeb968ce8f18057edb9663e5311ed06453ebcf5801ca6b88edcb9af22e4e0a3e9c55fe4913e5d6e1d28583ab73e1b69632b7f0c225bb14b3f8beeddab22f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb541db52c14418b181d656396ea5d341f7be4b603ba1fd85c49074ae57ebf50f578067ca9bfc5f2e3778df671d9e84290d5096c06ba0186884ead26448c17abbe50830af48d39e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee66c016a3bf8204d370719d91b4a701d560680166e2bb12c7fd4a70a0b85842cb30da5693179a4675151a7a59dab1c1730137f4c82633a5a853ec4fbd1f4cfa203a31ff91578160;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fd2fcb5a3b1c82f38ec2aba256229ed12219994b5b1a811ceeba31f454bf7ea96a922ab32b018c4fe457106cfa5e911703aa0bc55b36ccea70d360fbdfb685fced7f67ce6ddf232;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29310cda8658c6231dd292697fd1db2f06c738293c0d9855ecd723e2ee79a35ae0176c94b32d335c3c2ea53c1846c30b54133b1116bc24908f1bd4c39f5695a7fe6a239b0549a059;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7c1eb9501c4209c7800dd6162a849dc901fa2008187139d417dd3de856f5720a1d84075e5e5439545eee3f30a977e7e3ec3f850b0193d7ab1e6cd757474b4b99538bcc9df5bda45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25814d7cf494eb6c8aa4d5c9ba5560a50dc974b90e0366ba6650bab03e124cc0348ee1ff1daef8e7a1abcce1420587906d4d6c4ad7293f1c1eaa0163267624a6e5a85d7a666ffa25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c4cc8f279792de8b7ef40f5c6d800bb9b63f788f10e59c9052493ac0955d74ee25992ecf4b49701ef3cd793bdac49d1bd82cdbb972a73ff999e59ca2c6f81b38ee2db2ba3bdcbd4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf43f0c7bc62f50efffcea5cbc24fc024f98da5b4947a18a14a0424975a3e33fcd581eed90c60c0f5f06427b4d536648171e320eac7be82ebbbb5f9fb7cf5186cc6f785aa054a56f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26e65e14db6eeb59924f851f4838278ca8711b8e8279c38df6e0672fa0a32df3073d9c230df38c6ba827ca4eeb9b50c4a72f0845155c174097f5a8256e3528c2f624890a3d202393;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b36b8d23a0e0ad2f2aae9eef140994c0c15697ccab874d6f4db7b20793e06b11b2fdd565337bc6bf67b1f518dc41c4ceb9fdf032470c58d0152e69aea72302b413716bb6a68add3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97712befae42649b123dc69469f7fd749d2758a74dba63b67c42b239fe53001c120b61f2272784ae62f420bf73865982bf648723389acc0ecbca6a82ce15df0f51949adbbe92af41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ffdaead3894e2c813fff7256dfcedd326c0f67c354d0124bab99d78e237c73c6bef6f0f011c60870d807f4eb3af4d5e52fe6e1c5e6619c534ad9ab15c3dc3d412da2858938028f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc500f420dace6fd82867456707704a38d8d7c421f82a8ebfbf9ffaa1d3c7484f8c7c84caaa997264ccef341c44a9e95b922f7002e57cdda6f591740da7ecb3c7996d51bfeceeb36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h857dc6ad212ee5e4c8cdf36155e9415342bbd785b35436c48be349740f8a0c5df8f12e70048aad948a0d610d68f6bb9f16eca687866c81b24cb375c3ac2f254589724d52660a3e4c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d51e4447e77f6df314dbd6400ec3c75fc403886aefc6c7b03a68f2dad9b40a8900bb95fa2e1d1f7f6e97fdf3e55d0cb472561f4fa6de6a5896743f9b229f5a86cfb85d69a087023;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd01526fd2a30b79719322564ab48ea4d0469b93cc485b78734361d7c358e2872440ddb63528ba7c0f45553696c832b0a11e5c54c98a92fc837b62e7ce79aa288cf01ba58aa0d1c7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf4bb299e6e960a252862358c0bad31a7c4cedd9dcc91d29502c091a3c7e8c3724aef876293d134c00dbcbe8e6ea55c4e9d8ab36ae7e32a4a33b88d84c2c32832bc513227c087472;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfabb859d6b4fb5802823c719fd22d01269e787a91b5511225decb5931cb78475d863a4cfb916bae089c47164bf90ab30e8d2431c0047bec2228a50b072cd8b88a548c72672cd7009;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fdcd3c0cbcbdefaa1cf92fa40434896698cfe75d3418925c6b477f6314ee5c3ac51e1bacdd5b1ed2fd74a4000445f5dc7a3dbdeb3a89901bf94fe46c2798a9f41068484640f1c94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf02211226313944495c829b58e7b3fa5bf2ad9079571b2299b4f680b6d7c05a37f173b71358e94f840afae347e64e2fe86ddbf719eb830d7e3965e82a60ad79a6006c96515ebb036;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41d18c4c9dbef307cc9968c8d8583a92ba83676ee51a762ef8f87d76e341f1cc9d35db7692233032f48314f6e88581e8ca2a5b964e084c9d7a3096932780a0f0531fdb7311ab807e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32ae96a3f97a5e57789231fc0fef346ba9db8037583343b1553ed212684e99da416d7c8ee1b10a521c33feb6be89eebb32750f6473ac2eb2b8326e15577843568774f3f066d3c718;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h799ada2ec43d0eb7f75d62719d7d35e8a99b0dcd411d3cbf080037df11c84c1adfc815c8899aac013e0e3a9e4ab57908594919f8438aac9cd684ed5398fbb39509b1be6856eed2a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cdc42b215474ee5edd6574b83627609f325d2f5c014ebec124b8fef4ea7e9569cfa7b7a5ceabbd04fd89e70b49ae8be9f6c390d1e6b2698441a907cf74d239719c05ca29dfa6c28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he60cb1f56ff72dfeb0173df337e58da1fd38a0efb37439431fa3bd194eaf64f1ebff68291a42ae94121643e07f567e66c4a37a0d36a18706b6469362eb2fa5a4d53d0d92d5d7aa48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h658a442eceba59df3b15fbca779f6b13ee955c345a9420aeb0e7892f2d0ab02b388d155ebed01bc9e51547fc57c50b2ff74b4e96b6b9f25dc3a4cb8ecd1f6a577b305a6eb9ea1709;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cefde78d76af61c8f03cb2431290b537d96003c7e7bd3678447da1a04fee907163e5e4f9d779d1d955c7c0d6129221fd114b3b73c8606bea36ba466e2de479d8c0a4f3e119b7f19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeb90f2c1a3923162e5a193152ca40681a3e310ed914fe891340062687fdb65a2e5e0d7d3ab60359a3a7581ab4bd1ca87a0b7d7d5c63d01f6514a687065f43b6bc20711da59b4652;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haea14a23c5814aa31d91e39dbdd440d1410dab18dd69a59c06a4ff079a0bcac2db0d03963465646bf8240238df36c8365408193dc5bb2f70b16d67eeacb0cbeb707991008ae4c1c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf8faf4f7157edeff97e75b215be55b4d17cba4be3597bb961ecf2260983491c1c47eda5fe7b68cf70ad1cd8bc5fc2100da88c8ba9a6cc7ed2bb962b0d0671415936024815e719ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdf18dfcd8371d4e2da88907711e09d36d3f9e82cace387b7b733d63506768598db630820cbd62a46a7753096e4c89cd68b9d5e1c291b04960409c4596f23bef9119097fe785c297;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3876e895db8c952ee28c9d26acc1cd0725e0e163ddee897bd94d7aa8d5ef61ee74b5a3a26e026ee52f0248823d2b5db82586723ce519984d4a815ef2662f0596b82dc7d2f8ac436;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac938b7bcc9622d11cd935bdc58f00a23a108ed69c4240a73dfb525dfbce30cbfb593803746033bdff03311ca2cb885acb06385b9e36c09a7be027aefe1f5f21b666a36fc40e39d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5b98d4e7352216da1381036f2cbe4c9199dc856216b032e00698c0f6103d9937a2f377fdd3789d602c63394cb2fe6f50a2b69d71ea3a30a298ff6a78fd9e164787e4c6fecff0ccd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef11275e4e33318bf1693526bfb977ad1c4acca2ea48c809bd84ab1539e1026c00790f716ccce0b114fd5313c60f787bb3609f7b9c45f2b7aef8701630188bd3489cbe358c682675;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf07892bed3127b0bf0446f9be1da35f8efcf95334101700c81c86c8e800948e2af6089bb324cf110acc0e8940a13f33ed774bd1371e39d8f281ba4b06bf030e5a4d79c9a47927f9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55578eddaed937d94244bce763ea7a4a95e5cc9c96705a3934f9fa32c2614ee32d593cc0cda366c1138f2a13e4433bd3012a12a083e55989b68557a1624608dca1896b51e8d4b09a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habc4ce97c0b74e510b24ca11bf5df7f17af61ae3c4e2960a72894f41d8f0e1fc45d7128e662a89a2a9fee25b34d0679dab68986a3a6b0c54037939c1e2be5ed799b1e49d82608ee1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a2137df2bfe3d02a1b5dbe0931cafb6a32d306f735fdaf72e91475229920526284c6d7bb8c437d59a720b66e3c122e37ce02350c9edbabac6c2ac69ba876b2b9713f53e18841010;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa66200d19ffac6bb9c2cd417c0ea8ea4c60b25e5ed85ac2c09dfcf040a8fb083b392c426785b67a6a91ea827f0b8dde4bca1081cf6531e826acf72c8b534286aea4b810e2b71246;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaa810614d599f3b04a476cb9646306eb0b37801032e3d4271810dca651805132ee3c115a659e45cbd15faa49d28730fc365cb6fcad5dfe0fe041a445f85ba011fb0f0e4016c3704;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a5542438a1b4165abe55a811d58eb7829281105a24f46ff59160e21c7038ec084e85a08548188246c3de8c85f0928184b0b244759d406e2fdaa5d13471e648636980027cb5a8eb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8bfe657f3b46a9a0b58ff10616992a7b4c9d3229218085631e900ac94b008dd452b033fdd4999aeae7e3e8a4d0852852bc7bbeb0b8466d43376e0a79cfd3df25d45d7e28ab65912;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e4fe01a7974e8ca1a85a692e472b98a4cc4b651d2e0887a819aa2b805c77accf492ec11bc8410c560f117c058a9dcdc8547905709ee1010df5615cd8098526643cc75f0a9aa984;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2215bfe715db72891a802471c29c72408509e4532850c58d7898e92ec11d4cc13b6db37ca750c861a6ee32a5ec964a93c8790418645a6aea6a5a4cc53fa4b9426981ca2c599f93b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d006f6a2df9b1c037836143c37785285a44fddb98986c3aac19aac73be080a7bf10359f88eae94441194dece663386b46949077d16e0c35d9eeaaa7f6d8863d0d78b2a09fbb08fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79cc4e6a720515930afde59619fdba7ce407d751bf7ccb6270c474b8fa4debf3d61f04ea48390889faf4764596d84485d1614d9736302ec045416253e34a4603c7e4fa25b44852e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf34bb96a7da58f667ef821cc379b0a4856a20696b5533196f138ef0788082dfd169a46b71de6ccb45e779ffd2a9636ee6b26102edb0dfa900bacb15995d87b2ecd605625176d420b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he64e0e3c2917658c04c0432be61ffbd13332f80a79e4954812909553be02dcc56925c76bcd0ad929922ecc1520874057560e617fe754762f6f366071f70c4680b848afd73bdbcaba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57a13f5b293d383b24794d5453091c05a08137184b139c041a23952a6e8f06837cd44dfbabf79862db0da2874eeecd1b249b23ebf62f7451239647d4d54f7173fdb740be72132e29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb13ac7796a629825bfc1759e4cf9372d723beb5b0aa724e092380beb28172812fd9e024fbad5f40db1a0d2b9fdb8352196311500a5f27329009940574b689fcdbb6e1fe4bc7590e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9af644c671ac3e76a2ce7f93ae2fde66a9b3ed258b8773312cb43d722fa0a78cc601f62258e6678cb69f2d470c6ee5edb4cd87ba7e1c4cb99901f364c3ac2bc73e25f911a96e9a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h780f28ef2416fd02bf645f509c2471ea642bb4f2270f4e3492be87aec2e87e63d4dfd0eb8f406c8444a1ebd056508e16af5368a9a4b5be49086e7f9fcababd5fc3c13a86e5313309;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf735ce7f5b5456f5d218314d44181101a2e501fb37a5f8f071c834114e227c53cc110b180e0abd2c3a7cfbb474c04e4cc30f7cd630962881eaa49e7d1f95868586166ba9d171f40e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3386f487106316816136e9ff2bfd7173fa0e0d2a0121dee3797b3f901f4918db767c05a42125185263b022b5a636125cb64921c4ca7dba0bdeb6a52f1cb40901ce67ac04e9051cf0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae498fcfa6b8df4f64c0aae8a4d1be6f3f34f3e6859155e4ba99f122d7d762961e6522db53b5ea2b0ccc5f22026bf11384cf324347d012629f3d40485bcef084a2ae6280a30ae7f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h222d71b82628a4785bead8a909667d1355de135afdd6070dc90de0bde2ab6b2ef02523b3db87a70960a28816fa05c258936f34889dbd7e7fd7905f211989dd9c8fa48781fba2ede2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5983455e5827d8441997a984ce50e1b1b0906c816dc7b3663ae409ff94bdda2133cee7588c1c3445de408d8986ca1cfc0a1c74baf703f342663b87402e5dd7f2212430f9a14b20f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9668a9b1e6fb59084a7bc210e445ee24dcff4bf0bebed01c0fb20f67d616af1f8b9fa15a34aad05a72fb03f8a4cc5024abb79e6dd9659b00118d1406a9e412cff783c571034e75b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a6312042f69d8d89d02834374129c46bbecd6cb9859b305ec54c799a642fdaa3b7e5326eaa1aa5b5362def90ab32b410d47499454d8ef973e62617aefdbb4246951f4ba57de687c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63b6d4f3318c726ebae6d1f7f164fe3f17c78e1f10b691dacff502bb5b058d6ee0638b9153434f1198d448fc4faec6636e2bea280595b3d71d450771f6f322db7e022eaf1bf73464;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43630dc6e6e8c3020a6db4ec14c28db83b4b59374e2de1cf5ccf9f7590ca0124b9f9e1200da55f7cc982fcc4c96a9f9eb9caa0671ab90dd657f3ad00cc032a64717eb013c5fe6c92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99be365e486f1931c35cecb6bc5afde233976eda3d2a586afa7d65652fd4d19d475a98969b035265b68696b5ded34b0968e1b04c54cba8cd188399683bf9267f8f7fccc00358a390;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ad7896dd2d42bf8ccbf91391aefe53fd00e9e1455747122dcd86894c68a348d9e416cde0cce847c990f2a82e2eead434b18872e1f22d6ca79413b0af8682f240afb6596b10777fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68c917b9d9182f33618529569d1db93437a1d729f4d9ff3976181a5d75428f42b290673a884e8bb3d74e3cf96127c5a7443ae99f27e8fee7a92ea7cf2e078f9ca774417ad6de11dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha93792bc2f41e9101a6d4376473c2a7b0a31fd63ea61dab8d1d7b8d5e4033b444a05a0812138c06d886470d898971a75a689bb303fac195767511d846f170b7491fa84e33d60f9b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65255dfab0c87a193ae796303bcfda23e118820ce1bbab0240bc9919e4b43c0544f651f8001ceaa813e20e1fbadce9e2ecc4c0dc6427ec9484e7ccf118a130dba47ec8961e5e53c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93a813de0d394940a8316b34f1c26d799227c08a776fcb2d2620bf9e1a0130e1e8349a7c375693b9bc0ac8351cd0fe570115de401a8e4ede4479e77556883d27f4766722c97008eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcff496d7041d0ce432e4d8238c921ea647f55277e9b722d3000750b3c1e984d799bcf1f07758b2c386b918198c72747cdea6f2e10f75a2b102e6e0dfa6d32b254bea3bbe0aa318a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb3fbfbe5bce820369bad4445b3e7c8a298f816eae6a0d345c51b94f6c55f7ad63c3486da353df00080bca58907716487eee172e495939aac31a0ac5a6be36197861fa37d7b4385d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6db161f46a6f921928d91cbcebe0766f7a8bd63a2f66a1651c41a771060d7d4f71f2fd4b60989cfdda84930cf6f2457c99fac7fda41cd1c529ef13567819070db90bb46c081b4051;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed9d63f2db02ac7fa1c1bc42958fa10b62924b43ae9ee40dd5da95eb1df5e6fadb66e90c515d07f78fa7a8c1753d9dff33c4930758d9937af15e962867de830a0dd9a56b89e6d12f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68686cc40e42959d0e79e30078d9427a2940592ee304ca9334b4a8420a925489852575f2a01c5195178263c81c263145b2114ce8e549d53eeaecc2d5e46380a37a0b9c17d145677a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heebd509d36bad5f354be24441b0f1dc5c38f0340d6e2120d45a05273641b24eaf2d87f081004be97b40c2fbe1cf2a92f1302eadf344054e02137d9bfc79b78919ed9860803cf644;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96f0fa404abd835bf10bf739ec5087061b4f9be51e9a800928915febc108640ab455133cf90c24af8dde426bedb9fe0811fb053371861a3d8b5e7092694bf16edd23c1af946cfba5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9115cb80d0503273a68eb41af4abc9c2eb2c197316112399d658edc24bdc5b70310b1314b4bdcfe70120c42ba36485aa2ab01265f04ee82e9d41e2d909ab9d98b0bd77d3b71fc27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75b84c20e5178d6fdb58702b0392b6c9d45511fba7ba528cc219bd1dbd9391cfc65bb3e408d20c67cfc69a30451a23f6634e1ceb8f8e09760c44c78940e0551c4107be51525fe57a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7ff353f53f5da0304c5b57d9651dab6ddaabf9d72e314333dc1abf29deb1c3b312d47fb6f47ebf4cf949ca5a5f60130970cd4b0685713dcddab716d236159334a7dad41b54c065b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57550b66aeb5db44715d93177683f40b2aa1971f156b9e28b580a89342bb30bea789e6245175162f52b6f50b11026bbf41c6702c5e2cd1d363c0b9764f76763de269042f2893e12f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4068f26ecbd2bbc5fe176bb0eecdb2fc0850ac3e871fca023fa9e7040fb485569a7b044e4aac9c8aa62d183e7d702848642a34de69b71dfd2e6e1a6a5e8659a53c7326ef710fe843;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96aa832be8c04216559d15985a58bd7caf56b037932cfb353841e18c298a93e14ad64995f7cb85f24425085a82d5d02e0f9c5f83b7677f3482f96ecbf6d78eba99e8791fd2718fa3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1530f9c5382c97d5c4fea831528ea7d2947a68f272d603f599dab23f5a1a9ea140fb8c7199b767c8e6a8b14f7d6fa2db93a079226b398c250c03a5f346d624daecb853f30247d59e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96af414739ec96a1d7f1d3bedc2279a370eb16ee1e8a84d22012a18c25cdf146dfa70a9f03cb29e05328124c2b883aa0c897bb8e43e8ec17ecd61a4df29eb16f8a098ca67a2ac8fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5065d9a2dde2e8d8057f519787d548bfe3c63ce3b5740fba12ad0d0a90132c8f93ed52c353f54987fcf047c7e2d8d8f8ebdf757b47e8fd9f84e8902d465e3eae757132996c6dcfb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc037a2304e20cf6d31b90907baf6b4a4cc038c2767936eed98d60478f24ec8e704a189c0fe269af7b061788d6fdf98a13b6fcfaa1e2b65909c5187ff4b33cfb1e0cef56f3e7f2fff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1f5d5a0dbf5f5522119a4d59d8458ef151c35037b0f707e41885105bf5f8f00c77fe741eda02ba7fd59cbc1e941206d4112f6a2b8e08672bc12a227a34770725816228dbca4f5c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4442cf14b5ad8e557b031a7425956d0eedbd1e51e0a4e15397b282a6260ccc0863769b234b26bc5bba1e5d4b11c13250fd4f2b896fa981ccdcad6d22ff912985ce67e523b014209;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac05ba820b354bba0a3de76e577779374b14cd102208d766a21b2fdfe4c8991861d89945f801ca2bd1d1e4de55aa52e6b6c9a3976222636a37c8c170fbfbfe370c2f834daeb31b21;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d16b805e5f3442ab3243e37938c5d9d90f93e7d33a691ad0b3983d43a8cd79a5c23249761f66011d581d12536c20fc6fd2b8e648020a554cd9cea870dc845755bb59ec8154cf0bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h622c3a3119548a196b02c2d9d662f41ffe32e54c70012794a8668f8562c6889a296626b85a37b015df7e40def713ba3463acdd2cf284ef810d55b05a51ad1ef2f9060a24d0bc6145;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70d636bc325e79a5dfbbee967ca1ff0dfe7741f74abc27d2d5d240b2a17766e3e15f6e8e057767997ef8a6712886901cd900bf2247f1520e5c40b110ae39a80d89fe4a4d4d6fbcfb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbd35c602db75d5a02c21d00084b4d6bf490db7ec9d218855b88723b9ab9ded72ff68fbab224ab3467d93ccff9550e8a3afbb74234f12d9d84c51bf64b448b2b06193bc90d1c88f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaa6367de5a046f879a918881c886ac99e388f87e1608896a6ca733cfc772fd23185b04e7d95bcac6a186935851c6a13b72b9c881c0199de0f890ea9eba659339fb67cbfd67c7830;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9049fa394eae263f9147346a61824491020e250ccb1efebc4c1a6222cd58e5befdec2ee140f532522b7621a0d84862dfe41560e7e17aba100a46352635199533ef2c6958f0790f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda2e6f6f8443232e2d929ee2728b1064fd2cac1b65202799b0d36628ca9b816504cda52633f810f1dd5e9d3b9cbe570521eef2602ca39f4cfa2a68ba440157d5b36882c57e0b12c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e41acfb0a338d0471d040c74d298568be4ece46efa3e0131d3e1bf950a19b98f8c4b68c4a2aca8125e20c7df2c4e3c4037933c0eebeae3b8c0681c6efbf864f6889ed8530a558de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h303f908c845d078b7f4666529dbe000c1897ad78a9c09516a46b6f8309555f85d98015515f5c9cf387382ec22c4de19d68053f90157cbf0cb2c7f7947d6568e88897130afa61a8f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60912bd9d30937ed372b65ebe29240f7d4be15665d3294bca5514774dfe2798c7d3b8faa631e4961c347dd3f02d126bd454f169f98357935b2e8b045d37acb95a22e9b4ac255b4d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdef97d1a4d4952eeb7bf1cf2f15b8ff9190412aae9a8206f4882ea881f95bbcf4bc985dee1c7bf0f38b9a8166f61fe887805d0d7262fbd344f94f55462773cdbb00e198d68a7e4b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha38e61c7e878116a47b067988d9d51672075e04bb28839edad4b6ca237a78fb70d4f1a0dec0cfa7ca5cbc277dc8251abfff10e07b57fec203a0fa7b47dc12336e988875b5df5bbdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6dce8c1651f23bf38495c0eeb466d6bec53ac97ce56f90dc61d9f8182f85ecc63e43419ef4254634756f26863602ab3e64b065f9c725a09075e2a9ed6b178401ffb3c5bc07a924c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65dc871defb9abba80e58019dfe72a7bd4ecff9cb825baaba069d86b065c935797b89c5944536b68b4d056cfebd2fc4d46ce33ca269584eae7fcac75074e909bee749f2a786b6160;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27e7c5bff99efaf36017f116efb9d4b3f5dc93af51ede9604466aa637dc76a2273808271677f3480cdc502d43e15f4dc057d9bf5b4f7935a7117c8c2d94a7eb7dee862b99e5766c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4af7d579d6d29837a781a0990ebe452de75e6611001fa6c4d18b970cc33a82ee0f755026e4148f6faf48705a86ce52979d4732eb07a927f162ef74b6dd8b4896234bac7c8afde9df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3880103b1d990671a925d07f09a8c9f8820a86f7f4d85ebf6aad04eb32e45fcdb1c6eb194151d09d66ca4203e607e798f0fda870da04e4b25389019b8dd543455cf1d4321501ae92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfad23e708efa02ceda32141f2f3dc18026bb00d092816aed283420788f54f477d028681e413a79b84fda315084e0d94754e4103eb49674280653ba436dbc53184124063cc6b2dc2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4eca32aa5b3745fc5b0e9195b17e32d16dc66bfab9d75194f82ff737ebaebde174bcd9311862d7dc2191167f9f8486f3b30766494363f04f027fc6e1df0656e6a662801602f0751d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc07ee1be2c2244c167411082f0f68fee5b8f0475ea50fce1e0fb156caa77aad2880dfb2122d3760b53c00169c9ec5875262320393c92010a878a5b4dbc869f5cf2d3861635ec0302;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h234d864f6e693d080c43edb9c3dce28ccb53cb8966b573e438209efedd4015e6dfc186979d9fdaa2c18bd0b17ae4dc039f054127b9c5f9afae24aac547f466a3ba33d4e10477c348;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h311078ef29b5afd31cfbc8a764e1c2d840b305d1280e096aa7b45dd524ed072d687ae7d5f9e38e14ba70ce1881bab4666c31f8ca2cc6b3e55e526e39978de291ea173fc126be80e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf31f10286895af225b32d069a525dc75bc9a68113cf7ecd1867d2a049fffaf9797ee306bd229ce3d2b3d39b1756772261e16a8fa9e66d8b6a17c10de2e2f576f1d9a9514b9b6e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7274ec0a19c79ed08a5d82336d436e653d89b13fa5212430bc6c714a8a3f0e810a0d28629dea7f70548085451a92849731a8776e8e52499d0d0a0bdac6e7ef96a70906b8685a34fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94037a5b10df973c0c10e78e027f8c1972ca57ce84b50870a358a93dda994879fa14a4276d9d01184694606f74148a3fc4df676f8037900b7c6fb3bad6f0c357fa88d3013c927598;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5cb6d99f66d5397f1272e6a34ad21f475a71549a3df50cb726734249de068e441ddf2424411233d5f2031c8268201fdddbb4801bdc3144100d86a84dba7b59dd3ca63eb896cfa6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a14d99d72e80bcdbf53a3be0a7fb489aced6cac00f8f7de20dd92e765c115391e90617b32503ab519d2050964604ac1d0fb6e9fa3cc709caa13f9f10aa9fe30f8391cf724da8139;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed1612ac729c66e2012c7bd75cda0b88ea5a7c989eb0388d808f541c3f2b16c664496b54c43f8feb8a18794614aab6f6d7c54cfbbbf72ee0eff3b822edea1217d56925d3be288e73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9fa0396cacaf47db2c7fee3629f05086f62688baf76fd5ad0b4ba117bde0ec682dcee32496be97d1d0b36b3db5f42f9f4d6592daa1a5043e4a98e39e35ff5a9b8a51de8e9d41774;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7190b2d03510f2bd9026f4c20543f9fd5e8509c5b46170657f4b8e739d78703d6f42ee25addb727520b19a642da92bb07745aa9f36b51840dd2e1fc02e0602fbfaaf2e1d0e978c82;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd0cb58b2fc238ba0bd2bfb9df79f92e00b96ab5f7a8e2d1d3acece58b1b7f32b38b2cdf8ca47c3dca65de144921070c4993c7cf740b96ee60eab1113f71b4233e5ee69c71de4272;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23a881d05cdda43e262a5b7650e148d2ac3aa41dcf0d82290ed186fca2062ee295a51c462f73b5f5131784a33f7ca78cc2b768fabe2d6d4325f45f28a4790cad0284ccbbd2f330a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc2d2150fd951354638e5a5a91befb01ddb7910e923f565e3795a8a6382b13ed95cbc490a34f88f627fecf16185ef98db7708c17e50dd9a5ff8126f772f80c04b7f048214621acb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h129ffd1b1645b94fc103623664fa620b0ba7ea9faf56fa6b23980e48f7946bb93b7b676d7bd18e0b0cd03a3ad0c1f42657bc1099ff48e9555841f7104b049155377fcd709eb8cfb1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6566b529bc2a45c8388625b2e7d6925404267ee1a74ea7c13ad784daae722cbb04eebc4988ec41b11ae5814029775799fd62d2c6893948c1e5920c7a1f3282a4086134374a966e1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha602613519ebefbcc1b56b2399b053b8fd3447bd17c1e69cbc32dd04064e9cdafbba6a11c96e1842b853a2e3d6b3f064c7b63afff53e7a09521b095736b4d7312a8f598d3ca45fc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h128b530e40e0ad9cc4e002976b159a894da6de11d187190eb5136dd158e54c79fd11fb3106f615f4042bad14d6f6dccf23717137a141b315251d9cb95c53e70cabee98bfcfd16da1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ee5021d875468fe29cc099bb5138a2bc44c722dd7065947efe2edb63a86f2c6cf75725325647fdc84e1e6b937ccdd0267e20252f368592f3ceeb5a70fdc066ad32b49f6cb320fa1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7d04185743d40862c4703d6efd81a08ce11c7ac245b421583326874d6fd672dbaf5c2b091ac12b145d4617da354ea7d54cfe5190c9077f6e2c3de4396d6cb70bb21a2b0f7b831f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h577ac28f57e6b4100c6ed773931ea35ac496a5d1443b25307b0dcfd023a1336834aefa24cce226164a6b4a1060aca5fef07f010bc11054e89ec0da74f707910c9939dbfcfa314b26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3445f0a3ab49c70d697960649b2c4c965a73f340d5f011bebc0a0ca779befe499c2dbc0bf66fe8b69a63443ed4f66dbb50664430cd8881944b1aab0bcdee5a4873ef17468e8c6e79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93d6a9d95574131dd34a0f796bb1895707f0a6cb75448c629690fb5acdc5aedfc170870579412dd694694b9d774daf7be17f9423cbc84bcb8d1ad9179a427e122ea732f853f52b8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1ac74800ef06565a5f8b5a64bff56ea296f8561d39ee764eda15894b16d0370a4986a4159de1079ae09fe324997e5824b6205c7dc15cef988a6ac99c634d58aa6f68fa36c1e6910;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb839b2e5cbe66a102b444f46fd15968451932d9dcecf0f745bafc769ea6147165d1c56b088110b6fdfb965eb0b9e03e5b105021881cdc8505ff3c9e5ec251b18d768a1c9b2c76526;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd931d32f5fabeace3050ea032f1744efb2c1d177869743a4c6f87d25613f3c4a7e776766fe0ece3b2b504a23aa97215e9b0f69e5f9c71a6d9a689b1227ff859fc05bc3b53a4a2096;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac81825baf4ea047101d0c702a57bcf978c738a629c3ee9795674ec050eb9fa7687615bcfcf845c324a86097ca1cf263c6fbc6cba5ebc90b097e3e3bee740cdfba67951e3a7c3441;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c7226cfe889276ee0d5511b698dcdd3a3a23bdeada3c9e0a76980c5e6a09655de809cb4442f11c726660c1a9992b49bfd942c0d2e82d900b30df1348a446c34e5f899f8b95229df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d882cf1fb67ec743545d8397ee50a7abdd0d5165f4b959254ee6d37ac4a0a3cf6c95e7b229998fca73d0e853fd466c34f57a0287e4ddc771fa1d619ff64415a2bd526436e6e89ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ec8283f9cee6d4def238552435fb83978fe7f443fc60386ec35306ae4cf2211f8fb27282e6cdc9ceb01aa8983097f3f8185b58605646a7847f1e3c8bace2e89a127bec86533d2b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3becfde100f5b7cb9ee082fdc71245dd2fc0ca95e347bb70b9bc3fb45214267979dd5d4117bfe930483c4c4cc6d061cbb1bba51d3d1bd84df43d7b51968535bca842df6dde30bf25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h206a198c77d283e18f99d7f8b2332123030afddece61f363459aea5d82f0d0fd261f85d4d2956a3fc918fd9ee41946d2eb954d0b2f7c56af743493c538094f5b9c2b33fe10f89e8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4af5932927156703fb7a97310f3999a38a2463bbb0dc782a1483697f446529d83ae6dd841e6291933a2cd4aea2b5641dc9bf6e513a2d98a0d075a93106b5d79c9f2575e66b0e270;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd88e803d2b19f771011a4c9d2f39ff598182b099b919d4720017fcd35c3524945472a2728cf33aa9b334752cb26d3cbf8f9f8ab4c508f45fa4fc84a62a82db19f736b08101272b9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4508b6bdcfe4fe3dfaeb13c2389a5be9890a63df79a59d7bff4defa47265ecb95c2aba74a65ef325ee2192953dee6aa0560420c34d2140192f43659447614d25caed2cedab4c5f98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13fa43c1d1e91c826665702405d56d8cab1c69fb2281f0c707107447abda5eaf9a2384fc9f9b2933e8f342d5e2a9ef1090daba8c3699770a49930f8c7f944ca0135ab4f09039087c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5795814d4d3115566750e0733d7f8f11d38f0bc7432765eb0b6e898b41fa2d05e22d57ddf55693baeb06f0f80184f9c39ae3a488b4f99065428e738fca08db5ce24d52be5f650d10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ae96d42de3656ceae129b6e1a11602c43116664e0f0e518fbbecff02cd86fd20d80755bf0f37d2b9f9911b5b3f7662f92a540e3c2082799f62a613f8c91ffc9149d32b5c153900f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he45b3809d2e19916114625350583e25c6757853f67ffb01b5c4fe56a638cec6a3fbc4217306e0c383ee976a105672a0e15d42f66beeaec7d1e70a2335cb1328d4cee27b17ab3c64d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcff8545daae097ffb3a9ea06b3f94e6da66d65d9bed89a29878181ec00d33e49ba2303cf3cd59934932c14ccaf9d3816f3a93eb680b3b395972faeb049435303abac955edb8a3fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hada509cc63d3f221727a616b97ca34cf41d95f0e043390f14a0fc3ca1c0a4a6b277e935e744ce39527b56f5af5ab0b68d92afb18e355fb68b8bdbd4f8039db5821774f780e2ccfe8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2066cd832c543a6aaded0418bd459ea26691b4528f9e88c054f33dca7dcf9ee28d97df8f6aab235c0fab21e8f07f34fa94517434f9aa572def9fc3ca94c9c9defda675fc2eb9f5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha44b32f7bffdfb38901c437dbaa4503aeba59e315fe138013b36f190b8c900017d01c3b4d9283345a18864ab1e169cc572bbffa5d925908319aee7105e15fe8ec4ff6c5d339b63b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc7ae77155756b02d505c4a20e1eff4f7d147040975552dd3ec94597f70719ab8f224264b9a703be6d1b489bdd3745aa6352b255b6805f6fb3db0b516f9c460ee000c829a54990ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h690d6ac840651372c1978415da1e6550936268ec566c6fbc483ee40fa08af6030390283cacecb5d313a8c76ab2cec65a83602237070a103d92832438cf00d9bbff8895436758c601;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31e1780833feade81c88e1ddad6949632b0695fda846f7b0ea221e0222e69e758582020d5d90c73ce8ebe2e836c9ffb510f355c7fa3e554d5633b6ecb75ea2b5f23567cd4f4b31a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffacd3aedb456a7c5d46eeb159d54c04c10ecc9362c132d4c3be29905ba41cd87d6f833fd172ad202ee37854045f4626c0bd29aa5b1a21970fbd9856c9d5de00d4cf10ce3df5db4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcaccb0d83e6e1b548cfa86788be0358acc3a6fe216de3d165ccacfd8f6889cd9c6be2d791af3e6f4f9f6aa39b77217ceb5d326d8319cef66db56a1b5b5ecf3a909d665a4daf6430;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he987df8c2ce5ec29c36d5e5fd2ced00d390ccfe59d63d9b013e3c2fb1cd5174952e017136f5fa6d0e8d2289a24c56251ee14008b404665d09926f2726b13c653ffefee4ad802770e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84c2bc80bdcc13b733d6ca874fb0a62eee014e905047e1b71923776a5e2295334b38848a04bce3494bc5df57c9054cc479e38a4fab86c7f0400d06d335a38ce14dbe0f360440b576;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda52cddbf7c97d970a332d65cd947216bd733f39beaf9fcee04d31dcceedd3a862fa036de554cb19a30c2891dcd61378a586254829fd0caa9dc06ef54d932674c2ff4c5690e3f8b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h638c338f76d0fb016ca8e4b5a3b15893f6417ce4a4b60935234c1ed95ab574def75207d2b8ae71e8ead21545cb3ac3b73e36673ed7f6e62ba7ecb0615542f37d9ccf30c40d06d69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebe539e55c3ae7a4023bfe69b70931487e453da10b5376a3deb5ad4aace30be73a23e71e97cc0c728c6d296b778865d87a26d9888adc7219a95418cc720cb70f9b4693647aaea23e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73c64b089c79bdc247029b60835d3b1d4b04869ce34fb977e27d445d94ab3fdde96cfd629f853deb1e33f2ff99505cdccba05296a2a7a65764c2fff7b756045bc6fca1422078578a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4d040bcc300efe8a2b9eec7ae5ef3e2174a92286934bac30fa885721888f64f7302e11677a0c33a6b0e7587231afcbb784dc0ca5dd305d5364e1f1f0fc41f8fbcc84a012ea9138a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe75dc35364baf1f9846721c48ae11d44840429d97bd3ae1d1fa5d23265fc42b5ac4b7b626c3e74fae370c97321bbb24b9fd0a06b40491e7e02bd81fcafe114ddb8053e95285ed92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e3ae1f31684802c367bdaff9169d94fbb1558cdbcfd2df440b98b37617fb5ce13ae6464982df2cddc76b8265d6d9c354d01fd18f3923923c3351cf88bf963b45c37c813c1f36956;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dad8d8bc8a2205d6f4d036e6f15f90223b5df58075c372af419203afd8704c14cf2523ea0a3f83443b6f7fff30050af6d34732086b9ed2b891e941725482422ad7e4531db91c537;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83e5a1c03c528915185e92ab949e7f3b1dd3e40221b34d713c3f553ff533c58825a5755493227276b01864f0aada3c8255e3b82dbc5029d363a508094f08e80ee60b45b640d4d079;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc12c05f749d95cc49d4086f00f06c7ab4dfa7555630c0e7e540e84553e4126c303b829a6a2bec2d3e7da208f6e7c7faed9789138f409ebf05574ce245c216d08d8c18a389dfc6b87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h620f97fea75cb7d642cd166c0d15c8d6011d281303ff6972e594266893198f0c30d1547c3c3f12ba5d257d05e780e205fdf6dc1fa350228617b61389265175f4141500124abd9dfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd640a44f66e6a2f3bc08b0aba1312ec0389cb4504384c1ff9c4bf4609cc2f8180376e72471cdf0ce1425a0b075b2bb0fbd7973025b1fe9215542d061e69eda4ae51360c56db17ed3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h405ff0bb41ae59b97d2d14ebfa8bf94a81b328775ba63016356f273c4b68133300e2e3a91d968e92e7efb6256aaa47ff518fd22e9f75b538883dae520c629dec75961360f0138213;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bef7e6d2e647243ad3c9483b36b9c26906e17e0edb0a76c4984ae2cbb1140ba3555da8e96529f8f56ff0fd2990772a5c7c90fe10a57cd40993faaa7c1528066f22da15073a4b229;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63568a5cd4ca1c7b4238958628c1d0922364fad85c6551e779dda03c2d64c2d6d92cec90a4309e61ddad827b0f09b39201591fcfebfb5bf4ee62ce137bf72ece55a619bb66e35750;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3108bc3b3f58573aa3498223b1bed573c86cf2095de3045ba0a3b19e3a29686558c784a298b21970f0b797d8d2796564fd1f6a0ad44a3190a6c930fed8908504c4e6b25a704ceeed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h855d58dd56f80e0c472358bdc8c0aaab73c61cef43e51127a487ddb0a730f6c2102f4d60275c2a150b1ef20bea968b39f143c90feeedd1a4475e653d8a931e0e07e955adaa2637a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6525ec69ac60bd13bce0bafd269ea417da0c758e80c386ff4c0af990ccc6f1e6a23273ff64308bc32449410f2849adb6cd370710ac041a7ce3fadfef928fe6e882f1b9a68782c7f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90ec41e81606b34e0accce949c3ba7652b62d219491fbfff713f4dcbe84844dcaaaec95913fbe891f75f829c30b667c66c24fc7f3789bcc5bc1772f55ccecd2cfba21ec02e8b0c49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e2aba541073cb23bf7b93277239e8fb9c5d7858b495a8522ec57a1e07196da807f06c8b0af618385d5327fe24038e0dcc9afdeef367853a276a6ba92da33bcc218d4e480066bba5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h257dfb39021dfda5b1c0db33e1d74a2dc1f390fb8102b2c538de32ff47f62988d2abdb4ef90b72701a279d28720b9b44e79ed2f63598f86a75dcdc2f66352e71b141ffa78403515c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa0e914e10fe9b62735749de5c2772c3f18f0255dd74d18e816102ddb5808adc0295ad8f799b6b819a7541280e86e4aa4ac11e9ed2175eeae40f8e4076cc501dc8cbf2146b0516a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a9c76cfc78e31695014b33e08649cd2087e8a9d3a48d186a8934cfeb1f61392193a5066a60477c9c10514c47983695a1cb07124ec177f5f6286f74f3c5b2f3803b4b8c5f2099e60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba4bf3ba41c820175528bf53b5646e073494e0a67d03d740d7502c13e9098feccca97915011b0c9bb2c0fc1c73e336b82b8ede182212b8d0abe38e349f07017494c9f11799595ad5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf357e6699a4be2c504ae395b34820e0f6bfadf79fef859a7bf3e9d8586b3d8f0ebbee30d1ab937e75e4d4eb0a681b7119c1f2f9a98f0f346fbcadd22c7d9c8cf2a69e52d9c49dea9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b03d1d6ee9b9fa969f0f21b2757e60828b925b4887f8c0c4ebf72f00d4d5f6a7d030789dc236937fdfbf8103713dffce8450bea4d0eae80f7faf9370ccd31426bc0bb027882ea10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h947dabdf058e99740bd632d55c59259985217d29a4f7409a69dc378da713418e701e4049f763e41beca3c66d24d6f88e3a331b52a2821b5bcaa5752238682e2bc2e9bae9287d8e29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc25626d401286a43735dc635d44065b649dbf911c47e35969a1cf7c20946e770a1baf287b51d6442e6e0544f4bedbf61189f9e960e417895bc9d4a4ec90198f3c02063fbcbfebe43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1980b0b47eecd1f944814ca359725e92fefdcdcb29796d8b786dadc8f0daeccee182e6e0a1d3f045ab7294ea1c1f3eb31985c747bf5da458510050faa416de5f743c0a8e0a5da64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3122c432706043b6e241f29f26b56c2f99798d500dcaf39ccfae4cbe168c77d685f9b9c6af9dcabc09f037f4682c0c5772797b992f0d2ca0912fb6613f0695732ac43a624d6dc5d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3239c7954e717da0b66de6e6ed2302b7f7132b938980a7b73d9b3ca76e5966a4d56afc3a50f23e4c17447a398426519b485f8e75c6e8de764b44ffb4eb4bf71f3606f4f88fd4da5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86f51be37ae65bee144c539bd16137b8d3a586f394e220802852a53526c1573d596e5ec7319f34d439379e5fc620c21cb1b9aa1f8a56b5ef2ebb83276b9a2d4bfb48c94446b4dcdb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e0d5edeccfeac4fc48a9da1b0cd07f593f3a4e3006137bc2a19adca840d36210683fc654b29596a58a89e206b8a46450e01a342936a69a3ca3e5573f298c1ff24f1532a8c6119fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4522a4527c7e1f1fb1dd75ee61698919e157577a2563f717934ffff7f1c10820082889c0c6a83c63b795ae5aff6f08ff88796bd51dc3e54acb6e05beb8fe1fb1fbb343777a53cb48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec7bef74b6d4944e019aec6c718e31ab6bf329a007cd68c73b9b728deed795973ea0aa13d2ff739901a7d86c6ea5ca8d18c0e142aec28c1f024efb1f16f1fb80022eb33df49d97bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6a7c38d86234ad723ef7f0cf4faf361c88a8124fe2e0831ea0edf0d554a78e1a79b666508057c84391f5c95612b5e4e9fd5a21f5ac38e622b1f8884def0123dd6d94f66bd8604e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h904a16ddd4f6805b2f82e9634772699731cd50e8e538ee0e509d88aec4daaf1cb2f6e69b13d78567729030e4060d77bb4d5d3b0592d34ad12a61106c47600475f049b679245be96e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51023f6ab11e3f1c3716928191d04bed4af90ea933e76b03d6f6f0dd054715eda27fd72a2c273c1bb4b9e4067913f072c89b3b64ad819485408b28b5946f8a2b4a7ed06e674201ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d140f202e3a089b2fb2d70b2fbe1eb63e21425405b6b36dbbe460f692e9bca3aab7cff8147956fb6025a4d86899dbeee7187ac0eb7db739047d274c7b4d89dfa0e922960bd86c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf11ae79526d0f2043b144061577c8deca93ed989c1ecdd774fd1d4703bf4b3effb336b6fd4ce179de01b24eb147feff3da085b24766197eb6d0f3cec6794e6e3435d701ee2394b29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h842e2a34be21099ac76bc137b465990b58de5c4da379780980c002904126e49c29c58560ce76d13dcee5a874d88702f83849726b4d323571bcbf99fce69d87a3346120a57aa461;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d80f0358c4420eb051f756c30d5dea0b656a127e778de9dc8471d7a47e6df75dc5998af63f43450cc620978c5517d99138ea95b968edd756a2cc2c436417ba47e342c403753727;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5982ddac80be277cd3e351bbde4eacfdfe85327b00db3d35bc2802d295a40dc5a0afba05da06f737d4159b50406343692e29ed400965826557ae789527ee964041b4b7f8e1843909;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habf97b7bdd9bbbd12a52339d64f767a18907715555cedcbd50d07e9cf3c9ff432bd851384221254aaa7688d416c5f5ba14003f4910b5b693ed42788dc383f4129eb0904335804d06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3416491e9cefa7f703271d5cc28df44e57e257af12be9e54d9ec2f6b4d6dc1e9e7832259b1b855f30750fea87df1b76f1aee831a9bf118409450323e3d8beab74a6028b86bf219e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74e5e20abc0a4b42948fe7d275c5cfd993921d3eb48f7421d3b3f32c60868b8b39f0e7c4165754aa7cc5bf3ab3b516b7b03ab7cd1d9d5569745e59ab620a5bc5c399a723da40db2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f5eac9fadd8f43a2fce324089f939485debf89c1d80fe24186d230e1dfedfc4eaa678c6e0cc7b4922a862377d715fdc6452d70beb0ac0f7dc4d7c44e7cc9358a25cc8e3125fa0d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cc2d69adabd1045cc2b3ba0e6f851abd23e4ed75c2a3ea4f6712823e0a7751a54721611087568e096107534e78e07c0ebeb4b167c411c8bc9f6615921675cb576e9dc0db8ffe61c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h675eaed1c23921b03d76b51039c0373523ef13c41da129cfbbd5f7053af99bad8954c95eb559dea9501ddce63d31585b46d0ca469e0069b42e1ec4db2cd5b04480bb11aeb40b960e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42527a87f8252c1a24dae818ca56a054906a54ef6ec237d23c1b3ffc68353f31c4dc31d1f229f63e82b6cf65a518ee1b8ebfe62df6ae85a368c2ec76a74cba11cad10c104f80f420;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1379c059ccf9503ba96a75b8875f6908f92ba01a3b9760ebb2ce0052135fab3d5340d10dd3708fa74af03896a51d47b0233af6517e9e842eb76946b5afd3e9e04bc588f055858695;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa4bb8b11cdcbe818a94a1726b2f31c6f1a5c72171435d9f524e7565c88d59b7f10709e94bc67cb469d4b2fadd1255e8604956775332b3491fa18b0845c801961d73f2fd9034e461;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2dfca211bc1f807835b1dc73cce3f4819a2cc6c29ef2f5c0d79dd7a240af7618e81b09b7b96de22b7229998e160ef26dca2ebe32903c8aeaa8b0506a96175973507f419babb5b8a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61bc8b776a5fd8fcd954d778f852b09782e66d367e22f8efef2de40b7190833741af965606e31f2365b13faad70afda348761c2942018924e2b01c3e1deac66100cb695b0e27ebe6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha56370a1e7877ce0b953d20daa8633cd74a70d5ce127d071dede03d2af541e71103722e63de1c4e4854da52d341620ff549a91069ef09bcb379f680123d2c8bd94cdcc9ea4162321;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d5961acb732c74e556a02a01164f341f60fcd9c17df4354010b8a16e84c728d749f505a4b32809fcec434d905162205f9baa03ed9671007c23fdedb6608c7e31df19816509115f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf7091e74722fbd9835f4e65afe250807e19bf49da9dbc0e5635b40b9f77a2416b02474df892b94a71cb34f9c1cbcc8c8d728e1b0837cde48a662ea9b04d34b4140025d2eaa042f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcffbb402b594a9cc4616f08778e7e9abb1c108a9e8f70a202df772f124c16e0c077e89e57bb467b4f0e97f27f8f4c3b984bcefb3e56794408005ce5faebbd394c0d7f4fc2a59a808;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h982a803ee66cdd5a5c9abab72692dd11a4f74c15db216094ede4cce6d5dc77d595fb12afdc86c5bc9c8cacf5e5896703ef3a2e80c5a6553ed7176fa4ef8d6e54384f9cb9a0e012af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5de8e83784a4a186bb1236f93e078f44d70e071000dbbbe0694d09f19e7cbe42b85f0e1428f774a30bd9ae4c9df6eca9d5bbeff28daa2b98552e6b15fc953e45cb9ba9de86ddf55d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0d036dd63a3ec70749bb9d74d50fbd46b6d703592810054a1e42c46cea3ad8f7804375914acbab67bd03bb1f4307801ca664414762e067e8f3da623ac2185ef793592758268a3dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31eb9b2537b00d4b851eda5435b4e1d7fe251a71b2340cbf81dd40467907367f6ed9b9555602201df1fd8982c18ae24040ac38470ea40313761aec807596ba5784e88d35a1ff6d95;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4c8236f0e91007c76cf2afa2c50fd8cad69cbe6c8d0fc8d68de0c8db0b06663c9ed21df37f3b86a3e196a1f55ed728e5013fafa191f30633e9bccbfe8af543f685153f3b1d3e344;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3beb95d28ced45a6520eac188d0049bf760caca4b38acb81b61da2f38b79578ea4e6cdc5670fdead495b21e28378454c5506b51553ac4216c76ff61d5f795b6ec6106108f806cb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a65ae3eea27ec993cb9b3f5b544c6b1377594b2275c2b5e10eb1a27131fa61e853440a2e57d9bd210024b736f22c8239b7c71b47c692febc7fd6f71838c59ea0f934b8eb302acb2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7b01cc8cd7ca9f85f4388b8312ad2589289ce50de9ff9c8eb36b450ca0b1881c52e10bf6b8c572f522090f2216a8ddadc5d681bc5318b0313a7d0bd6d2cdd4ea054f5d6209cb8c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7d438aed93fd2a84ccb41322a22e5d0cd704fb19444e466f6580be070766b92d2804d88a185c5c9aa149ec6cf885d5f060f53c3a3401d5b9b4eccf3ce784298f314aeaf29a8992f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a300b3c765d62e49fb2c34caed916d9540ddd9f0b70a903cc339d3bc7f7ad89e5463f50a038b2e11e556e980f5072d608df83963aa3f18b1cae54642d3784657c0de7b5f0b6df3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5925c7c750a7d36debecdbe73223d548b2c204b5b8c134d6605ddb4b213d7c6d8bc4b3bca465a42569620ba7c3512b8a6f9647a5b62a9645ab680a3f6f3f9b1102db24c214306208;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc83ddc1515ebbac87a1d17db447a0b36c8912cebb01b9f57ab0f12d9676f41f41dc30c3beb16eef0f529e0861b2b5da2bf771e680666ef93bfc39f1c85d45f1a01618b0869f20e7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb69d11b0da58513a4a2750e149fb7387c6252e6df1a4570d72dcc2e5f00f8a8aff2f287785327531d973f8865087d3b09573c054146f02dc451c2e3af4bbbd73e49d0231958401b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc01c17bc879187d76cc65809716dc4a6c9ca4ae83d6574c4ce0f820b2bf77570ad7394ab811c0679d77499ce15942eef1e3c62279c5d146f3c22ae0fc705a2f105b1e865f8c921c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2c19f7b8cabdde219bf474cadf81c4036be685ab0ae63ac95c5d8b09a607f3e4f228a401f1014d203cab0cdd8074c03f686dc0668d731b7b4695795b1768a078809ae479077c5b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a769e6f28ec4b85040f8448f8a4744796c69e5c6c89e9890d52206b3907e178c22e3d28ff46a3b1916dd46613b6eb11a2ebc3782a2e444e5f81f0470c447046d6cd037d1bd2f652;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40c7d3f643cf884fade99f2387f1e867c3baf2e047cf9c99b1350f4c30883936e0364359e12e66bd82465a3f4d589d8c48ad0d471a47e7b9c7de7c17107d4a7cf4905609e5d5b500;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfee34732e00cd6c70db83b73bca5711dd751aabf9615aaf461ae5404dc8a3d154a9f3eb4a06e1ab827935164b96c9181558a0a41b49c44ba9dbce9cf0c966a77bdccdf4d2192a3b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7374ab10d696b98877694845633785854b82ef68decb5b12acd730e55b3ea5ff33582b6a60ffb1bbb8893cac7f222fab312e0482ad896e11d809d1517c3090d81a5d5d8d1ebad50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93c7915a254dcf649dc68500b2c2c86636f910d9d3ecd333ed2e4d4820533a0b373bbe2851461a2bc9ffd2d27726151ca1e9489f98c1ae2c187e5789efccb210aa4255c167ea5181;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5472c319c0de985c2bd551c177eb1d79e2509dc197d5a55f603af3323f58fc6954efbdea9df6267f680d5ebdf4644d41c97a8c56cf83d4e47a23246715847cf00a62cded403b63da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h747264a7e607d0ce3a57f673cf60593bf880a4adeb28829692a92b1b3f5cf976ec4203df9dc00ab11a5307867a4ba07e9d71814a686e41a9c29d630e803807127ea2b9ababc086a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hceb81b10a2effbdadc1110f87bbc036fbeab0a4003590dce4466434b63b19ebf18ee36116590c9c297a9344dad00815b09e538c89bfd3e650c719dcb374f88a86f19f3ad55935dc3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4920e1d70b015178c9c3a918d5adec6eb8a7d5eca7fa0802a64ae69b4b21cb35c1998ba94afcd397dccb71484182643fce1683866e0dafd52abb124d0ce64eb0c1648c3b9e9775da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f68d7dd5ff6078881544bcbd260130b8a77e7ef4c18b5818521fa73a70810a42e81a4e46a992f836ae72f7232beb3d069d5d160aef07f70ab50885ae6ce3bf4e0213146f734f79c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc097e728d99ffcace0ce52ae9681a0daa5ecfee9abd87b4459458f09f8f11d78fede62faa14bf15f322a492b7a194d0019c3ed844d5b579bc3a6ee0f40630e5402062120713049;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69b7cb2f87ff989bb9f5181f146d127118a9e71a93de009bdc271489c6419479f80fafb3597748de1a98f26e4d94b9cc2bfb7dc9c9fb7e9fb133f07ee1671368713bd6eb66973b3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4783a9e63fc520011a054dad13d790c2e131cec8fe71e79ed3a5c161a13e86b12c9caa14f92ed44ce386ca7881f60441902b91e0e0e4ac84e6fd268f19079ff0bc1b376adf5cd97a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16261ae10bd05766e3d00540ab5d40b3ea09a52086921944baf4c73ba60a0eead14064c3c6dfe485e5db2f8e057fd4e6b263b7aa343874c4f749e8f2b5c2e348fe23064f7e24497a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h989d72f01eceadf6a737f97cb90b6e88d71d274b4ac8f3ec1113b885b4b0d9029df1f8778bb5eac80963f26aa883323a9e53522fd6b7134ab0a6758acf236e890cae4a5fe52b2e19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93154869d07f56ffcade7311f9bbe1be29df7641a4c56f4c2b70bb2e4d36d871fbc08d8e1bc5b29040e9f11c78770328232424d123c79278957523627266ed01e96c2cb098b27a29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5f629a59c4eb9856f6dd946977a1b0d27f310cc779a6d86c1aeccf2ba49af8559382b1beed113bd4419d699030581c4619ae482854e9a55a125916620944a59e23bf13fafc2d8c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80fef333af0d42caa2ff86c81d35466bdd5efbf843a51b8fc345f31d59c945112a19abbcf98a66915a0c4cc4615e9688eeb38e51a4b2d75ec8671cf4542a0f5ce477875379a075b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he91c9e150264fac0cfeb857d108b3895d016b7cd37b2ea867655988e5b9d90118025d57aaf31371364cef391b1a0b1d58efbc42fa7fdebd43f94e91febefc83d9802e2ed47fce7cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habda45894d92547a65f81ffcf7b8bd9d569c4d6add9276105fe239742bd09914a310fd62265d5a5ccf1caa9fcb7d5b4ceef7d17a7f9dabfc10cad07de2fe892a4fb56783c8eaef1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf23dbe56bde3c6871cfe8374dd26bf0be4bcdf218ba3f2af41b3d3c88201f446f7da4f1e458a671383463cd6d46ae69d5efbb01391ee759d5c787c367f79407caabbcd47edf1954;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb86c90ead36318d9ea54f0f57d43968bcb894133e9c8a9aba776008b39ee538abceca92b2d8b93496d804c6d854e6c4e3dea3f757d2ab5c2f9f13e0c44f3b3e726c637c57dc74335;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e967aa2610dda94bebf4b6fbe15f1c17b54b23a113b41300ed60e13164dd71aa9d32ffd01495376a3c2c57fe305e4a33c78053ce5089d00434ab4b600492118ede6209d8756bbc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc09a8e95bdee07a38fcde86e4ea629dca0ffce7effddea1db9d635f83d5e5d9ee02530d03b959b97f2d1c690517e3cca08b9ceeedc6e6620bbd85def509eaaa8b2c8a167d8867ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dc2213d702e89b6c01418ba938d0c7ee512dd7af92b9ba2a11f3e01d66266d862a416034467b684d367b3cadfe0836d5dab10b137cc67cdd0a38b87e17a0c52db4c345d2836c41b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70aa2eea692cef651f8f698eb0c503f0a503ded934e49a0862f3a9808c21f301f044f722ff0f081f2f2715cf3703ec4fe6e403fc461542a070b60fd0de5cb29a6ca8ec5fa858f58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff5230f6b021b104da774513b17fd65a085f3a7601e79d4c98bdfcc202161b811c42b50207217ac1bcf0601403c3154220d2ceb94e3361d6d6a65f8baebf510a0b002f3579ae8060;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5bcc6dd13c09dc323379f9246954e85caf73010b1f1db2e03b0db73a6ca09127cf281d20dd32765c31f46d646cbfcee0f85916564d2ceac72a08d589a5ba0b777f86417d6d4a847;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68eeef485210c310ad63a3c31629459cb7b8e31ae4c0b5e92e0f7af1431ccb26c239113fe79d5efb1f9a48463b20841f75e75639cf78ce6a3e54ec8e9ee7f9e5f01ad90ff1e737fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h966301075ddf18c16b588f6d46ecbe76201be490e69b6eaddf67bf9ad48c3fcf70ce41642d6c1737977ead451efe309d81c8bf153b13b1811b0335c71de317f0942cfabf018c9044;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0c0f4e3ef60f6a81c7f6dad1fa95d4a2dadfec1b3cf9afa43c034d0d57cb5a4d0f29aa7056bd797981cf9031f49b7e5076ad2b4a6b4b479b2f325d473304b60ede6346cb0a3465b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3ca46da5366c7b7201815ad8e79abcb1d34c37eabcfd5c1e760909f4c62c261b93fd61552b8964d3652f0b254cb93162573cca6824a607c4ed35c805d34e0cf02c77dceb5f57815;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ad89e27730e690613856fa3006efbea431d117ae6825d5875296bf5c39bdd02b0554a066e155f64ecdf83156efe635f68122d2aa9a684ce80fedf1b38eb7a30001e59c740ca4d06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68fc66aeec40ff11ddf4b7e0ebb9e199f585ce50deee643b712302f8e511081b6cb70910f09a20c74d1b50d414a4808c86e71294f9b00a7f231c687012014390d1bb2b4306dc5bdb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59690172e4b105932f378431536a43b1c58fc538f0ad3be3686aca793e5d5776c319f01eba9039b7df8bfa459040f8667dd3612dcd1252cc2107b4a7110c8ef8324e52f811977455;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h949a940a52249c0d87dd1a143c9c69bbe1843a330286127a65727851866dcbf9f5cf51cd74d96b7d909ef95cc618a282dbce72b514cf6e06f472ac74e33b8e9f81e17553abe370cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h551583d4b1adff875ed548d9f9398054c6e46816d148a87d26dc1f0c7d7cabe268b47276ab48001b58a9dd7547acedade7eedb73ee40c58ba4b0c3be41c923057e013167d3f4fe2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0129e8deef342171dfc90a259f50b27b925da7ccd15e51416b9dfbb8eae3f04f4abfda46785d943275b17c1919a1f896491559d987772dbf8ab30da98f7afaed5937f603c6da476;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68184c9605e5ce5ce770ba5415bb2a8f85837d52c9c13dd85619dd55fa51d10433aaf71197d4092b9ababad07d0a6b925b9365384eada5d03abc07693334999d6ddc4715c517e3b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb91e0defef5afe18ab06b9946e3d855798569edc4da171dc19921faca546cfc3406b1056552abbbccf613612cc9ef9bd5b33fc6df825edf256f8249699414ff37fc7523ce4111580;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h305f9dcb32b63b4298c2ad4d505de33a9626e1d70e6e588f0650b70929e4be09bd765cc7ae05993f09e506ff82cf93cb916d18624748b6e0fd6b62caeb1477276a4fae079adca7dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h933d20b01a004e1404197faddd22bee3a86be72187f7722ea6c2bb7d370a8e65c69280b5dc7e9ab5b64214a4d26073a130c69e15f21f4fed4b1ce8451a27feaae768085417a82865;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4e83331226d844a8e3bd14f9d26f332d8c5f877368ad9a66c649bbec2bf91b8fb40e51eebfb612cf1ccbe7caa2b97c3205b64f1e2b245d346416ec3a875a769545996460a05f2bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h201a6197708da4c93eeb58ea67dfca16e47ecd7cc7436a3aabfa7a1d90bd54a37ecff7d58fec9a3a38a6e22dae23f8a0d3bd1bdc8b58246c23cf8ba828edb72f5647c8114ecc26a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46fee7a19c4966502f9d7e8a80a1f9619596772e7d81b19a1ecf09a5b83afd10a28c4535fc7889031e57e6487e4c984fbdc89c5d9903b73d641522575fbeff46a798173ae356df7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b567085b299298abb9aaa2f0d4232f9a0c34ad907086e807950bda9556e520aaf4f76c49790dac4521eaee85056dd81bfe37ddb15c384e2ebc5ed0f6c317c15f8610da44d127346;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb2ec244ae87608d9ae20a4d571564ccdf14d7ad344f59354eca1dbaaffa7dc823bf82f221bbd5b62ed91f26bb558e89873b343f6c066589871544f063df756f2cb6c2bb704a6f56;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1181ddb75cc74cca45cd7fae76bf4796363ae2d1c332bc63295b920e7c1eae803959d3e0cdecf8562770a29e14b9bf26f509726138342c1ac01019308be6f6a0f1fcf4feb54f0096;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5d5bdea0617e306dc7024900e7fa243a70a1aa3f561ff9db9e3edc6804f43fce2e98e55009e689e0616f2907eb2f45a2ea87c6ba3406f3ef5a4f372b8c43c7b616097776104aa53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed3c2b1feba8c78f8970fd7db8073f287232370a58c962d93e9f491a526e8f2f3b81ca256f09823a09bcd3b950caf9333ef23ab9a07e14e671168a9bbbd60d615294f532953734a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h867584dd9c4bbcdbc1682de6626d5468662288de6a801b3d76c858e82422edb17ade62274e2685bd69a10542a2638f09484cd1b2bfa27c91872751e8d09924a57506c8d833bd0c12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5772113e120472b4ffa2726362cbd372fc0c7437cd66a71335a428cd03a348151cddbcbf926adef6eb39e8a2b26b8e616381b14705c669ed3d4870a4510583bd6d5da0e622a369df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6aaec2a2e6766e70e1e880147c91bfac4f98cebf5c9395061af6aab7c5fb1a19df29bbdb080d57f724832bd2deca2c2a700221f4d391f5ea4cb8cfce4bd06f6d25d21a06dc7d011;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58bd7447cb10c31c0d37638054fbaff2ad051b04cf880929f451ff656ca2f5acaf2cb7b53731c97259809afb8389d534d914f3af5370c31198bed6cbb80b76d7b1f1f3579281d0f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc200d7060ab2bb5f7f69b1d14b65a36d675f764833b5e15e90e165e44f7864a490b35038de76145f5afad9469960c2a5d1140d7522767b2db75f06b2d6d8c50dbae65f612082261e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a374ccca4c96c3f348ad2c2152870d92dc8b40846d4f06da75bd15034023d6548e5bb7542e2aa4e467f2c033700ee2b097d58471d6a0180300e94b52db7dc76d741ac9f2a5a841e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76d967368cb32177102b2839eae63e24eaa60469c2132b9830716fb96e0e57ec797e1f7937dbd48f274dab689c4884bd776b874512220c52a7cbfddf2336bd4406ef713e133b9940;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h304140f5ed78a9e79a777c5e0ca8d8bdd4cd91a1da6f6c5be8c569882356c8521d6c9f9ff09ff2df691455862a9242666994a3f6c0291172155e32d92714ad67cba8a3b8dd33469c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ffb733f27e60c50b42fe6d5fc4e86475a7aadfc5deaef89066f392e9182fdf1255d649d468a86ba1119b2c5260b597bdae93d1d21937f99fb21d0e6ac52e86f4dd323721088e30e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdafda59674bc968b191ee129553221ca0bfbd4507898df5ef859a6f3da88758f4358fc3d22e90e1afd3223de1a4e930b10fda7fba4563560f1a2ee84245ff1be77cd8a77d82108a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ae3bd7e59cf4e136826901a15aa7543e858de9543c8b5d789459bcffdee2319740b1cf68d28e005b66507e51b5b3bb5572175ba898c000d2a9d9cb9f5e620d697c153dd87a38a44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ee869da7e90e48cfa6fc70e53d56b7086f9c35a50801f5edba5a7da912f9369e621125969ee9e5d911396d8d6a6f6195728a2a8c6da29e47483041f15c7f9beeb7f60314d5dd0b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52b8fd0221bef24631c55bf1ee0d18808ee6e923bb0e0ecaeaefe27f1b49abfb5b03f8a556f2e8e36bc4bdd3b6e9ed2b63627e9dadf180e7f3a5704768287240e1aeb0c2c93b9c3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98354e657827d4a9b4e7ba7d81ff8bae11120c1cb0adc589ee5d9b3c75056a46f2282301908368b7a08b4f720197f979db2f5a700a0fb9e55e6e906e34893baaedef1c7e19bbf04c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26ce98133777f7335dcb0c44fead54d5a6512cb6b74158e7fea187d6e083c642a0c30f8560f81b80f0b3aa42717b387faaa6023f32a973d75443e4e6fb5680fe8b39a8500bcd2b6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fbf98ee35458a8adafa6ced9bf6cd2972fd23e71ccd4327c690f7e8a41037ccb8ee845dedafa9e6474c813d3e355134d9db1c9972cf67707a68a2f720ac95fc1643905031402f08;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fc267d8a39aac4934629e0e42f82dbf51bcc6374c5a433a462be6f6eeb241e9c09e4c4d55ff6d8e90313c9c192800217a0feb16530ec6d600ea15b138d3f8f37d887aad30087eed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haca3ae716d1121642693200dafa99791a97637c44ef5c902af59cf5803a229157fb1fa0eb36510c54def7b0549733ada4d11cba4cd2405e6c56af9fef4be1b188000ba938b69beee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b3b876d2e939ea587a522a1d67188889143e482468b777b95fb1e587d2836076b9c6c085c4cec2c5023c802c1d84c5f287f9df43bb548e1e990c0136d2f70e69f150a1e95bae7df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1411cd86aa04942befef96236f549ea7631e9ead86d7ea2b404087c49b169a5dc743451e9bd13fe1e31f1b18d4ded26d0389e87f7424410e1a3a8b7e86b5b52dd76908fb3081ddc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6c5712c6c0d649df5bddc748b3659c49854c6aa2bf8ab80168bee670492a83e8ac1c3c01739b00a0b6f9702946c681ebb3e23c40ae35f29af965ad338bcea7319e22f11b3086bf6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cfe8fcff1e218fc1e3602fb550c877280c774d1c4c941172336d105c34fbf49a145eadb6565b631abbc6803c0cec386075a950766221d0c0bd3213da2304c3fdf42a10825d18c53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dfb455416f374d6d8defcf085e81bf8c9739e282a51dac66c184cbdf40e30a7aedb27db6fd8531397a5f3b90cc4272be5b7a246a06d61ec1bcdb73bb771665d03453b2ba5aef62d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4446fc9c8a8d30bf31fed9e5ae5e041c11e17bd3a4d961aa3e65b640c31a678ccecba9f70e132f93004de1c8d63ec85aa0f65cde00364dc2932b5cbbe1faf6851ca13a94890c21f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84f9b378574b9c7b782ac89a733f5c1665e60b22a6baabea7d255599a7d9c4d219752a918092a57f3cfda2391e27923656202e2289f8f51219e8eb549bdb5a6ef8a1d40c377471f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf409c6c2042a071b828a4ca85e1f8bee89d845afee49dbbebdfebb059c16c1c869ef0eda02b1c60bfd2c20e43fd8213106abbf265d44f53e2736034f9fc77b62505ce9e654c90d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9be62ca78aee40fba0a1d4df34083d191faa7eeccf29ebb78b2a9f683ace28e8e841e583e9e58478d991b7c028036167d33fcc11906578e49aae3738d732ce8e99c3a4c68cd576dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80d3a7b93231cbfb4f5e7dce5d491e2a0213cc7fb09e608eedf952a6bfc986cba37bed089043a50b1be93f0fb0da6977726d2c60be3e2a7e4be67209ef8552b8ba8d66137fe63caa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e7ab88123ac04519026690231b1f9c81e28d5fb32f2b8ddbd1c8dbc718e591bd05bddb804782979633c85337af288b6c2b87546d7de82ca22d85eee3213ae886e8c1776e7697819;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habf48e345ca9af44a97603c75b7de2d6273f45afd3a131e638f1b2e0a67e9688b120fb2ba33905e9a014da6abe9379ec681d86e74c1d1f433d56964bb09519f6ca9ca7781d5df937;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h267c8c556f0d9651f517676b292f07ce79caefe15d756ec2a57f23ff968a684699b34da2eceb0780eada28c352b9fada3eca67e3f84a034bf26136d19cd6c6e7da882a54bf089ef9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2be0592344f29c89ac8d1fdf874380055f491ba382dd5081fe9613d537c7c9be4684c6d86248428382e9abc4ba3dd285c315282b18b7152d69cf3a7bcaacc8442735958b54613033;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5019e77293479778df75bbb6cbb364b70e11d63a18916f7b05a3c7bd33b06ae8f8b954aa4999ba554359679f913457d466fcf285cbcddc9170e83a56f479ced82b2816e3e9314480;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11be889aef0826b6b730fb3800a5c616143f35c72f67306cbf575d7e8ca854865b11f266bb13aca1ef04280c74019523cad3ef1bea759afec977fa368952492e47d90062a2cdb2af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc215af1b7bd7f715931ef7354df53568ed68f90177b4473936d03265e90a90562c079fa21ae2253146f88fb3d455a81c48deed111656ba8ba8e9d0b76bff71dac3e988a538f40a3b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7548ea1b329ddac126b19d1a00f11eaed5c205f9ec963713a27eacde4568996affe6eda833175d0f6c5f11f5e9829dcb1f86ec6db334ace16d22bf8b8afeda41f5b964540b90f107;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f308b8d2da5e16bdbf1dabd2ad7dfa5388125ae7673ce6c2d4848fa68d40459ea2431a3b369b63cefc913c4cb42a55e1cefdf50c1cf464c1c81daf7a96b5b1ee00102ad21bfde51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha892c3231c2efb0e0c1f031552190ca87b5ab684e9d2e0eecfd9d250ae3c228bc2d0c3aa81ac86c0c745506e032e75c680336bd3862ea98d35333d46b23c36f65fae4a0a4e959f31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb913894af89338fc5e5d172de4264da6630f0b60bb7679f1fe8d35860522532da016a9bee8eb79fc3a598f2a6ea6f02ba113a2e5ee6338c3dc99709ac8db79690b0b53944c3e508;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e0f60e40a56fc8b25a483833103b6104daf193630d3c893636cf2f914f65cb75e821d805b01f7ecc1c9f179c4a4903fb40c564817b887ada50e75968e7e17d960a7c5ff11b4155a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72388c160ffaa4f8bed3437ec8361f488207d0ace8b4c4a72ee21a5de8596c427e6d229da1c9e85095f6e330d85916ffeaf3507a929942cff42b8e655eef2df56fe45cc4fbebbca5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85fab778e433a262a531247efe3b4be66a0d785b6e504a929e17a00e18eb821a03382e8bb8cfa54b5c23440d7a3fcf1f79c85d66005e3127415d08a15d18038fab78f92d30934a78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb7b50e5af1921c65d0b7c1ccfabae80757c4f5daca7c77062f3f33a03ed731506b768e076c3d3d9309a9f7c6a7d36a7e2e4fa79fad38f38c481a9664ea79f7b07b8c96f5d7038a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2be3e02727646cd007d1e3ca3d8720077da31a8aa2f296f7fb751fadc891afb00298d665d626a77adfff42d93a041a961d75cf3cc09f2769ebe105e5ed4c6b05a5b0302e729df432;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5d24ad5d3bbc91baae9dba368269920aad2d9aceaa5f8c07fe308c4e8cd303bfe57846e332084fda71ba53638641e22537812da0826e73a9926c8b288d1eccbe8cd46655b820b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac593305c95b5cd43d9979a7869f08572869cf4ca1a937c23ccb6e9c8732b3ce2e94920c2bbbef032ef69a908a86bbc4cf67dc6c7c774bbae363dbc7bf9843a7d56214db8b8569e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5208d19361b53464ab0ad7f9739479ec44e1505e4751aae3e651fffa23708e889ef2e3b0960a4d6a8cbc0fed5f4b71e5bc48d46a8078fd10ed5402258bc7ef2d3f7c0eed18f62f69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h501c780335530d6929e6fabee1fe491d7a7be672745928f169ede7670734aa807659a14be0ef312b013c1733024ed9112b64ccd88772f8435ce7897bbb49a22e05fa9790714d7c4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ed1853df8362bc537a6a58ab4387ad6887d310b9e1a7adab61277f1bec31a4254da6e9e1310fe65a58bc31fb3ed6a05d9d255ec9dcd6a0890185dfa26582c38992c972cb2b16c75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55f5b16da1e8e8a54bf02f34bc2786a0ea3408bbae8eea17a658caffd258db9d085d2186d210bcbc9d4b70f6e86dce9513c5c679d66972061877218a4c12a8bbbc7915fa038d2809;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h780668afd09b4b246a755021cae20d39221c771f4ca8ccb840198de68a24b05224596686d951834af8d06e7276f50e890bddd6450d64d668fc8d4551dfb73f84cffa450f4ccb11ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0c74dd4a19f88925a9d13865bcd0072a0870bf3d278de478c6c85cd3f18f313b3d3ddf34249b36cc0304a6736a099928c9ec2ebb8c9322e57633a4a3dbc22f42dbfa3e96cd648fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb095754d2b09121ec63c6488337c0b13fbd019cf52fa5e97fb3048c667e5d1c212ac0ab582b2d42141f951b6bcf8fc93dff3fd69378dc453fae1e002130ee007402d1c63209fbb17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h536091d62780deff1d47741a0ebba2838ee0bb13c904fb77384e019fdc666099f807b1759baa86ea891005fe48380dfb73411d4082aa065913fe850b22745433d1cbfdf67bb1120a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd980fdbc6bac0fb2ea7fb0fa2416e6803958376e8b8c7487be4049ea60e8f9999f52f274c379c4a1833943de6303aefd079f6099ab2ec9cc07aa0bebf1e70cd7115c6ab29be3d977;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ae528ae26105de771ad6898d1f4a8c1c30e41d64c0d3cd2e86dd0ef77b9c3720b556cc665acb497ef74cfc9cb47a2e0c425e7db0481dfaffac5f6ad92b5c4c377c544f85d02d877;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0093fc8081c85ddb596164487f078a234666e4d094620494a26101e88db54ae64689013c149e72b400c54da5fbc96a1fefed1e48c3913a29161cbad26f084f6f1a71ecd932f09e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6b4c0f90c6d2fbca86346bcafd52a905de9371d869962ed1f015d9ac35e82cc035ebcacbbf141653fff65b046ae0126b9b69d264c3bccd3d8668e405a0a4b78d88813b5ba90d4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c12cef002b592c4755c5c13e3f8bf7bfb1fc73b404266a45a0414d90ff99bb11058031b73c2072d746ada9dd8e9d14861b0bf00e7efc0b659baddd5106a67c95f12332699ad4c4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2949154dc853ee34214e2042ccd8c803b7454f65c451e82839828e14fb8a8b084d702c96b450c112ade8863ad6f82d335a7a8be1c38d5ab54680428bfd9fe7d36e7bfdfd9b76ebd7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5565ae1e3aa67d146ac63a6efd473a5309627e449aa96e63e87a42c38e391834b9cfd0ce32ef1ae2707e27c534c64b9af09a13e1fed714d39195c2cb7a9502b2059aca51f782ea42;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h486dacff1b7289d925db693d39722ffdc3a10cec8490ae5862e75c80451df0b0525ed94e3d12bff685bffaeeb633cdff975425a74c387e047f0ada2462ca8c68cbfd23ed31134da6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he907b37eb07182d1f00be969fe450c1b00b748ef0b28896c7f71d6419a144dcc2922c992b52157ba985f36ffd389bf159abb848f2b6ff4dc12db76775388101ad2665b3973a12597;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca124a955b1bac6906a2434e18fb2b83fae25887b8b9d7a0d82a27f16e97454276357aebaaf0695414f1cf24bd634ba66cdb6698089dce5289250ccfb5078b41acfe6799aa154a50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h789ae1b49c52b8246589722b5f55a16b8edfcf233c299d2f82a69e3884b890209a652217ddeea23462949d8df74d87134ac62709f9e834668068c1512b28f21444c6f973c51047;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd01b01728940218103097d29cc2f2916f6460b64ee51424c28a1e6efde36c1481eb8f56fb53d5a88715b040131d95d180c5f6b01f62b6c4edefaaed74fd00f481b76e962f1ab434e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62f4bcc89bc20312c20d8756ec0c47df6d6fb2a683ced7507bbe8447cfeda5ed59d8dd17d720d5783e9d03dbb07d317a58cea8eeddd5a4d91db5b9324edbb2c6d4ec75ae39cdd2d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7eb5f863982a39412113d9ab5a09acb619c65693fae5dce24f5951de6935e88bf1929a99bfc7280dad3b65d411d6d0b766ed032982815c4127fac814830bfdcdb5de8c08a2462967;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h616105c13aa5da5137318d3d96001a4aadc49efd56b186a8e06465cb4438b16a26742d1221e2281156a9fdf5d92b0a74c6d12aad1d8bdab34cc0ebdb0279913bb9f9d3864093f419;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27ecee1a884c354f9bbfc42c9cd51a66e176fd6080c50ee8a520182e05854fc9de0351bb413fa4394c0ac93db308dedb4aaf31cc9c776a7e2ab7d6c60767d76ac3a1d6227db9cfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcabcd9f893c75ae119fd54bd59b6a5f4c73c3d8fb159f3079079439a2ba569f46a2b3b30e155872e88385a631cf2d0b08fed90c362131e2c17491943dad7edec496954501536c133;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ae32140e589f3161637c5e1186919bd459d2608f3a8e95884880a3dbb1e22b7e2f729b192ec80738b3893304b003f6dcc3c6076970c695ca164f5bddb581754212d4ed56269c202;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h592578225fee5a261fb81f3626e71d7300f52f15434f8bffaa45d56e58a591704dd63c457c523a1bb9fdca01459b8d82098926dbd9d66b6d025c18dc1c0940b3765882daf841d54f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ab4396f66c1162562e1c01fc7dca6f0ee0094b57138894b94a7eb12ca60425fa9c98fe846fe1e851d69946c7e8c4f58ef87000e88e95ca4ba3b6a45a59ace8fecace310b9f2852;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he28d08de3afc19f18f1136e25e117c9b46d140c4287e1da00150c94c0f2e72562ff6ad20fb340b46354bbaab362fba98f0986f414da087cefef059b6e8c1a1c414dacd4346e3b1a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45fca664b1ab29e544cdde433b8d12aaafd68a935dea47146724efcfa330dc117858f302636c1ce25315d6ae31d0ad79e00de1e461e49ee1ffb48c7196341a3b3787623cc0f15eff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffa22b69c6da7eb6504a8b6f49bb5ee63ffc3410d5b72224f6007079b9bd0dff02a84380c8752917a0b95d1d03bb29229365dafce4d189fe72aebaade339f46963857a5b1ea92ce7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa83bbbfad4ba9381d2f55bfcd1dd28e87c0e2bb5bbbf04ed28e987ac2bc0bbd0533dc854e16a538a4c4c23e5783e21f4502d7826d6da83e6a60f0481a6d86762235c48f3bb1067e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1ca4e4dba76ca5f4826bb19f5f8d6c6c133bb7eebe781f708d626009788c0557ba4ee0a3b39504163e9311ac8332d1dccff73d3ec8a2f243d34d3253b848c99a9c1575c4ea67db8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79b7deea7878bafbd038044665e1f9de3d5d60f35df073f1bc9166b8f5d8cb8824be9c9142dc4beaec278cf51afa3515d615f0ce2e75ee6519e7f3de1fdd16ace7bd1797642775d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ab36d3af9c1fc20c208f3e17dbd196676c5738dd1808485ca59ec5a0b0d14ff79c4faf7d73f6c90ac6b3f98d83dbfa549eebe1cc2f28539c979bbcd973e386d858d3f922b40ac5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cba2961377cbdf6b779db3792d020d026afbeb4ed811d032c5d1359266453b505ae2363edd6c0e99d0c2f5be9e2ae679af60088a0102dadd2bb2e60543941dad08ba6ca4401f28d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7dfe08dcdd970a1f79345024f1e3889289ff908bd2bae44f70ae289694b4d965d9eeb69071cbec507fbba892ea6b1864fdebec3eb8353fc4a08f994f7a9fac5499dd4405293b375;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca1a7a12a2eb4f91cc2f264de194977d2f010871cb58de0437c8c5908210d68001934c548fb5d72c4deed92318cdba359b0ad6083a941e4404bc942146419cfb2fedb0ee93d71397;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb62c54cdee230196da3ae409c947eeaf9b2a356ff495c6af178f5f14ca57b4255e3b45b1272b64e62f4260692fc3fc777980017f6e0f26b8fc839bdc664873e79ed3ad512aa71b49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d04e3578ed249fbb6dabc6fbdde64b18ea51a19b5cd3fb5b3907fa36e49b3a4ef4494962fa8c31cc659f1f5da37f6a6c28f6676af125b541fd7e5f46875dd4356a6455f9efebafd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87c8f64dcdc45734e3bf1b465662612497984b86cf272db93d0ebedceb30200a4951ceda194a1da0b61cf676f0eb1bea7b924de50bae5e6e078c8a7be943bbfa690c389f47687a44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ffa09f58df1ca30a55ee0570951a4a022e450763bd04e7692f999c65f0c10b1dc1da6c7880e88b16148f5281934d6110928c38cba8a293aa709c3b82adec213e6853394bb5fda3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f32c84c045c8656548c1dadc091600347c952dbed79fcab0204e813cbd68e0654a56e8500dab80d7435a0b13147f86d82eeaa56d1bf90254601d6922a10307fc72b2778035ab033;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6bce9cd2c753da15c4a4521b3ca1b0d9e2dc3088a665d64e68aeaa6c0ee205515c481507a924216c83b1bdf986bbf70fc1ed64bdb1413ef0da791ab6c0a601050caad454e7da52f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h430d1693b6689f6f9aa827c32d9366b0f063f7c9b0f0df710c63dd4a0d228727205b97c5c13cb86ab59a3b6f6291b958d2474fbee77565f556dd7322cab501bd959ebefd2dd03f61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95336b983edb0fbbfce8aa71219d613b9f24f669a9e6f1a257d5b4f2f901b31f57d05df699017b6fa926c2a1d67971790b953f4e5772331da8991eb3e85e289256ee5ae47fdd4230;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h284faecddd8044f380c7db92a7b0c083f3f50f3dfb770b91486841efb706de22c0c18963f0869d7f69f645eef7d671d60caba8ecbb092e09aa8c9b3d13cb40ccb8ab6fdcd321c4cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cf99c2d6efdd6169c130268a26eb580b9256eb9406bb85dcd88fe87cd907ccba50ebacb43553e1b079c85ae4aecd9088fd8d43acd861211af3c1a38797d137f905fad20d65f2c54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73fd5c0ecf33837fb561f4e492dcf9b3bef745901ab94493746dc04370abdbb72f91f6a5c088278571f090bfd08f3ef8bce341d34198dc6c9d85ddfedbc6b60f1ccd0b533598c305;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcc3f9f8a1e5433d679b72c161dc32786e81a0803278f77f4a4fb3707989ee44e64af5b2eb5524615bca37bd5f7a77b5078b907754d7aa079d543f6961a438bf9bad30c139c7d1cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b4885d5725ae8e5e5781043927d50aa9d87923e51110fe2b5ed55557b27e753ac978efbfb8455614b499f1bdcb6f963a55cafb220eece64d3dfc8952ec68f1a660cdd076ee2f580;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8082390e650599a25699d6b373fe1afc2693e3c97bb60d4cdc8cce570a312774017b49a37800e661f33e96bea875f39096753a7d9cf35595e9c4907bb7c830391d50f9d00dcc8c4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f981d1808477eea20feafbe851ab8593050176bc6deb6e6153e6c0f658e44c3bd7997c9f83d5fbf62cb1a02d0659a732c9685c0fbdf046ea84d1c3ee3e7fa8579317273ecb4aa3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb4df3a5b71fb1045947835bb53e0a0df315588002b5008414e9f6de4c05c8ba463778d1039ab89e303a1d82547b6107bf47f44722f5ce40da6564dd3a5219f541da7c935fdfa947;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a608cea216953efc5c7db237708a2d6f9e4f6a5a48fa73d800444867aefb53d1521868ec3d6ff9136fbdf6c2006240897862947a68d1b107e97ba59d02429ffcfc6b8d1b984ecc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94cf93fb737c557c49c88e00ba90863e4562a7a2e6fbba27ec6c55feee7cc5b986d28e9eb1ef5e0c0d8ddb8a79a7e9b36e92acc7c618ceb60a416e697d75116bcff6f388cc2f7719;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e989485b5cdc2aea8a2a6d065b3c98cd698fe7716ae7facebc3fc2c0c779244e4cca7d2b2d474ef4ab709afd2db1906b954caa1dd94fe8c63db36b11e87555934393e9df4ba239f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha39d1021076a5b8a748a7ec2c7ca6087597c3a04d2048c1437fedca8df66c797209ba3be42a853d8dc26dc92a9456eb8ad00f3554c91128e8cff63db19c74b54da655051bcdb6714;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd81eff20647a7d116c8a70526adcac116fb175ce936a79ca858df6dea6dbc938e2fbab83488634eeb20e8391daec8a24a0f3173fdcd47cd670dd4817757d473c6e2f54b2ba00cfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22773dd7bd88ab0ec874b5db6612d21676ddeff8d9af6951f2cbbf208fa49315ddfd01d1827078d04c75bd293cf675ec4dc07b0bb55314bccabaafb21b1671de676afaf5c0c1ba36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc25c870f301a29676670480d9700ec452630fcb755bb3a017d6cc8f599803affe6324b91478deb2c21d5498e0146f8a68a82580620f45fdd7d6707fbca7a134695f83e6c1db2a52c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he603e4b6ab9a83a2e56a23135cf587fe9133b825ae1b3b057c2a068f89f80e0667a7c08721a793450b6395f1f51bb039973e002041f2ebb3e265ae838a10d707831d4d96d0958610;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aaf469576b54e34cd096a95b02417f85e717aa60ebb23c2bd7e9a695d9f78d270554893f340e4ab593f4dd22447ab1534834bb6a04846fcd374a91c38208204c9e46b0e2e9c1942;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63067378332ab830416342c32a7fbee0e2767174739e5e26ead7f88edecef965a9e8339ac93b76862ba3227572e00074ca34374833c415239ce11040679a17fbed469964b2342fd7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73302a2b636f6b1c49d593e5eb51105b5e9c649aaebc92ab8e5ba0756348bd09d3c6d1f9a5ace0c50b11a4f56c8e8ee27bb017c75a9fe2ad25241ab319a37b1d93c0236210aa75d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h269e613b97159fcd2f80471022c1ec07dc2d5ddfb96fab6bb24856b640d3c29a14a9bc8e079b31088533cab239a1bc30a79af1021fa62cbdee5a00551c2d082bd1cdd0152288cbdc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47c5e75464c8845a1176a61ed2506eff4cabc85030b870dd0e06f2ab5216c2c3909a8c794e98dd0e28dca2982258feb5bd45c704d8662d44404b3634fff49fa3d328ee9a0d37fb85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h964ed033b276e46a04f2d026499df01ed26846d808ae6001782ac2bd5bbee97b9d26c7e17150b7a9f316128a3f97d8534948e64189df206f49a242f0d36d44c01ad90806be470c94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b613bb4ebb8fd4b9555ed646c91f32a3fab1ab2f8cba7fcf19148ad752e1f3487a5117318d85978e5928d96832d2b70058f35a61a1daca6363ce7508316eebedc064e34bc92ffe8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9f18a39564913c3f5065e01beaaeaa7234e54989885085566e124d2590648f294c27b72d6be81e3bfbc78cf710dcc5641854648502c64be51d239ea2d5d2e7e70c7e43cda513cb9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9fb5afbeb6c1f980a6b5a76e862beaaf3f817449177162fe0da69f2f777c99829729b2140dcad81fe5fecf1cfc33da3e0b03f92ba977c4692ed0d03b2c84dda122fa00e57daffc6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf05bcbb91113c7a747758544555186184c5c0fdcea4c6168c584c9ad3690503e1aaeef157829e12c05a8b25333ac735dfe6ce7c988c0262ef9c9fba7470b39cc554f68f8ceee28a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ac79ccd2b84c54ea1963387689c7789dd2cb3a51e113f179e331a16f06e96fd4bf1d1e75db6017464322f2ae2852f095644a6ba83aa37293d16c0c42e607edc4e0f44bfe3f9eb3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d16416c77210b4954b6dfb5c788882c591cdbc0753f6bfc0049356aea9f171bb0b5ebcead96a07d201e9476fec57a1500e473562e60bb7811157b1a0db2ac536201d07a70fc82d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b453a3281480ad8865a4695eb4343d398138917a2a9e383b2708b40ba818eee6ef642db1365ef862cb3de4acb80e1396422dfd58da6c6b0a227f6d365d97b447edf36686760d173;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49b7faad904bdd5e9838617f05763dfa93cd141fe6a395714934b09dc7ab2384cd7f7564fa26bf6fcc47b415b5978e23e5e1418753d689ee348f316d8d656448b6698d1b7ba9f91d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54ced56abc738571f28c38f37df593a2a75892a835f2997fa8e4a18a30d6ad3a619c2f36a77456d7082bbdeb18670bb99bc0e1a47cba217e6c9660b2809968257e6a6a21ff75c8a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52f41d2275d1eb5298dabcb4f08ac5f088393e564697b23ca6008d4e09d9c588c343176ec7980e7786f66aeedf9152145431f89dbe9c20086ba00eef6cb24beecf3821d8c46ba685;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9590c564807a93395d24c243d5f007a2d3d72b3659f27febb31c342aeaec9e2e3bc769dfc5b08c926c3884e459158b6499ce4eba101ebcc0797d658e62910ccbf22c3c39db07bb0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b1739b7af3b155fa8bd675fcc533e8031550ec645a1f2fd35a5a67577e9d51e766933e7d385dae6b62ba4a2513bea9a46e9af529a1a399a9f2ee9ad71fb2d0ee79f027a7522e165;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h822fb1b258fb7a06396268512abf9f77e715a454dd67846a2b1c84bc9b4e87b2deef16deb0104084b54366487d836056ed288338b1639fb25ee4a1963562bbe31cd71a4469a9fa32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76d1c7367fb7a993b59bbaafbbf819c4c3586287becaab237aaca7aad9ee404ece553eea902c8de6297f00cf0135a6e2c4451b591ecf6389a389914c544329ccb4c803e3a8c85677;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3690a1273ac7f9eaa88905abfe6323204e94fe49d9b0a3f1bdc225b52fc50b5d6db2b5a9e1d9323012a434cb75d82a2269af200d9793fc0e0a281b40f030809aebb16d03678258e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h910e6e7b1cc7ef3e05d6cb4d6eea5689e5d61554061234d5ede14ffee7b001cf1ab57c94d5ee3a7b3a481948e2e54ee57824eaacf9f92890ce9438d2711a7bc3b1ffb3323318f124;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38e042043989ee12cb687553d31ee3e82a92ee524265a5628ab2a099e3ce4560111b070e84bb5020d4bf1d1d22c9774a1088c5572d1ffe89f2d44039ca1ae4e33bae698602b40e2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30ac2122dbe9d756bd861545d4490fa169cbf4fcd96f57ea93d18ca645da7e89f5d366613232b46bdb5576337f64f8b718fe4a6ade07d1fce582843c6f1dc285dda23a606c62a7cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h444940046836b6ad169911cc71849be278c17ef985b24e6cdd46b7c8ed319f234137e9e595ab36d9fdcc3b54a6fefe24d07121ca3da4dace97322b4667f8b65b437f8577d8e323f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2782e513a584edef65330b977ecd8923e8a596f4ccfe9618fcf607c64986e0ff8143859eaf934c7b1db8a2c511aec64d7c6352aa37a819ebd4ecc16f01ce584fdff7de747ab73845;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h890bd1841dd6003ea54642ca57a179cd034554e58ad1a2aa481fe912be45e7175e3a05357cac0c3237b2966be06368fdbacacde7d91265b826ae281deccddd919a0965246f2bb056;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78b887b2d5c4f5e2d2fd57a794563e7cd88bb4049d08d14c04b8aa95c5f138084820d9a5d14c2ce9b8ccb10546c9c5b5ca8710e26a26999c8e4e9f3fb7ad82572c9e86edae4bcecf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdf66f80a81047a8df25ac074a3ca8c991a170172a73a3b9f24af1b7f7319cdb65a98ef027794d5cf0875e0813b0e0a8c63a87c4ec09530f5cdc83f9feb79363ce58960ff6d2f844;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he81da7e4bea560d8834666e545e50b218cbf39e4519fd8caabff4cef4d1d6ec9c44fba79bfc3d81d2fcb221c6269cee7794d1d3ca8668b9a5351b1090240364b889e338c91b89d8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0af57004beee47e5165fcf11f0662133471f9e420c59d34ae22df200ea959ce819e6e30a5b16bb4daad2457ca3a7ad02b2f0892cdd26780002a20589f6ded22e957c7f192c9e22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbc1fd54c8923c82db8c9faadfb026dabbd6dea136a6e31fed38ecba694f3d142c43506a92719393c1c7e0e5282d29ebd6f38597655df9e1e1336c2d8a8b786e359de5b744a7ad46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd07def3aa7c28c1719f58482a1941ee9cd6ec921046df50c871fe5d5b1aec52f4e75701f605566dfefb6901c5b938a90da61b2d323cb831a8da93eba153a026b701db00da94fe28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb30cfaf982d7ece820048d2ce81cb9cb8e08e1509e0d45ce9637ecad75600a853d1f4a9db4e6c39ffe07d05377d7e018bc2cbbe7a25f0d92f736953b3e235c7bac4fa9547a97cd46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47bfc73b2c456b1dff12bc3bb9653e379164397912b5bed8ba947a261479f9964c2fa17b6c98161bacfe5c37dcd44080a25e9414a1a1b4c30e1b32b13f2bbf068ad50f0e8b6670fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb3905ed2af04c70780f53c283151e7691ab2125bde4aae3213d38028bea4885646e99de210580d3c1aee02c1510ea763d4e9677ef475580acdb26ba20aac75dfa52b86f0fed8f50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf738491134406e647e76b3d6ca40ff8ca7c15f467e0d2e8a6616db10b5820bf075c14f6542efd622ecd1f795a7623d54399cee478dfb608f0d80033ad18a88735d48f97765a55694;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda2e0740cab5d118918876ba7a113111a5b7e31424445ca33c501a16bab97856500425cfbd469870eb320d601bb734929b0d359a323d69204d2659d23221161902429d184fdefcf8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h606f0c2e98d430935b3f00ecea0dc041d3f9f73e25743ca91fec1d7adb73cd34bca9c27dd4ea5dc3ef924a073d68759879914fc4459d754a30c9ad7a6bb00411a556359d755ecfdc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5b10b115c38aa39becc0097863001d290b0a108975c6fae7434b15375b4ae2927b3c6d3e44870b7b5514bb829cd7fca9c5648c9f3298915ff9ecef8f880edcce622ede3762db663;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafa7e00812c16cc218324e783cff7b146beb51b67b77d75fd1cbc91379dd4f17e294e719b89d517f4e11a33685767e037693cc532be3f6b5b36f90e0835db6fbd52ac5669cf4238c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d9de6b8a0168a20a4777bf8a26d327c2ed5325315f3c0ccecda37af20bc4fb3e386683b1206860200e25d1dc12d23c71a50b002ddd9f9931a9da4fc24e9f5976e95cc3f7a6aef79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde62e2598319ffc7472a34aca56140a63bd534d22c53f95bf11aad5ddc280d74264d7091082ff0f36ea8040a28092939604efa3cd97f687df2ebd433a7dad2b079cf699e4946af27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a9d77a26fad3fe681c68c2d0145e813baa9b5eeb73e29a2bd40d6b908104970dac03c055c69c1816582cb061f7dfe575735c616ffa673fa88c17334eded491a4903c4979363cd4b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda61b4351c6cba60528372dd467ef27f01f893d82ceb9977424ca82bfd841cf7d438c67011f2b9823bda17e9f925e017c119d4984df93b5e69b38676b86d84cfb7a8ccdcedde82b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h673d1226e9fc5308d4f106651bd3258dec52ae279804408dacb63c77ca9bb2733b669dc7f85456304203ef61820f38a8284755c1795b5713409ee89dd72e1179a0aeb0ce226d1efc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb7f2e803f4e7ef7d79c2091c4c9647aba420c04fb777e13086d2155c240c178892204995c28d1758f7d9318839c5a010b56047396cfe6722a93fd8b165ac2c67b83f163c18d441;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4ab83f01909955db7fac0a41185654cc95d6b06b1427fff889bb6cf1b1a825dae087ef43990167b63c86f7a7f20425bbe4e006fe948b9f104fefd632e72be790c46dfa38373a663;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80f6c8a6b39525ca53d6b29d324bd923c68d74913be55bb7ce099bdb2796fc2c02b9ed212327decd6d7f731b7903e625d818efa341adb7c4f20142b82defc2a09af82753440df2c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4be7e5d14b035cea2908918a884910ff58e36b4ca283dee17a0925f6c0ef03370d94c2728b21fd31fee0eed700af764d573c65eb7a8bc9fba5a445fc6d898e060140d7561f915238;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bb5e4635df487ea398a5c2f95a876ac7eacb310fe33586969f6d93d95767f218abc1275a124cc6f6db06edcdf2f2bd0c1097ebc3a84e8920e14c21627e9f3871861924986300214;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6897d91dbb5834094957a177b9e12cb76a05bb682520668618f8a63e67430ae42de173ca5ce121c76fef3cfba0aff49947872bb13afbf238d4f8a065dfdbc707b4498dbb7f04b50a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd78eda7da63442afaa94a4201ced9806eca84dab833dfb0f8e12f1a11e2fbb2d3bacc53ce031ebb89c1cdc6b394c33df311f12f25cf07a9d2c0891c9e622a37fe181ee64765c56e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bc5baa047145a1d2e577c2709d8ef1aa9a557d4a7a7c491076d5083877d02a37c9af36d58292ea6d2242f29262de25b008b80fe42b439caa9aaa62ebb37664c79954580f64566ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h156cd7727ed63b73e6ae986df8adb8f2b40e60eb3169888e297c018fd980b6c41f2ede115eaf328d30aad907cb7d02d18eee62c2c039255dd1bae01791215a1a9f28267aa12c8b30;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ebc553463116475b98e9fd137de62d3e552e6532b2aa7761dc6170c7ba1ce4bebc6cd1547650ebb5e350b84b98fd1d076183bd0764704fcc7b73f792ae84ad953f777d08a46a45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcda50e593e4724978c6176d2c59de6dcc7e539a9f17a04456208b1feb629cf01c1fee68d1b1d7284716b23dbdc2ec5c0e586dd60f08f75ac22593a9da4038220cb520b098656715;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28341cf41e1c292103c9aa4cfa990dfcf6e974cf2f58260561151888c8da6b38ced5f6972120a13cf34abc41415ad03180e9e7383dd8ec0fd2555d0037d2f1c4fedec1417d3c784;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac929345c59873dd7b589fe1a8426a761b2f2980bc6825eb48694443d5eacd4704cb760749444e45f601fc8d7981537a2b0240c6b74b2e9ff4e248897957afd21958050979619798;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf44097ba307fd789a5d27214f6bcf4712bdb0379c059d652b8d753fbf3d226b1423b281790752ec34bbf2c1090187246e4deec4c946a44e61bf906001ad4f10f5acba431c46ce91;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf325fc258b3d6bb03ac6bd9a728398fdf4d204a127fb19ccbb0a8ea8868b0f96102da7b595fee66f2e03d14f4153c4a1f557d8b0d2267dcb09f206a8f3d964b2e783d3a29374bf88;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb283a9da61a5fdbfac9a0cdb67b10d0d1236277b1123e4bb847cc0b0762982e9100eb49d655b4e5468643d33ba4e683908c5fb9b962d2573df54b01dfb82d716505c148ee8dfc5b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h315d3f7fdd7b65967a47b00fe29d1718a7142b7ccb2e34410c5bc7b916f87f886182f7a3f5863a31fb0bf93244961f2e918def550daf57ef21388c658e0ec92e598ea5fce1a0193c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c1cada50e7eebba32aba6e32a8d84a8f9f69dd370917263ced13fe5790783a8f6c7bc695288067011dace16d1699584674b78376c17ac94fc4f02989215e6ac854e5cd81b8badeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93a4b94e76e55fed62f746650c1f814fd8697e813709bebbe304dfdc301cb7a2913ffa2bbe779fa773d31fcd0bc916d52a409ecc23bc8af2cd4742e5f237ede9ef4d84f5f4e93ece;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80107b16253ea4755de4d91641e124734106907782a476717749e9942019bf3929f52a8d2f690f550d6cf8a5457973f7fc4e57488dc06e9d048e31bab275eb8cdba7d3279bb00193;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a3e352fe995db35d343ee23cc8140b66e4eb1fb3a03ed982f871e3a70e4c19d5a9ae2565df70ef5d4b046f0c47153e01a2e6aa0fa0a67758b3e3378016511179b2c0e50d6780621;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h429cc2fddd5ea7c68e07aa34dc579d720e3130e83cc4f6bcb52f4bb5dc4b0f09314da0f2fd8a52379ae61a11622b9afc4085f4d71cde4fe8fa7de864e824211974f2a2444d70b028;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc263f38beb5a17a415850d316f63718600fb4a2aa69cb3f0952fb7c8cc70759b4729fb14ef41dc0e8ee32bb16d6e15699bba2e0be556950b415e9acb4eada1a7b810f227f247e14f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc60fb8dc628f63b127164c962a00eeeb59c709691ef24bf876ead613d9150ac276392670969bd8abdf6aba6b40bd6817f83d5ee2fcf4b3b08f0044da209f4860f0381411e503d8d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76aa2965147a00bbb680c51a42bac41ba288e9fa1f1de935d46dcd9d511bed0546b1484e00907bc4d8ccee3dfcc1b17960bec16167c939ec336b71b96c107f4132e4883d8b69c99e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1106ec2d987cbae2e29f695f6a95af4370d9fc96d4e9c7543da98cc70f16f3c6797372a598be670a64dbec0d3ec71cb09302a1bf51bcc1cfac74b20db0dfc92a9e6f3b9143600c6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ef20228844e86912626349074389f53c8e81deecfa263dc54d5e214880280f3b3161fd4a7ccb1f012bc31dc4c6801f0f8c86f85b9c2e9da555c91839dde941a2be587fc156cb0f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea5dff17f0580e4d8366c5bdacf59fa315b6d68e1d9338d5bee89b9f93b6010ff923f458d7998181af5827061414acf5dbacf04091f1b20a3d3219a9f1fa2e25ac20513a3eaa4195;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6da4988941a37ba3112b6cef8c08b3091889402dc295522dd00b1ad695f86c365931088029b7d939aeb76f1d51c2312f4a84d632b2aa7d0a81fe0d704d6d44480f6338ef77fbcff5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f35785cc039e777dac0c89c0e84c8735d7c2860388d05c614f2cc699fcd7bdd98da309fbdc79feb20df6a4c3899ac11ce83f98d8cd44b58d27f2c44df1a78bce649e7ffcad5c095;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87e80e18284536cec1280494a9a881ff20f0014b1a254bc5e570f2a52e670f674f61b114bd2a4614ab8152fc9e65a1cd568a96e7035ba8914cd647dec69946e50a9b978a0a0f55a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50ecc1bbbabb259dd07bf6416f30b9a63f7621a7871ed3b408a8052f42561a19bd29cd4a1b6626129b2523ed856d3daab4940b40a57e76461ba702c463f809f595751ca70651dc04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd575601d233372f4b6ebe56d893be04e79a6a122db5d61b2099ca6218218db4d2fcf337f9ed3f87f4f1183f581a75dbace88434874a830a141233ed9064d510b598147614cc3c38a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h891a40ac75ca4aafe71c5bf9bd43b8ca1601745509460cccc517d78c9a4b68f9a0eb68ba208938ebe7d99386c52b369cb86169c4cfc99a5411061a99ef961b8a31526d0cc804f106;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c7efe0e4d3770d356ec8768c7e9f5bc2d730c289755e7ab677639591ba7d5b869a171424405dcb02821612f5b86ff0bc0f990413a3fc52e614612c5769809af8d1419427b44c8dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71d246d6b8bd7fc80b328bd71739565e7199b32ed3e5a4ea924e4e5991cee0dcadc12292429944e694497292e9aa72ed75e1694403c5d41c2ac5e8472b4779ffc2b73abc7772d6fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c29fdaf9d2964d96efaec77c0b32ef4964b2728bebcf11624c23a469f49c41b0aedfd129fb079405d890222c301294aeedfbe9aa4a9a4b65841fca3a5987cb123b02c3d42e0f7a3;
        #1
        $finish();
    end
endmodule
