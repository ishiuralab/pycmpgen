module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    compressor_CLA32_12 compressor_CLA32_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA32_12(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [0:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [17:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [13:0] stage1_4;
   wire [14:0] stage1_5;
   wire [16:0] stage1_6;
   wire [10:0] stage1_7;
   wire [21:0] stage1_8;
   wire [28:0] stage1_9;
   wire [24:0] stage1_10;
   wire [29:0] stage1_11;
   wire [2:0] stage1_12;
   wire [0:0] stage1_13;
   wire [7:0] stage2_0;
   wire [10:0] stage2_1;
   wire [1:0] stage2_2;
   wire [5:0] stage2_3;
   wire [6:0] stage2_4;
   wire [3:0] stage2_5;
   wire [5:0] stage2_6;
   wire [12:0] stage2_7;
   wire [5:0] stage2_8;
   wire [12:0] stage2_9;
   wire [11:0] stage2_10;
   wire [11:0] stage2_11;
   wire [8:0] stage2_12;
   wire [5:0] stage2_13;
   wire [7:0] stage3_0;
   wire [5:0] stage3_1;
   wire [2:0] stage3_2;
   wire [0:0] stage3_3;
   wire [2:0] stage3_4;
   wire [5:0] stage3_5;
   wire [0:0] stage3_6;
   wire [8:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [1:0] stage3_14;
   wire [0:0] stage3_15;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [0:0] stage4_15;
   wire [0:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc615_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[0]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc606_5 gpc9 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[0],stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[1]},
      {stage0_7[2]},
      {stage1_8[1],stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage1_8[2],stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12], stage0_6[13]},
      {stage1_8[3],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[0],stage1_8[4],stage1_7[4],stage1_6[6],stage1_5[11]}
   );
   gpc606_5 gpc15 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[1],stage1_8[5],stage1_7[5],stage1_6[7],stage1_5[12]}
   );
   gpc606_5 gpc16 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[2],stage1_8[6],stage1_7[6],stage1_6[8],stage1_5[13]}
   );
   gpc615_5 gpc17 (
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_6[14]},
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage1_9[3],stage1_8[7],stage1_7[7],stage1_6[9],stage1_5[14]}
   );
   gpc606_5 gpc18 (
      {stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[8],stage1_7[8],stage1_6[10]}
   );
   gpc606_5 gpc19 (
      {stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[5],stage1_8[9],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc20 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[6],stage1_8[10],stage1_7[10]}
   );
   gpc615_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_9[6]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[7],stage1_8[11]}
   );
   gpc615_5 gpc22 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_9[7]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[8],stage1_8[12]}
   );
   gpc615_5 gpc23 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage0_10[12]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[9]}
   );
   gpc1_1 gpc24 (
      {stage0_0[17]},
      {stage1_0[3]}
   );
   gpc1_1 gpc25 (
      {stage0_0[18]},
      {stage1_0[4]}
   );
   gpc1_1 gpc26 (
      {stage0_0[19]},
      {stage1_0[5]}
   );
   gpc1_1 gpc27 (
      {stage0_0[20]},
      {stage1_0[6]}
   );
   gpc1_1 gpc28 (
      {stage0_0[21]},
      {stage1_0[7]}
   );
   gpc1_1 gpc29 (
      {stage0_0[22]},
      {stage1_0[8]}
   );
   gpc1_1 gpc30 (
      {stage0_0[23]},
      {stage1_0[9]}
   );
   gpc1_1 gpc31 (
      {stage0_0[24]},
      {stage1_0[10]}
   );
   gpc1_1 gpc32 (
      {stage0_0[25]},
      {stage1_0[11]}
   );
   gpc1_1 gpc33 (
      {stage0_0[26]},
      {stage1_0[12]}
   );
   gpc1_1 gpc34 (
      {stage0_0[27]},
      {stage1_0[13]}
   );
   gpc1_1 gpc35 (
      {stage0_0[28]},
      {stage1_0[14]}
   );
   gpc1_1 gpc36 (
      {stage0_0[29]},
      {stage1_0[15]}
   );
   gpc1_1 gpc37 (
      {stage0_0[30]},
      {stage1_0[16]}
   );
   gpc1_1 gpc38 (
      {stage0_0[31]},
      {stage1_0[17]}
   );
   gpc1_1 gpc39 (
      {stage0_1[31]},
      {stage1_1[8]}
   );
   gpc1_1 gpc40 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc41 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc42 (
      {stage0_3[30]},
      {stage1_3[10]}
   );
   gpc1_1 gpc43 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc44 (
      {stage0_6[27]},
      {stage1_6[12]}
   );
   gpc1_1 gpc45 (
      {stage0_6[28]},
      {stage1_6[13]}
   );
   gpc1_1 gpc46 (
      {stage0_6[29]},
      {stage1_6[14]}
   );
   gpc1_1 gpc47 (
      {stage0_6[30]},
      {stage1_6[15]}
   );
   gpc1_1 gpc48 (
      {stage0_6[31]},
      {stage1_6[16]}
   );
   gpc1_1 gpc49 (
      {stage0_8[23]},
      {stage1_8[13]}
   );
   gpc1_1 gpc50 (
      {stage0_8[24]},
      {stage1_8[14]}
   );
   gpc1_1 gpc51 (
      {stage0_8[25]},
      {stage1_8[15]}
   );
   gpc1_1 gpc52 (
      {stage0_8[26]},
      {stage1_8[16]}
   );
   gpc1_1 gpc53 (
      {stage0_8[27]},
      {stage1_8[17]}
   );
   gpc1_1 gpc54 (
      {stage0_8[28]},
      {stage1_8[18]}
   );
   gpc1_1 gpc55 (
      {stage0_8[29]},
      {stage1_8[19]}
   );
   gpc1_1 gpc56 (
      {stage0_8[30]},
      {stage1_8[20]}
   );
   gpc1_1 gpc57 (
      {stage0_8[31]},
      {stage1_8[21]}
   );
   gpc1_1 gpc58 (
      {stage0_9[13]},
      {stage1_9[10]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[11]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[12]}
   );
   gpc1_1 gpc61 (
      {stage0_9[16]},
      {stage1_9[13]}
   );
   gpc1_1 gpc62 (
      {stage0_9[17]},
      {stage1_9[14]}
   );
   gpc1_1 gpc63 (
      {stage0_9[18]},
      {stage1_9[15]}
   );
   gpc1_1 gpc64 (
      {stage0_9[19]},
      {stage1_9[16]}
   );
   gpc1_1 gpc65 (
      {stage0_9[20]},
      {stage1_9[17]}
   );
   gpc1_1 gpc66 (
      {stage0_9[21]},
      {stage1_9[18]}
   );
   gpc1_1 gpc67 (
      {stage0_9[22]},
      {stage1_9[19]}
   );
   gpc1_1 gpc68 (
      {stage0_9[23]},
      {stage1_9[20]}
   );
   gpc1_1 gpc69 (
      {stage0_9[24]},
      {stage1_9[21]}
   );
   gpc1_1 gpc70 (
      {stage0_9[25]},
      {stage1_9[22]}
   );
   gpc1_1 gpc71 (
      {stage0_9[26]},
      {stage1_9[23]}
   );
   gpc1_1 gpc72 (
      {stage0_9[27]},
      {stage1_9[24]}
   );
   gpc1_1 gpc73 (
      {stage0_9[28]},
      {stage1_9[25]}
   );
   gpc1_1 gpc74 (
      {stage0_9[29]},
      {stage1_9[26]}
   );
   gpc1_1 gpc75 (
      {stage0_9[30]},
      {stage1_9[27]}
   );
   gpc1_1 gpc76 (
      {stage0_9[31]},
      {stage1_9[28]}
   );
   gpc1_1 gpc77 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc78 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc79 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc80 (
      {stage0_10[16]},
      {stage1_10[9]}
   );
   gpc1_1 gpc81 (
      {stage0_10[17]},
      {stage1_10[10]}
   );
   gpc1_1 gpc82 (
      {stage0_10[18]},
      {stage1_10[11]}
   );
   gpc1_1 gpc83 (
      {stage0_10[19]},
      {stage1_10[12]}
   );
   gpc1_1 gpc84 (
      {stage0_10[20]},
      {stage1_10[13]}
   );
   gpc1_1 gpc85 (
      {stage0_10[21]},
      {stage1_10[14]}
   );
   gpc1_1 gpc86 (
      {stage0_10[22]},
      {stage1_10[15]}
   );
   gpc1_1 gpc87 (
      {stage0_10[23]},
      {stage1_10[16]}
   );
   gpc1_1 gpc88 (
      {stage0_10[24]},
      {stage1_10[17]}
   );
   gpc1_1 gpc89 (
      {stage0_10[25]},
      {stage1_10[18]}
   );
   gpc1_1 gpc90 (
      {stage0_10[26]},
      {stage1_10[19]}
   );
   gpc1_1 gpc91 (
      {stage0_10[27]},
      {stage1_10[20]}
   );
   gpc1_1 gpc92 (
      {stage0_10[28]},
      {stage1_10[21]}
   );
   gpc1_1 gpc93 (
      {stage0_10[29]},
      {stage1_10[22]}
   );
   gpc1_1 gpc94 (
      {stage0_10[30]},
      {stage1_10[23]}
   );
   gpc1_1 gpc95 (
      {stage0_10[31]},
      {stage1_10[24]}
   );
   gpc1_1 gpc96 (
      {stage0_11[6]},
      {stage1_11[4]}
   );
   gpc1_1 gpc97 (
      {stage0_11[7]},
      {stage1_11[5]}
   );
   gpc1_1 gpc98 (
      {stage0_11[8]},
      {stage1_11[6]}
   );
   gpc1_1 gpc99 (
      {stage0_11[9]},
      {stage1_11[7]}
   );
   gpc1_1 gpc100 (
      {stage0_11[10]},
      {stage1_11[8]}
   );
   gpc1_1 gpc101 (
      {stage0_11[11]},
      {stage1_11[9]}
   );
   gpc1_1 gpc102 (
      {stage0_11[12]},
      {stage1_11[10]}
   );
   gpc1_1 gpc103 (
      {stage0_11[13]},
      {stage1_11[11]}
   );
   gpc1_1 gpc104 (
      {stage0_11[14]},
      {stage1_11[12]}
   );
   gpc1_1 gpc105 (
      {stage0_11[15]},
      {stage1_11[13]}
   );
   gpc1_1 gpc106 (
      {stage0_11[16]},
      {stage1_11[14]}
   );
   gpc1_1 gpc107 (
      {stage0_11[17]},
      {stage1_11[15]}
   );
   gpc1_1 gpc108 (
      {stage0_11[18]},
      {stage1_11[16]}
   );
   gpc1_1 gpc109 (
      {stage0_11[19]},
      {stage1_11[17]}
   );
   gpc1_1 gpc110 (
      {stage0_11[20]},
      {stage1_11[18]}
   );
   gpc1_1 gpc111 (
      {stage0_11[21]},
      {stage1_11[19]}
   );
   gpc1_1 gpc112 (
      {stage0_11[22]},
      {stage1_11[20]}
   );
   gpc1_1 gpc113 (
      {stage0_11[23]},
      {stage1_11[21]}
   );
   gpc1_1 gpc114 (
      {stage0_11[24]},
      {stage1_11[22]}
   );
   gpc1_1 gpc115 (
      {stage0_11[25]},
      {stage1_11[23]}
   );
   gpc1_1 gpc116 (
      {stage0_11[26]},
      {stage1_11[24]}
   );
   gpc1_1 gpc117 (
      {stage0_11[27]},
      {stage1_11[25]}
   );
   gpc1_1 gpc118 (
      {stage0_11[28]},
      {stage1_11[26]}
   );
   gpc1_1 gpc119 (
      {stage0_11[29]},
      {stage1_11[27]}
   );
   gpc1_1 gpc120 (
      {stage0_11[30]},
      {stage1_11[28]}
   );
   gpc1_1 gpc121 (
      {stage0_11[31]},
      {stage1_11[29]}
   );
   gpc606_5 gpc122 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc123 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc124 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc125 (
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc2135_5 gpc126 (
      {stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_5[12], stage1_5[13], stage1_5[14]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc127 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc615_5 gpc128 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc129 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[3]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[5],stage2_6[5]}
   );
   gpc615_5 gpc130 (
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[4]}
   );
   gpc615_5 gpc131 (
      {stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_9[1]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[5]}
   );
   gpc1163_5 gpc132 (
      {stage1_9[2], stage1_9[3], stage1_9[4]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_11[0]},
      {stage1_12[0]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[4],stage2_9[4]}
   );
   gpc615_5 gpc133 (
      {stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[18]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[5],stage2_9[5]}
   );
   gpc615_5 gpc134 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14]},
      {stage1_10[19]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc135 (
      {stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage1_10[20]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[7],stage2_9[7]}
   );
   gpc615_5 gpc136 (
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_10[21]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[8],stage2_9[8]}
   );
   gpc1_1 gpc137 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc138 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc139 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc140 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc141 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc142 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc143 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc144 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc145 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc146 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc147 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc148 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc149 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc150 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc151 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc152 (
      {stage1_3[10]},
      {stage2_3[4]}
   );
   gpc1_1 gpc153 (
      {stage1_3[11]},
      {stage2_3[5]}
   );
   gpc1_1 gpc154 (
      {stage1_4[13]},
      {stage2_4[6]}
   );
   gpc1_1 gpc155 (
      {stage1_7[4]},
      {stage2_7[6]}
   );
   gpc1_1 gpc156 (
      {stage1_7[5]},
      {stage2_7[7]}
   );
   gpc1_1 gpc157 (
      {stage1_7[6]},
      {stage2_7[8]}
   );
   gpc1_1 gpc158 (
      {stage1_7[7]},
      {stage2_7[9]}
   );
   gpc1_1 gpc159 (
      {stage1_7[8]},
      {stage2_7[10]}
   );
   gpc1_1 gpc160 (
      {stage1_7[9]},
      {stage2_7[11]}
   );
   gpc1_1 gpc161 (
      {stage1_7[10]},
      {stage2_7[12]}
   );
   gpc1_1 gpc162 (
      {stage1_9[25]},
      {stage2_9[9]}
   );
   gpc1_1 gpc163 (
      {stage1_9[26]},
      {stage2_9[10]}
   );
   gpc1_1 gpc164 (
      {stage1_9[27]},
      {stage2_9[11]}
   );
   gpc1_1 gpc165 (
      {stage1_9[28]},
      {stage2_9[12]}
   );
   gpc1_1 gpc166 (
      {stage1_10[22]},
      {stage2_10[9]}
   );
   gpc1_1 gpc167 (
      {stage1_10[23]},
      {stage2_10[10]}
   );
   gpc1_1 gpc168 (
      {stage1_10[24]},
      {stage2_10[11]}
   );
   gpc1_1 gpc169 (
      {stage1_11[25]},
      {stage2_11[7]}
   );
   gpc1_1 gpc170 (
      {stage1_11[26]},
      {stage2_11[8]}
   );
   gpc1_1 gpc171 (
      {stage1_11[27]},
      {stage2_11[9]}
   );
   gpc1_1 gpc172 (
      {stage1_11[28]},
      {stage2_11[10]}
   );
   gpc1_1 gpc173 (
      {stage1_11[29]},
      {stage2_11[11]}
   );
   gpc1_1 gpc174 (
      {stage1_12[1]},
      {stage2_12[7]}
   );
   gpc1_1 gpc175 (
      {stage1_12[2]},
      {stage2_12[8]}
   );
   gpc1_1 gpc176 (
      {stage1_13[0]},
      {stage2_13[5]}
   );
   gpc606_5 gpc177 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc178 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1]}
   );
   gpc606_5 gpc179 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[1]}
   );
   gpc615_5 gpc180 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc181 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[2],stage3_9[2]}
   );
   gpc606_5 gpc182 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[3]}
   );
   gpc615_5 gpc183 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3],stage3_11[4]}
   );
   gpc1_1 gpc184 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc185 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc186 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc187 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc188 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc189 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc190 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc191 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc192 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc193 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc194 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc195 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc196 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc197 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
   gpc1_1 gpc198 (
      {stage2_2[1]},
      {stage3_2[2]}
   );
   gpc1_1 gpc199 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc200 (
      {stage2_5[0]},
      {stage3_5[2]}
   );
   gpc1_1 gpc201 (
      {stage2_5[1]},
      {stage3_5[3]}
   );
   gpc1_1 gpc202 (
      {stage2_5[2]},
      {stage3_5[4]}
   );
   gpc1_1 gpc203 (
      {stage2_5[3]},
      {stage3_5[5]}
   );
   gpc1_1 gpc204 (
      {stage2_7[6]},
      {stage3_7[2]}
   );
   gpc1_1 gpc205 (
      {stage2_7[7]},
      {stage3_7[3]}
   );
   gpc1_1 gpc206 (
      {stage2_7[8]},
      {stage3_7[4]}
   );
   gpc1_1 gpc207 (
      {stage2_7[9]},
      {stage3_7[5]}
   );
   gpc1_1 gpc208 (
      {stage2_7[10]},
      {stage3_7[6]}
   );
   gpc1_1 gpc209 (
      {stage2_7[11]},
      {stage3_7[7]}
   );
   gpc1_1 gpc210 (
      {stage2_7[12]},
      {stage3_7[8]}
   );
   gpc1_1 gpc211 (
      {stage2_8[5]},
      {stage3_8[3]}
   );
   gpc1_1 gpc212 (
      {stage2_11[11]},
      {stage3_11[5]}
   );
   gpc1_1 gpc213 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc214 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc207_4 gpc215 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5], stage3_0[6]},
      {stage3_2[0], stage3_2[1]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc2116_5 gpc216 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc217 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1]}
   );
   gpc1343_5 gpc218 (
      {stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc219 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc220 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], 1'b0},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc221 (
      {stage3_0[7]},
      {stage4_0[1]}
   );
   gpc1_1 gpc222 (
      {stage3_4[2]},
      {stage4_4[1]}
   );
   gpc1_1 gpc223 (
      {stage3_6[0]},
      {stage4_6[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor_CLA32_12 compressor_CLA32_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h12a41657a0ea9292e819e1a213f32f210c1007243d15686740aba28eb50cf05029839581aa18023a4477ddfc6f5ba2c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3e2b8004fa39b92e972bf53229b1913ef23c6bb948424235230b8e3481c325e19300c475ba640ce0747dbc3b69f27354;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha5e3c44ca1c542ff2d7bcccf7cc9bebadae49fa064413e5f87edab217a7ee50e162ffc5ce05aa556e0a26650b70f3061;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd8fa1f203d21963b1aa15be12d4295a56a5290c3caf63b3e1d3a71e645634ae316b5fd7eca48d6301e02605222e5d392;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hcfe7dddcf4cd240f6330f5bb63b92ef5f8c39f714415382e42d9556b25f32cfafdb5ab2b4c36648f481b379960d20676;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h49eb23cc7ace78b9cb6c95e59f0d5462191e589efef430d5c0f3aaddd7713820e7dfc55e296d52b83576dece5a7e1038;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h47a4834772457df509f92744d64a059b9de5d9b94c29fa89f7d91d6ad258e4ce92b7fdfd26d5ccf0be333a24a011325a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd18f93acc16e28423f93290ecee886eafb016ff104dcad4451f7f307b6e8aedf1f675b8ee0b8c9189aff201d8a8093;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd16693bac766fc336690572d9267c9dad28cd81775d83d1c6a013e25b7c67d39c5d8821ed47ff6c0e743285227c874f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd0606cc5a0898fa3314c6606caa59c82da7f67be5e0a8f889b33745f94e532f02882770b3ebbdf28bab8dd71c7714a4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h84a13c2e8fd433cd299c308a8573aba51e4e1ce98b3a463f2a9dc77d8eb9f44b1806b3c53eb4f4bca6de0b57d161792;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h243548deacd5fb03e33708badf60fd4166744f301cd9747dfab60ebcd4e346401ded1661bf38045116f0d6d4f9423f10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h28d930de16c4c63bcca8d2e1b7373379d93891a32ca0c1c12a92d599d70d66a25e7899c9d5ed6fc27c0ea4af6fe4a538;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9c602870057981857b080a7d8bfcdcc64ce5cb5e1bef1fb77e64f28983e0add14eddf78d39c8e1e677d0d3715d7cd37e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hab6051e077294adc823c55230900be578079282fd70c7526107389579aeea77ffc93b3b9b4ad2e423a391b520a8ac764;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hdf97e535bf76da6c64329f6f9e4229831ccf38584014035a53fed03c4634a2cfdfa1d723f40bd9afcecf3af18864837a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4efa5e3359d9aed28ade601653c504038e9ec4d81cb2beb1cf83f78c57a71bc313f463aa389c686de336c3188bdbc24e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1986c93c700629fd74a95b1af18d8c0b53df34133f82f878f428d520e243c72f6d9fca790f67af4ac599b4fae58455fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6434f4fcd8d565ac4b13b19534c472713c69f60d6dbe5dfa4ad65a788f6a5da0ca7246c230a1ee236a7029bf68e3f0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hfd24f894024a1468259ff1288f77f044af8fa2c065c2d7f0931f67b62d910db1637bc1f4b821cf6255b9c41c9300ecc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6aaaee1ac4069f9b88c0dcd9fb01932f3effcb2ca4a334ec726f4c249d673dd1ebe00fc3275118e1c93c7f4c92596110;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf15fd5101b44387ab0dae0e3d8c19f6b36dd1f608a0ca1380d24158ac44cd42b3444eba4276a1d463db0b402973a81a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd44a2c75c16bc457cdbc0496555d76296a25c61b9e6245446a7802f4ce2ee53e5b3aebb2768725bffbc7f6d02d563432;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3effb4f0e584f79a28e293d740101e7c47d3f6817dea375de2de3f6b2b3b54eddfc96aad15e8322f023385c5fcd0c935;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3772c4e1af9abddc2e15540afaea44e800653fe4511d80f5bbbfefed32d1969dfa9af9c729d6c63b4a1d0a64f7abb98e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h19baccf3e8e98f8a20e22ee1e42a2d81f64a7683a3002dfd43fce392eba0cc9cfcdff30e7765e7d8d3c52442c897eb3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h134be7d7e08d8b68c3d7d524bd06c57f6704f0f7f567ef70b8e0924d309af7b7d102f81c4fc37424ed0ffb5503f0acf0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc5990b3f336aebefc991021a72adea90d1924d175c21ff54eee4f87ebfdaf06007a9896c0bff1b3141a880f4d33bf15b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc10e472a76f42f03fa7da99493b7bc86ee76d4485e14cbc8bedfd45aa305be685e61584dabe4f3542b4e0dce2fc9703;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7ee2da67cd08dcc87ed144cb77815431d9b8174eed707cb5c795304e33921a22bb41eec64069dfa0211b1ab47ddad42c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h48a07af024ba7933dfede8c49ffe3de6193296e2e89a7a3dae676c644b333edff50022450dc02a51a6a9b260d9bd3c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3c29d895e94c88a852c93a7b3aba08161200617f344792a1e19e3e71289e5c5e85f856e3c859933ac0a3280d07670621;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb51cf8bc6554cad67d2b77ec8fa1c95ebe109e2f16eab33ca7ca1b250ebd74ddb7ea0c49f55c3503db7c970c3db7e982;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3629143d48daa3538b08680bfb7bd93fbd7976ab69038a75987897a902189dae6291fda5b2bd37a0b1b479ada8a08027;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he79d21e521f1704d8f92d77c21e69b18d0aa37941dd8bba1daa024060e64261b2c50ecad2800ae39c7a6dec961fceb47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h17ee1edaef0770fc39bd2470334a654d5a6ccf88bb207350014b11f6d544fcd3c5be85b751774f37f7e65dafc2688a21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3791d6c21cadc6a9a6f28e21daee8b3ae4fcdc2f3b0bab7958eda52947caf9de46234d5ee108e8d7562990bcacd8363;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb1a9731b93ecc9f99d0eb7af989fc9387002b795d5b3733527f9626ff9116af93f2d1998eb989fa31f75dc85b68c246;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5f4a45cf44db0b685690885528b2ea8d174d18d427869a87e24cc001650ea64e2ce061d147695fa170d1214d49e1b8f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h62932050625469d5e621d985aa291969c78d97e8b2ef3cd72b2517a186bac98110668646fc8a402fe530f4d3c06a638d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7d9ad501fc5701e885298cf8a588af5bdc4f6ced71e3bf298734bb189e1320e11161fce59af980e9c2e116afeb338be0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h142980c23540e986a7ad55e36b1e13b1942069d76e0215f01deca62c1ddde8e97197a30282b8c83a48fb0b371c3889f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9f271ee408f5c6d8351eb4844d50c0048b3a959ea53b5c85c5ef7d42b0bdf301e1a91cbb018e8abf51d2baf944a8c0ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd1ff1218f23acf0d9b8a7c1537287c7d0aac57eb6e7b36dd71ee69aeddee6de0397d492c0e6176cf2519040dbfb64ecf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb6d51c1a5a62ce5a96ef8f6d683e13df80df3b107b59320fc3c62023e670c3a577486393232534771e6a0569086f6e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1c18d88dc067c3b5a1698b6392aa849467fb53d8cd890c485a70af19a8313933d7c9b2d5331bd816b7ffbc105975fa4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h56ffd910d6a13d831461c3c9d2466f742fc3a12411a3f2e7aa313103649f5d72465fd294c1e112f76daf064aa20f69a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3c978875ba10db5845d3a38cc457a00f4f5c6bcb387d183d96fb5400087ce2b6a0079f4db36f12e673c0e8fe07c0636c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'haccaabcda4e4c3cccff6cba69ad6aed4ff876cc96bf8b35b40ced7202f93d7a39a483d75619144645fcbec8c82242f5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4a2109d36ea14b10f9f2c5c0f98e3625f6da020c951330766fa12f7b170d2bd4fb4e09210e15ed40fd4728b7c70fd512;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h61a789ce9d152b1bfb0092db9abb6683d3b05f04852f21421cdf2c1b8e5a63133d5ef7df9ef49b4b2a7e528bef0f0bc7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h24702c57a1d19b42661c24fcb02c9edbd0c2a3ca36ec849102c31b3cda375dd5b7270eb8e9cf6a47f18f160e6a7ae4fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc6d0636c481a3f9e979ebe1fd65ddce43e9066c80fdfa240daa8d3e09fd956875672862ae143b0d03199259c0645c5e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6c26932bcf920e84b0ded969dcb08d2bc916fa5cbb58504969671c8bd288b692b844c9a64d31f18a4347343f2c62028e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc1007d9ba0cc56c065eff2dde4d1fd9e81051f7a9daa0147ba27eab17af26cd63c919e095db6bf3b3fb881e7b3a84b2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h600780dec18f8bd6cfa60974c68cde3200d07ebc4a350c4dde59593218086516f57f2842a764e335b9d7b74a53cc4b3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf9d2cc5f047cc256ae504f305694c9661615a17b0a4b97c419bf43a3e98696c6505f53021848da28433a284da052ed6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf368c57861d4e491694bf6c2fa803b6057cb074fef2918224e8f8a129018b45104d9c3fdacda81dae193b42001c2dbde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h91a41b043664a26347315b804b1bf2c6d895a280e97b1e7def1b8f3414efd15e0d8ffe04818ddab7563b3ba799553ddf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h374131f71153bec2ed822539e251d8b4de8a21f14d15dda7b7277b9575b2e9dfc2be45abab2c21c3eeaabed0842a78b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4debdf047ae80e064333b3f5345d29a412cfe158d50f70e6b5b8e17d850a96377e6b1a509dcdcf7c5ccbcd31a833a309;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf80a191a1dcddcb27523f6e77846feea54dd4e551bbd258c1e4cca9207b371993d6ad20c31dc1b495fd2a2ec9509be48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3f332e92c6bd7f4af715960866e51972e15ef13a4123e0b9a09ca1f5f0b97d2efae9a3aa4d0cdf1d30f20ac21ed51830;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7165321cb60127e46d19cb197aadf0660fbcfbdce9f6fb597322d55d45bdf72ca62ea33f6dbb77ceec8ef30f1922ff25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7e0a6d41d6d24b90443b188cf367537ee579cf47b2c2717a45f063e4dd77c8c3e1cdd41f6d2efa0f2da8d4823356fd48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h39024eca8ea0d3fce9dbff5da5824f03685d9881090dc20cdeb429b6c10525fd1e8093ae1d01ccc31b8d0f99bff5e7be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha96ccc792b576517c4e25e577d87a06049a4634fdb1001d7bf63b83688ebc94b466a2a38dbb49d6e3d04d5ab3a16853;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd6d2335401d378adcf6c8fb18d8049738db5e111ec1498273be3041fb42607455acf489bc785ec64be0abee2e15eadda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc508d77c4d8f259df5e457db193795925d000315be2ecfe8ad1c51fb3509605299e5036f5c746538168eef63e3738c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h61e97769379fcd9228360ea1600e4fd93924297af789aec029efe41272a1b589881c2c23d92ac0d67958eb3ff13e7b4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h631e2385d56c22c9af562e5fa96a6f2be26b3669d8c11ce3a6935c891ed0372f60d78ae3d3cffbf60a7358d1a794e612;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3bb7b1994c9e2791eee8653ac122938dd12656fb1257b1058f0a99f95430975b9568e3b3810a278a3662029e2f884b2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h12025851e0708350a25b2550668c6821f64a66f3ecf3882abbb421eeb8361b8a04dd72b12446d846a0017b5a431c6381;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h45030901eef06f053a6d8a41262355d0cdf8081b4371e33fb6f0fb988b2dd1fe3c7c00e44af72c65b59a3bcb2dc8f977;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h69fdcf1c79a950e655bb416ef76f93993f2222490ea7d20ace694c2df97294eb0d33d7e638d4c136c276fe1c8ea26dc6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2dd42222d7b0cd9e539d45ab1e97896a465ba0af36726903f26e7ddacf3f1fd47688fa2cf2619873166890cc7775ca6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h934e0ac63d68dc7b142c0a363f6c17c932915d2e8c52108d97eb4cb4c81a381e7613dff8d1cd6c9c25c974723ff7695e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4e3a33caf642065292c43806c2393961e32baa79b5cd57ce1d007d97e13ee2396ed09726b6de18d0fa32e22d5e15fcf3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5d134a76d1886cb93c482e624bde47830a0bd5b0b371fd1fad66da1e76737dd65009e75cc71f06aa9c311b22526208ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb7ae042bcc57a1f6c4cd610c90e5bc74452988c5e8c8ba29183057f4f6186cee8aa8e2e0af0e01dc178932c588c027c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5f32f1fc14aef2d7f26fde71df58a06871d5736e676785298a1b488c42f33752cf084e9c870ee86cf526fab7e89df2af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2617f6c5a41fa1e52a96570f2a1cf67f49fea2030f7278c6512c4697e8557785921ed89c9dc687478e4ac6f5ce0d0a8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h14e2336ff7b7dd582c84257f158898ca1f2f0eff8f7631df86c5df880f76dd6caa471cfb97a3fb7e45d4eef3ed44f1f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h23552a5273c43e7856c411e1f87918624c39a71b51983d83d45ea402e5c08a46e85c1b84c9ec792a2f16d3b830709d18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd80b811f4d3432845299bd6a40644debd5efa20a193592479924f7fb5cfc7be361cf38e1c0e9cd62407e0883278940e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc31af450449cf14716364fa7f51b1e03681e869d58b8462c05bb55e89da9d4a799894d9367863e7d140d9fba8bf97b88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hdb7d9830924d1b60d8fcf952cf3449518e8e3962ca953e37858fcd727982b791daa178dbfdc0765a70a9d70e97684ab7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha12a1a8cc9e54ab0ac5add4e7ee1d1e650c1dd047150c6ee8e208b9d0c5448bee6c6c86f2889e2285aa84af875604d4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h97ed0893c9f55c0b4d5f768e4f462a5213a3990867512655f5c3b13e8549674b77b155b9882db5bf88374da530400f08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hdcfa15061a9d533f8f1fc3e8ce3d7cb20a37ad783f9fd4c46d8bc0f4713ed1b2f886fb4a3e4ea6fe4a15f57329ca681d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbb3ffb72bfd22a62828c8e8c58f0bc9ac0127df3e1f5d9a1aa4093800dd68e29cbaffee2ad3a46b61e0083e8e0fc03fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8b7291a2639fe5d910d3c57531d43d6f9668b75b65a9a34f2b87dc0b31606305d5dda202092cb1f1c9c4b713d47a33dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h38efc78345b1c0d8c1c9c308cbf4955495aa41d8252138612bdd5d87f54f8367d2c3c756b8398d4ac73f6d787d9cbbc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc8546527df484ad603afd137770121659a63f44f403fcfd3c77690aba6c06e39f8d100d1452b3ffaa8a88428c45b90bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h81bab927327b673b504b10aa90dd61ee2a34cecc3122ce874abab1f6485ca39535a7e5642b275feef5b73314e4c2e76e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6123a9728471c6dc08dd08a00206b0741bd6496154634e34523d937aa0ee00593cc189cec30b153a74c003d914512fb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'haa290defa547de9a781d1c8c79e3009f6fb828d95e18f628c839056849b728f0788fad15c9c819809b6de86d660179ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd8655eb53608ff11a7e8009f73bbe5cb8d0de120cd39b37e1f8da2cd4ecd73e1ee62441a18efd3d9935cdd26c3ebd77a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1aa9f8bd6482abff150761b9777e225f3557f1cb850961c7654120742b9c08d6beb17f972d1eb07cca2ae1dbf96e710;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc0e200e50f84f95d3cf3167284e4b7facc5e896d4cadf78a505693dd14dfc40e98b0de307d13cb560548591df0e3db13;
        #1
        $finish();
    end
endmodule
