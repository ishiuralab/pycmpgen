module testbench();
    reg [26:0] src0;
    reg [26:0] src1;
    reg [26:0] src2;
    reg [26:0] src3;
    reg [26:0] src4;
    reg [26:0] src5;
    reg [26:0] src6;
    reg [26:0] src7;
    reg [26:0] src8;
    reg [26:0] src9;
    reg [26:0] src10;
    reg [26:0] src11;
    reg [26:0] src12;
    reg [26:0] src13;
    reg [26:0] src14;
    reg [26:0] src15;
    reg [26:0] src16;
    reg [26:0] src17;
    reg [26:0] src18;
    reg [26:0] src19;
    reg [26:0] src20;
    reg [26:0] src21;
    reg [26:0] src22;
    reg [26:0] src23;
    reg [26:0] src24;
    reg [26:0] src25;
    reg [26:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7a394541c21ac2e38a1cdf852a69f2106dcde82ae377ea93efd78bdb6a6bad47a7dbea06722cc83087dbd97320632c633e5607610a8ab5ac3a2afbf09dcdcab930c1bd74dd883f0f75e11f1ec2ba96971f5de31faad875afec0e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127bab552d00eaf0a9a0cbbb0ef8a0c031396aaf28d78b8dbb83a2101ef1362020475c56bc548114f50e882c9acb94381a5934126f5e274e2061921c68a59996e24f040e7c72c6ef5c707503265fc74bb873f423af72cd7465558db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h571483d5b3eb2ae181ca0bf403bf99a05ad32c4def772e337a15b165e5d89e6aa755f8bb380a3480d81592fa0c934988c31c4c1f148eec68bb953730d2e0a85dfacda14c9c02eb3d42144160ee754a25a96c3ba7c9c68a984971c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc87659411c1ccbcad1b543a623bc298660d2141bf10c80126deeda635eb4305992f16869d4e31246a890e77a8e9b1cf5a1e15c652a00bddc284ef3e45bf3444ce2a28cee39e63d33c18c5177de9689b98985bc127364c857e6a8c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6d321c6dfd44f5dd740b83050f494b71098fba8bd9dc1057eaf0e4520ec8c1fecd8b44cc1b5a706562d78e7bc1bbe58d35e8c2c8e894d6a31598f3eac648fc861c2437d48a3ab50fb8fe794ea955a93d37c9c904df3de4471a369;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc08bb56288410e00cb9afa0f869e0a294b75eca33804b1e7c8e8ed450fa5c0820aafb79d777e24dbc8d32d01f7e114bef2212d3128ad4b6801955d59a36c0053a516c9150156223fb703bf8923e65e3dd6a39384b7eada31e34ba1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e49eb7eb587163aabb51b7f3a769c21f74d2526a9ebabe032490926ee72eea8274b8f7c7fcee93a8a4edf08751db5d06d7830a9419b74bc2e265d9fe445213e96f3e6be0001affa7f238abd6a84785cdad835a82976f05f8a47b04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf1cd96878748297de7331a08821b184144d3b7aac8104595fdb3358261651156e71c0ec5b637be5d6795a12b06c4758669a788ecd4b8cbec63a33727e30bdaa9ff904893a9c2e9e4b4df62bcd8bf3bd879c9af74f096522b74c39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126277222e309700677acf021c7f7691df8b1f99378696b893652cb671fed9955833cad0e7ee54396bb06abf934b162e538067958861e4825648adfed41d932cd87ef8bb1dc829487c278091533e7b930a3822813a59f8393d04b5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb04e42b5ccca07c4bb7ea6ad66d5c7ec456feebafee50340bf62f2b6fc8a301f1307ae237b699a69fa4f22183d5cd422e92da9f638ef336e59e914a1ca75de5dbcc3e0ec31d15cf99cfd5f7f3b04a8fff7c545eee0eeb599565d80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c714cf1481697b20b1bff933b4d9189ce104b6e8f1d1f1c6e59f3dba49524bdb1d27e5cbeca9fdf186935390774c1c8d809c408904a44021db643c0ff23501343c61ec53ea4f52bdeeb86f40b960a01a9f455a54d62926b550e69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb17c687c7325d7e0084939669cc5ecd21008a1e765d7182aba9afe54ab5f980ff92ff123f752d8b9f563f7ff5705309149553fc1ee3509aede8815c595f5f5d232b66d188afaa7a6ddff01881ac155d0a5d58f7fd20a48f0d9e102;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9ca7e153b61c6587c8a32c890b2b6722e1e60ead561fde94a08f13acd4ff00465718cd71a0a80d8c5c0e54599876cdb6b1f48690a7e1635295369d25339ffa5d32f4026b182797a94818938e885b4f7f19268413e3dc1e7545100;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c7c6bf2c559a682a7bdb59a14bbc56fc3d8d6b01c6ca6d3dca04db53a0ab9d5af50f5725db4cc0be56733b7e3a191fe5274d1ef380016d1ab4ba808a9275b4460796896d8924fc16a12297cab9f3cbfad742f924117d2e55dc937;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24b0c264bf120bc033c824b054593dcab588ad83c068f970e070d723c05fafd85057552a8d849544c32c5b9ada95bd2c47797627953612075880d0b4839fedb79a9e30edbde1c3732586865b69328c8d0fd623afe34d2ea9a79d6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d2427702a24ff42c482601d730cada43489ec1fdd6f214fe22babb1b82b21d683b728f5cc4b6ebd1a614cb75dd4b1c331e779943d608675a17e254f7511845d51ae1331e7156ed7116c98509b638b4d18a5b5d7a77e12db8edb46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197f9769b145c4a3d2f1133aa240b79ee8f73d3c875911b1f0499014ac0b0c866d707fad3cd75903c27598f0a6541c21e49289c96ce5a96eca8323f26e87cd4fc66817570bee8adeb869cd36d6d7cb77210368b2d035be69b0c5326;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf475f3ea10342aa09ae7373da9b69327a364ca549f0995e50b949e5db0c173c71b2ac0b032474806ba8effa30fa7ab7b8e88c7c9b3c1d6994bb5384a56a1ba264c86a03a619805de37b9025179734c4abb896ea16bb980a1532fcd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c7d40974e42812cc649c76a8c7aa6f659e67e28891c6aed3191c20f70fb162e6739aab36cc1b0525b933b42f9f1f348c5ca3a519e66ebabad60cf35404407a83a02c20d458aaa18dfd48c3a315fb1640181661f85bc0c0c0e6283;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9452b66eb8250876a1f2ffceae3d216b709569763ecc27934016d88af4b1aa0c0e272e7e91adacbcb81d504746c84eb3b1f9f5563ee168386439525ff42b4a34ed416ff0fd92f75947276ed042603eabdc9e039a206ddaeb533d0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95a12d92efa27da627d05ee69adc4ce86de930bf88dff3327479d86242665676338926c6b6526973f9a7505b7d25bf1a34151ec1f0e5f2d3c92cf8bf2c0c7a79ea1c346622d503b79d79981b8f775f847a4b0367af40c1b2e0899a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afeaa0ffdefbf3a5d58f53548c7fb5b640cb7136002b7201a015c19552dccd999ad65c534498c95537c7dfecc9c7eaf52a8398a73ad05f7c5d8a24a0046b4e092537ae7db0cea567b76ab9867934e6f80e5111ee7896d3e024bdc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183d91e2e6e3ff09ec624c7eb083a1889972be1f0da4b6cf09d8d7eebff664c9817cb7f4151cb2a1d493788a833fcd59aebe3353134ba2d3313e754f3d3122003cb38d977f819fd5268aafb54eb62c47fd3ef173c08a87ba2ab0c28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a74e74677a93e38dafe4e1907a0cd2784cbb7c75155f1533bd03aabc80f610f0eccc833b183908f0f570c78fa2f8a2ddece53b4cf564e7d299050ca411021b63dd6683c19d3a8e92666f5884a6fc45beda0113028f864cf97d9491;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0fbcbf2fed09b11e664cf1e9795f6aa6d1908c7b41266bc2e0493f5b79fd970e500ec44c6ab9db6465b54a22387653065ab87d36a17801db0a820ea749e7765dcbdeb2477b091885cf6f53d6489b1b94e6a23063bb2872fc55bfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ceb7df4d8314af16f397cc932ffbf6b89648ba4c1a94a4024c233c756606cd6e3c0c4eef9aac6495b65cbc1e29b22c83f625247f9b93280ea6d44d5078f7f3e36f95e983bd1e82bcb66242853f3616e7566e0d5a397e9148bd2ef1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e4989a92170dc321d1abaff18806e923d669154093cb4870aac6b18b44e6c86ef1fc0d5d08bb49c967ce3922b970a4b60f6cd5e9d8735278e61d088f4744da70e2f92d771dcd8d15c7065a28e5daa07b7ec4c912399f1a75cd5ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfab2cdfa6d7f27733037c5af9fa7be17e847fe5f077af8426d9de105855751cf8d6e3aa6819b417677f0ba0f9d7108e13a37b5bb128b31d1602a7a46247c70fffd521fafa590ea381372877a86ce5632bedad3fe8c86678c5b9c3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4a9cf9b1f5806e7b9555ccee4d5e63766347d68cf1b3bd0ca6aa986abd905c4c8e50c387dbe8556d74ab671b40ed322029137e8995dd8cb85b61363999a360a32d7fabba9494f56cc1145b59f34f4827b1b8c898aa1036a3a162d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4cbfb786854cd4467d7c05354dd12cbd701863738df2bc57ce0b5ccae22e65d6172a7aa4968080af3f6049197c7fecc64cc78ad5889cfce2ecb00e6c59f2c4ad801ff06ebe25b5a681211e83686b66d56c17c41bc9fae46a123e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1b927d76a28681371adcb8e228e97b7209f44d7be7516baed26fb870ec163b3de294002be773b14c8a618ac069c8c921fff78f742714867ddb86323f9a364feefad1ad8e24414f762d87242e361ae1b72621f3bb7f736a57b82ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa7d4d7c7bd7529f980ac19645ba9fe541e200876fae03a3afed8a32e4f69453b7fff177258c57d9f881ab92a2483da12fba3345bfef1a8b4cef2f0dbdc2db9b9b04567315e31b54ca925fb37727ddf4614a54dab3b9cb7ffb3412;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc129b7a9ff2c0fe7b2a7f07031dc2c49e75dab2fb6a2c6f03edde44dcba2d9afda779d4d517f8c538a9491485fa48377364d8d4d2ec0f6cc1fab464b32b23dd854877f6f19eb62c025e72e582abb373618cc625e3b90b1fb0bda8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bc1231dc679ecb732fbee590bae357e113f7bcde9f5b8efc8809d766cec24a97ba3733df07b705090bed9914816b0f3faceaa0b2069b7b9d53656890437eecd14deecd9675056a669ed06aab1a7768307de8f6e6bd2bad90ea3fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12132160551ceca6eb61cad41613c6c56184b5e347d2cd90a9c72d6e8a221af081bb72269c221a6de40493448b566d2254aa56296da04bf78d0e56ad0368f986f9fd18a32555f50b4563e3ba8e7bf15063c6f6d6ee3e8b87b225256;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7aa87f6cf960ee4cd6f21dc00a8db7a2795a7472932557a0785017465acc37f4c0b19bbeca90a1c0b354c8ecc883f9d1c8c2430387182c30e1c4ef1f3ca4aacb6a7e75e8ba546c03dcf12ad070be418385d450590914c65e8aa36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f218f5c98c32ea97fbee0800373b764d813404eb2e07fbeabf5ae4d488a395842a87e9fea530a39cf6db0c117bb799744892581d36a503fb114d3298b036a126c84ffa9756e0d7a984d75f1710c85fae24fa2b20f7f89dae9ff47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9a74822eac9705f528d4165b71dd0fcab30682477c8803fbaf3bd10ef3c4c781392b02ec047429f53d9cd15d61552cc32689a09007bcbc557da7b247561c9a8f1e4b1f8a4c90d4e9b5dce734971854da3796d31c7dea39a675a2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187be56ff4059ae370bea6f7447a570fa8444aa1f51a04ee9258d6d803d873ad9c9795bb009b2fcbf11b35bf2a783df48daa28443a623c6d546b71db0127f6f1367d8700f5dbbf9d6476730171abf1fa5429ff7d2032cbe15027ef4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea3bea8bfc971036b5e1a82688420a235d5dc7842bd7f6c4853b806873c62ebad7f27fbbf864072e3d2e6240c5822afbf1614043d79a29eeac3e7242171843ab3b7e4aaf6b2eb9f3f7f05bdffe36ef83079d16e5bfeb142276f146;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22772d8bbd44edf1c961e99ac0f11091c91b161a8a68b62b303d9d25a160977d728fdd81a70e92e3c848a39837db739ecaab4e17a78d3062c2e010ed883fa86f5a7d7b7547378c77a61420645fda58b9bd6caf28c5f842fa062d55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18aade397e705f8963e9c76b0287f751843552087025a54b02175c0ec743559ac2b48de38c4f36aa96558b0f3023a865d7831859490e24032e837c8ed3694227417e0c5ce950ae5163fd6607bb95a9efebce626b48a85cafb7f4f92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf709ac0e7111975661459b675af4717815451f20c16c4a685eb7090b0e27f81be4db1efe118580b4a21c0fff539de726f237d5e866bc575b6105a3e309fd356f96df89e1b266c6df43bd8a6bb82e64382313da18680c9dd75e52b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e36935e7fe5fd6c8de1eb3baf7740e7841f5c1b15f4130df1d8807a415446bfce3a4ac62a280512b641163dcb2dea404e45e4177664f3b6cf4c28428ea831e33879fb742a6021aa5e37e97d14c2441fbfb967dc52c07c58ba9808b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14edc41eb62a63a6ac4a6577418e99fb61c245b2bb4ee911710846bb116f83c78f97bccb69d0b6222eb32dd2b37d4e2206e3296efea091eba8467675501764381a124d92ad578351340ea5a0a9515d84c9f25ce17529e13103a047c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146065a9cf48c8853bd03cef6223da9660906b5c00ec32abddde1ed08ac3adc9aae44a3c0cb64c9d912c2d0459461b29c76cdb2edd6e3873e446c3a04e0d3d272d8bc8fee3138885c69cf98b3d140d2eba04d211805ad83b1f1c8de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c88e9d0844855e598931a87a74303698dbc84dd1659ffa8ea93d4e04f5ddb1ac9d12492018e371677145f5e12a13858a38252176047ddb50991c8e02e44c817ba94cf6abb4ec2df693c51018908731d2b73bde64eaeba24e401f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd5568deaa77525bfd619230bcf92c53725aeb8673395bf9702a409bd84eb7c32cf76fc482f83b05aa50b53b78bac16b12c85f96d519dc3ee227ba1dd08f93bc43f0d3a460ea66201ac0779d2d3af0e1b4041ec103a77c50d1225d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bd767fedc040d239c38473f00fd0e08d62df191ef54a87e3da41031773ed7f39046e5dd4bd171e84d14e0c603f0a0a723bd24598905785b7be25862466d00f0bb10975acb6420f0e5a3618abed37dfb5e5a9b57d557a3388291e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb947597b5607e9f901f79b529e693e435102db4d6a8ca74d5a2399c203a9aa7e6002dc72324dcd2583a171345371d050ed7852978bafd522b13de32766b8abb18d28b06901ba8f43ac583efa48da550d144e8019c00f8d9cc911e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1932435717f5626db945ff8af03fc83506279c4d338687eee89b7a45d6af0c92d6c725059ccb62db4c1402a09262fc440b2477116007cf05c3022fe801c884d29d3ffded58acec9f9ee6696d3269ce84c1093922ce2ded39d1e5f21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc30e2ed94e557d55cf7b60274c6abe68801be77a8f2264b8d55fa5732cbcd3702d15024e7afae0150add161937619342eb2fb959cce65b7be655f3ef4a8b526b49ebb40281aae259ec882580968212887d11e45fb0f65e1d17d0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5b63e8176145dc569465ce8d80a946659b63cb0b68c816e676f7b092bcbd1b77003f14cdcae06da1ab060821dcce20be3de0788ca2df544729aa1eadf8a14cc13f255cf067689793a0f6b97cd03a4919acd4bc460dd196c575ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf810d63cecebe97f1e7a644a11a336ca06e5800e2450878358f192a066f3c6c186ab5895fecd013099656d9073a8d64bb68296c906b8fc8f64f60159c31521ed74ffa7f5bfa65e5681f56daa49820923be42397c15088ac119966f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148db0cb1eb7a17eca856c31dc6001eff802dc0ec53b090d73de920d7a06108300f9b05da97576e2822fa0c7987424d16bef35d0d39dbb7a6855a27efdf96dbc7af5201fcdc9b044fc7e5d9797feb41b56ffedda7d3e738d3446706;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44e0ed8cef190d362fb768a8b0ab8ede2db02fb26f99c942aab20305fe54a1311e223023ae6906a5dd6b0a6f0e2793f8f7b0d7f8c9a02b50a0440e1b692afc9d422b9b73879e627a7e1858861661e485ce98c1953dc43fa3f26518;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc16a69bf41c2b8418213c29bb5925c053c26f50800315c7dabb847ac99a0cf42702ae6f5f7e0f7a67274fe90aef532b2e1be4b3a6792b76bc5c0084f2eba13febab58bd50878ee340723c928993c938510d2fc2f37cc8fc9acdd4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a883474f439a5310178618d5c60c3b17100bfeff5256878eeb37c9ba273f9e84c0bcd6bd9cf44b44beaf4dc04bffa089de98e6363874279eb409fd7b66becd58c853f5ff69ab0c792b6f8d1545f38f1b155b977e7ca1b6bcb2ce0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da33b45890fb482b45d4b6feb27df296175d1bc63ad29df7e19ad0ca017e61971ed6af696e78010d2bb3babff77cd04c349c2e9ba0352f4ffc39385163c4109ce5610b8d71c5e9a758068a174cf918a00864d7752dc5dae80b7aa6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h721b12c30de6e3330e5b3602144f55e0a7337b04f13d6f8d7a9dadc7fb552c0849659e8b42b19c26404912bdd2c8630979f1539a6aef89e8bf0385ae11f8f9fd217ae6f328af141fa4def276c2fd8bc065ea8d79bea40dd9ab76f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c02368c4def99a06c88a47fb4a564275b70ced75c762f97f014c4eb3740d0ff557512669033d07432ccd447a5c531edfe26ee8b65d21d38fbd3de16f5e398a2bab16b34f3aa72133e1228e39e883a9dfc22f1299c6e291483ca20e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153c45c8daa6d6f3d8754c80d31214bf63e2ad60efdd09662282ab512c5620b2ff95891ec7533d5facbf90b49bffdddb4ad9f4136346d716ed80f9ebf08de7451a67a87e76ba6ac342627c1a703c28ea56c56973ba8f90a4bef532b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1d4cde078c3e9254f1ceccd11cd343dec270a302674f107c48e8f86b0219704f7e9e88415ea5aca7af7c81340a2327e684928e40ab2a95b98d366b3fd1253fb08cf536af86b8b84538cdff3adc004f0295a6a501d348b5f893229;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h138e5a3ca9c1cdf711b8e300b51cbe8160cfed4d95b71d79749255bb6204956f444bea9c61b1536797f153a20af98b2084527ff69fc37faf83b58daf341f2289dd83527f077aa6bffae22ccae5ec7e612007f23df755bbcb57089c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h859ae2f5d8654c327b23184e4db9ed080653fb211876983711297f9c447b642d46ec595b94b46105d59d27abeeb13fb0ca2b96923e1a0ce5639c3aedb931b3db83397fbfa174fb60eb795ffb9655e4de20c7029bb5b2cd58709f48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a6534a9c41ac3427b98847f2f36fcc51673dc0b1f1364eb75becc4cfb45d8cafa4840a4f15d2197b13e1abd28785f4da8dbc89f90b74d705eae39d8542ae113c44f57f09a34456db55070f93ce8bc0a5d5c3df51f5c4adbf4fe8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb47476f5abe3ed3f24468a7eb5254759d1659e902b9024f561cba5d10b8356ec34df1e9c7a68d0fbd8fdbd77756b6d6cf6afcd7fddf94c365811ddf7e06b9453b9af66fa075e60a02e652d0c4e40ae95aee9287fe4e8eced820b81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115631581cb830de79ef5bb7434dcc789bde6859bf09349c777f701a2bbb31ab0c7e26f8ed51f89a4b8c65b4ac0c0cda9b90a129bb3f782d0fb417c73f10fadfd26c36c8f96661fa4db4ac92c1fa9d551e3775c5a2484645e6c11a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4e85ec9c25acc3a0722c2aed5280f4288ff2d0524e438124ecc41aa3c3b111c40de50ba70cdb89b64633290ee1ce34dfef85906c97e0259fe24663f8e08d4118f3d06b7184f364d923c04bddb36cdba105fa25cc4fbac1fcc126c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1372641705c6ec83bbf99a9d7ea8d2f8bd1cabafbea0b614d3a8b529e06e5186c6e119f4ffe23d9f534577b7492e6347a22019ee13cfac863719a2ecd7ef18d0b16b47cf396e30cfaa13ce11f5a9ad2965e37000ac293eedaa308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19710fbfe9d1e49ada5b36dcfe0dab8536e1e8c69332d9c2e029602db1419bab7f3f487d05e3a4e5205e2fc2ebcfbf78f2c3184c80d400c23fd6fcfa6ca666d0387bbb4fae90c8a4562968fe72180902707642440355c3b87abf5ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31ade2b667e099f0c4dab063d51b786e75fedfddda83aac02a2906891de71956d93caf5bbd179ea5a44854d546fbe68127d904b35bbc63938f3ba05312f8eb826cd21640be399956ed0502a13c3aaaf0bb99625d061c841d922946;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c4b01cf464a1925a15b2975331c4e23e024c883f85c99ff96ab8157f8d6f470e56c4221e6ee41f38d0bff39deb1c4249dd4f7129293f413ee68554bf11a84ca5bbf1f127d950d8b1cd42256ee4315fdfd9b6fc8f2d6f42fa877eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfd789ec31bdf3457c85e9a66426dc4a873e545741deac377125144b817251a3a79d64524dd2a134398f6f9eebeeb74eb1992135e3e5a0f270d075b5382e24ed95736b2b9ae1e04ad47ed5997665a4084268f7afbdc905ec9eddb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfde9a0cd611c1310c4c23b0c82e9fd43c089211a9b2e9908bdfac55c20917c9254c905ebefce6570feafec489af42cacd708a6296403c37b1d2542381b8d035c6b3e8ae5799cae72f0bd24d13ff6e482bc6e98c61935622ea78064;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad4129226ca1324193fb731aacaf95d349fdd65791464e31f6d4579e299cd57b92ba83b2ba3fccacb91e628d48134583a3f1094f9f7ba21f3aa7421e9d51139690727fb9475d64a32f3883909d32b47ca0b8715b4a5a0f88094871;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1600ef66d16fec939cb723affbece4982741fb7b70e50c3f58e53816bd579ee7b3e306009f196841edeaa343d215855bcf3987f58f578403dad8cf229f8119cb73fbbf4e2b9be527662c554445f70eb51007736eefba16698a69a78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1e009809991248c94c1d44aabb593cc35097c92b8f0064a3ec14b677ff80044b06d8a4f9a91c9ba6d7557e6a99cd1ee4b29ff65376fe69eb886039cc313c6ec26a414216b3829015b152d8af13fcd45d3d16204c07fd2b60281d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136d79d51d07ac390d1fd8638421da89d91c99788969ef798ac074f086e075d68929106b3d451475ebe65723b00e9a97317925aa3811a2eb8eced1397903771a51a955e6c3121682a13fe1402ef5d567c8b7eed9a733ab5ef909aa0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1d6a010637eb43e7698dfe0c75f9833e4398d285f3589586e1decfea53617edccf12e434d83c837708c71aa041f4d5ab435ba5ca4c7e59b0afc40f5a64b204f8f9c5c3f0f06b8d01f1c3250cb59adb9d549a048d41e744061d4f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9ff0a677915b03a471dfc8bda44901077f8f92779306f409294c6906f860eed224159f32528effc726f34214ffbb6b4956d6473802799d9b03b139ee2f5ab569b1ab0342432b40470f7f041b71c8facea2f412b1399b411f632d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1430fbf6c26daa0e9e9928dc2a6475bde4618225d897acc45f112402da24efe29e486c00292b90bd32dc4c407c340e37a2207679d54ecfe4c3028d17fec1bfd3670766041aa631ebf7cf987b6cb85bdff546af75c6181ea3e6c9ba3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6fd0be497d70a8f512926f782cf3c4a64ef1f75a73876faab0b9b0f08010ca0b0400dfe8496bda852e172a18faf9fc71372c5de846abcdcce024fac3f64743e3863a0d96fe04638fd86122577510a8a9f8c4d51d3d15e9975e0d3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a80eb7103a777e2955d786a6c71330f900020c157deeef4b3193c99018624c7a9bc916380ed814c4b3cd8a5fe47c4d5a8244c865c6a27f83ff008096c89e9d92098fb886fd63bc12b79340da691dd4375ee195b8413456b05222a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f5cedb101550c99c989272112d6cabdaf4807285e483cd93f63d95450bc7bb3c3f2a2607b9fa4f0a650c8f498f0b7b9a8932d7f89b9c60099f20ffbf3a7a5be306051e7fca8f220341120993de964a78ec340c8b9b8fccb681461;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3e244c8aa67dbdf35914032ed2c336547825dc26e309c6a9633341f7daf6ea31625987170509390c0356837ef8ef70db18bda5228533e1d26104b0ce014f8b37558dc12dbdce209faf25efcde3b1f48cdd8c4ec6e395704d4b712;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h890f9241938ca29e30c016d32734e76b56163d6923b6ba7ce9aa2f0bb73f001d1555a5892fbfc136b2a4918d5208fe8872278fcdd32cce1e4b5d5a9fa301642dbbf10a48065f2d0e051ddd0f56a11a14959fbc47ed690c8acc9c6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e44f39234599d0cd08a6666c867432a793f1fb82d323b7250a5a8516f641ce72b651aab0d2a1599933021f7318ee6a84675a3334d7ea58e39b30f1eb246be0f3e0da6acad43558c6c5ecec1d287d8fce7fdb87e8aa54170af8ebd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6eaa87f027618c8cb687381b1f3765e3963d19baae665031c4a124692a6cd43c971613bb590ed22e4ca8e6dbbb36b529d328ddaa936a8893ffce3aa1eff237e9dbe98416b36b70016faa185d2f1d135454afc44fd81bfc4991a76e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ce7f5379974ddcfb5cd005cb9aa6b2e960002412d9f2ce3841ab6e0466f3f2c8cf550286d9ef0d630e02f88f5619ce5c3102eb311f7110c3943e12c8682fed86052bf8785a5fd7913dc7f70bfce8a411a864981b76258a4edc941;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6d851909e5a83f2a2c8802bbb22bafb97e45ae12953cf455310eb5c3bd7aef44bbfddc6a1aefd9973dfde759eee8caf53b1b0648dd591161610653643be545677a8225932e988ca055db2ecdbfadcb33cadedb1afc0a63ec997e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a456fd85a992edc43f771b25b825143e4654c218fd87b5f76ae176392cba7bab557f364ace1545151df723432ce91e065d7938926a1b5991088da4a095e32e8d0f58b9a9699b0a028de40bb103ff9c980ba48e4a85e20e434c33c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe724f504013f13243cc28200defc64f389762a5f87b2195eefb22e43d9e5cda709f70692a01a21e1ba4beae6ea3410956144e17faaa1cbc637417ab0b9a97755d6978c4b1890127219ebf7ca3b6e1cbeba6d980b9ae078fc0dfa4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bad871cff65c392b68dd40ce7887977edab47e9a3ea2c45cd0023168f3fd152f9f5793d52290c43031b2cbea73d536bb273ada94876fdf1189636e6842ef97b36d731aab35b248ae1808c11fc447805b200ec3897079cff594839;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0815514a1e7d0ee4ba7ee4735ad1974022044d231d18012d4358f6b49c79dff1b7ce908caeb414f98ff4224a679d44ac8897379fe153f4740d86bc1767f34ecc9bceaf59b99c9e5573de85775664ec11e7b8339ca461680332956;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3db76da321bc009f1f57da02e9b42b27ff3baa95f4e704d839a4c5a165483b4a46e654b54fe2a6c61afb1eebee201dd2b37ca5718f1e92c393ba66c393923773d5f7ebb29434093159b3f3cddca213d593f388221ba01e2ef71a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71697c5580d114c2f7320bf1dc34f18e902d6559957bf7463b342ed2ef7db9408281c23f9beff4c438f38aabe25afdacce7c9f89cdf0f462e0cee7e5c4a71e33c53f505360e981f0a857b9dc01d5761098ebdea45da89240ddfff6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97102ad6aebece272217d2dee5a6263d34bf6e84bc5e6b968f22d4eea82812a5a2eb2ba5c443a5f9e9373d624cb3dc81c71ab780b673e49035bf95dc45c63f764b508654cd6870fbea23cdfcfeba1c4cbcdfe39c211e20c8876fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e324eb727e87c624feeca505288173c120d6cbf132fb4ec88cf1b900a65bc03105e1431e683a1df18fcae4871dc654d550609b95aca55501f57ed494b9212a78e0da0828f0e791e2631f7380dc2db635180673589de3d18419231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1e16413f73a908ec053622de6f71ca1f12000041428a7b7760e6a0a4f71bbb2d5154265f733a2a8d3ce7b0a49af43dd1deff273182efca5cce909b309cd0f16e6e56d65ae09b64a8c903ced10f532c1be03d7af499e0bbd1358e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2d03a5ecd3d3278d2661299ed8959d5e0a017458fb67800630d04353559f3879d0f8f0df927f417e5e52faea66db6e9f22bfd042d60beb4df87c65ac69410e869a8fc5474b475a0b978ffde35ca172820869ac94adbf7d06406ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cea7c1493e519aa625c784be9ab66e8aa253a0e948a6006529707126ad794c77145a86734366283d21a39a3624576f1c49277b598badedd3f0b3dff291a2bfe5da5bb0c7023f8f48e958d522688eac5ff786973f1fa1eda67d95f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38a2470ac9bd231106e7e484168391c0eb2461ebac6d11c52699cfcd304a43f22af57c884a728c4e9f82b53dc3e549d3ae39ba52d40437e887dfa5033e196055242ea11ace8b6dab522c955d6f94063a3b30248bbf3c871a4c1dce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h231b7aaf3205ab1bea7061381370f4163ad960279c49b86206e831d69eed7ee6177fb3805e95e25a3895a73ea4210680397546bf725f1322603fec1cccc0bd40e2ec8353f7c44733d29157dcf42c9f11b450134faa47065ce2e8e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb7ca5031560b8e51e9d3c95b103dbb922c1ddb5f8bc8c148a8e16abd75ece3ab1beb03f7848cca1933ebf14649dacd086dfa60f1e5157f52479d433283d355bb3117d4031ef50919cded97cc08cec5c286061cf0babc325ba05aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd27ba1e4184c93179c47f08d32951e6461d7b07cef9b8f4ba4c2c7eb01b02b6f709e069b70c1d8c42e78bcb38df3c665db845b583dde3985289e6a366bff34907f9291be63fc107caa59947c2b7bb1e698364824a9bde93ca32837;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h388da9e0e95dca2aec740d0bf1313282cd038ea6a1b11a20eb66c6a6f2b7604bfb390e5db44547c9b56ae975360fffddab300e89393e824bded532bc554136e865ad629c65f39a1ddaff66ecede7ccd9ba3aefe91d0c77a013bbb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h341c6094c6ca3b2475bdc48aacb874138627ade5e142a41336c6fc2590b38e47381a177c92182a99f389dd079e3770c95f7ba5f941b2f02bf0597e106181f79670a05c4472c2a1fc53cfa2985f4474209bd6c8ce060b257458887e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc153f5568561964845878217c3851f8bc1001a5c9092646f354d585be511d658d528ccb8da03dcbdc8edce8d84f13d2a02907dcf2b513b417ffad6f5d921f9ebfbab3a53091893c41025adfa8583b3acf93b3f98f55eb658d1fdfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1631f0841018df86ce45376f8271f68b9506fdde601609a084ab8f7b553a9956c5078b995a1e3d622657e5a3dc0fcd9f683f7d107972dbc25305430a9db1a5fef6b674129b66b02e78d4941400d35862accb0c5869049c8223fc35d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142676be99892c98d9c27ffeda0503f5c07d9bd8614337da71d51988490ea6bfca52bff0ae3a8119ad1c73caf92f87ec982a7fbdd4d40d3ede24201b90fc8f8862d671625bd3f39fb3cd2fc126e0dc48976d528ef3f50b6031e5994;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1210acb3694f6f21462da373d4236e41624ff76f6451c8d14aaa11b89242df451d33651879c91d06daa1a14e7f43fab7df8bc42497fdc973bed27310e119a68fb25f3d34c5813720da762469e5eed2ae85943b31da8652590727612;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1480d2e5809113dc67093ad0b8cc80712a40a0a1f7c2b770a467fd6339a6342e020a49fcbb67e2dbe0fb3fcbdecc255e1418bcbbf4ab4b254449d3bb9ea03736cb86eae812da547dbf5ec66e9908df899fb6fb85498365d9a3a3c74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6cc22b45bd0b2b4fc78c9ab1ff3b078fed628c8ea42b47821b0b65943e14e1c7756393b80062a3553382bafa0a800f61f2c07ee1e3a7c44e0e4baa4630755b31c403bfeb9bec3a5323bbd321285a063e7a6a2d01a8d6c90a02b1cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c4617e217746ab59d16f984b8da00b168c4fb7b36d6eaa0e6149b56e20d567a82c5e608836f99d49c981b582b8d898a23952275b6728fd07f989360fe9990a0806852905a1352af2c13d403bd4681e7bd00e65927187e7b1f698a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0b46cc0fc91495ba7f0bb8e6ece6842219d1b202a1398511428d9fa86fd0aaf2ce4baba35d5fe5e2ab0cbcf8f0815b7d6fd0b9deb3501d91f1c19f7d591e131776257db9ace98957d970e21bc80e6b162f788b1e79af38079871;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fac9496e99800f325fc9c68e6e5e59e607625d19d59ff38559e1145dd7cc21629e985badb4a1dc4b596876b9c6f587cc8ea472a7f3e2529eae22279aeac66a121a592326355004f19b6b2713b524c072800a156e5654b204e0506;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196cb3616841af270ef07f1605e591c1138e26ca71705a18e3277f7fdfe0e22f314fd86e2f3bff2b45b099039b19484a613290a5eeb98856c95b03e48fe5ecdc8e8753c2f6ca981abed9745bd94abbe84fba83e920a502153a53ea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h562d95f3a91acb841c8ec6f591381a2861b6dee006e51078250d5bb3bd921719ea9945d44ef6a0a983b0716482bd8b82b8235bf4f810873dc679b4913cbdfe6df37056ddb15e3ddcbc122abbeb618a15cfd0289521711eb4990b85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea7a55f52564a25b2643ce6da5aef741e66d41e9a9031a91b0b5390f3828034d3b98869f6b74caef768cc87834f7cef21b5b2d5c772503ee44bf3494b4394a2cc6c997beff84f890f38e3f7d0f89be080cdfa48b9535aca3838f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b44de1bdd913c1ba46caad3f89d12380e45c4901be2a109c4343f3ed16c4e3fcfb026ca87864649cd515016b1efaa60a7ab9f4d70a23e2b4d397807d5f37f80a8b5dfba8331a17f7e419d57fe13a2071910b081c252bd8a4af112;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89cccb6c573a1f9974754ba0ce3b5a71ec85434a047033d0fb9067030fbcc27dfc544e07ae5c18c1c0d45c37e3513eae85490316398123c151e5d9863fa57fab0c7ae43ef8d0abfbca64ed259190d679a81b5f33d88a2b95c9ae87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he345506c526718e2d69c5585eae28a3aa05ab54e19a3b453a2550b4222936d3be3cf1f5fee081caab9e7e3cfd37a3b50869692db652b2a659c7f3a7fe7d49e0afe9d8cb62a946fd911e0c54417df60df4cd4f96ce7eb96e307672a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd9d6b3f32c7b505bf4fedadaa79f710fee952b3b6108d639266635dd69cf543b4dbdf6974c6bf63429adde5c9a831e5199ce68b93c8957c90bbe56eb0da269f4fc95d695e73acc875e6764442ed3b78b9622fc16a4b392f0a2dc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6f8f56a17d656101f39c10e307e1e24ac1ebb8fe569aca49c2f111488776da4c5c43759b61094ab797bd851bf251af84c7e95902b95f3c1becee0836d2e9274c503b017b7380161672c02e8ab4064821b244ea0150a45d964e762;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2810e470c6b22b47ed06a02cc5de33639a76fc73654331f7b2013fe131e12c25b695b190eb56e9d9cab1770a1a0170f3a614f796955d65487ef3fe488d17e8fa9513458828a072f472ec67a5e7642c757d3572b0dcb9ea5c864c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d731e4a43c4ce3c9869502575fe465978bd7ac76122f9b567e1ec6a7ea9d54dfcdaf92a4c0eeef0ac3cc8586d5153f70dc0ddaba55d43d65e26f3ecd07d1d3ce6e4834ad5565522c17540d3eff6bf4b29b033c308970a7e4c7379;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fba86e185ae4e4ce2761a3ce9161003b0908b582477a85834217990cebf49681a0f44daa1b90ff1e3b55ac1d60dbe9eac5c021d1fde9ea2813eb51b512aac720f18c5b02028e26bb2a044507414ad38708e0a860509c58eb7a2e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ce9bba8001b934d381150629e96ae3bbd44d05f2dc7847fc5c73d2017e99e9caff3954b00837975862f225b50925aebc8e99327d9179866d7379af8bfa019e5bc3372613c57551ee6c91c2e6ec08c682122e77f4b457696b10a29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e45d9fe9d0444678c315d3d77c8ff9e64d6bc031d91c263662c1c7b98fd56ea54ee6cc54175495faadfd6f63b3c66e103c9478bfb20e6c852a3f8087ae07cd773f1e33cbda7db0a739e86e2cc85d8838b5562bf1e8e76cddb6fde7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77044e296d79b6d5159b40445cafd41d1b418b4254bc2080a94e9f2ed8117dddf5ab3bf29d05cab9d9ae8fbf1f41f3c057fb4c313b2f68515183c17cb2fa18b2831593742a51f78b89a81743eb1778991b63ce4ed5e1fb9cd4a492;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1ddb68ca2e6a9c8d66773df31c5385dc80f1264f75ad1100be2360a03f6a5b4d7821aa179d9c6ce61408ea3d77003a1c590e7372df63f892932c8b106ee2c2d7905f32fa76e84197dbfd4fba08891e866848d480a1f1bbab54610;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b614d5da3d58cf54fbc66d444c0cae29f33d861f859c43de4e7a7a665c44a855a2873adf4cd979d4148e4119773dc1689dec48af288409ead929c73198697b793a287f104c1a7ae3fe2948bc64645e1d7a94866a26b417e48aefb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd021559fb7852b046a8358eb511e751311340bd65d670f780498cfeca53d11453f5a657ddc4b9aeb96a8ac748e44aa648d47f352c7980dffd8419ab05e92ab91f3515854fa64368917109375efa328cacbdfb339cff490b9df8dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d89a5da6652db0744aed32579f6401fd56d3ef01f8e11c6003611f18d9b459ca5a0b91124c86ca5f6eaafa0cf58d1f38cd60e1b789ca70c77b4845b2163f0c98019ee5d4b4e0ba9cb42776f371896aa310fc4ff28111896d3df7d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0fcb583ca1adbeba1069b36d5f52e80028d3054514b5b863c59652bd2f95e8916e249022a63ac020d2b4e85dd8a096304f19bfcfe85e639d7daa0b49de25d829e5f74e389aa213009445cd05cc4fa371d788529fff7d94462554;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf32a6b76007f84cc303391a4aba4126096024a66da818da65151ca694ac181655193e9b8b7e9d3ff12aaf318907c73e420cccc13cbae219f8668ad1b1e51918448e547fe4b197e9ecf30e580b6d3ef1e0a6b2fc61606e0d52d7b21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2828a084d1fe5ea95afc51c79a1c22c759ab0926f4c4c5e24bc98fb3f328025fe9071468537711f81f1852f0918eb3609823d4164ef49443ddb766a82f63311108c34d126fec3310f631b3eb2935b337cdd8667fcb035c05354ce0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fb0b098ff515f72c84aad8422fc8348f8728991d47dffb4aca86265460161361fc8e4445555ca158568c1a9ca5e7c04467b910a8a21ab3f08555a9c203d131543df7605e4cb71cf2f970dec15a177cb91b1a91deea80b3461a281;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69662388a0bc33d68e520f019f27806386c51a0c1419175f0ad28f7593d0f5445c0680f586d8e8db75f95456c611c8b0ea45c69ecc0dca9c940bebda4b5c93c25b1c838cbf0ed23b4b2a4d7406e1bfb215f232732db08ab633bfda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf73d5d3e8e56beb2e607fbf2a4795ceb793e085d93eb36af3949334a9fa667b3a845b8a443ac05b901cded89173ab1d09a8b6d8c460ea567bae8f3f8202a6d3b1040a8a0566e6312a017c4f15809febead94ea184fb0237d442fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1484d5a7cc0b71840b242d42cab7adc865464254364d9e463024f7d30aab3ff10659b37ff8f7c3f76978afe919ffae0e49e6879526754afe56bf3dab80df3a8ef01f03917c8bdd8d1b8a5197ac10e81b0f753217b26b197ae40fb8f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eeb0f80993cf653a3fae274e1d241caf715e0053469da783742cbd917debcdeda0de9837090db836510a478b2ebcb5fefd3ad714e1b0e435d4ae437faf5f1f026a9fd5a16abca40c722c63310dc64537e5a18ee7c682da12f5dc99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8876ac1129d3e86dad1027604e9bf1bc2b522f78ac840fcc250f34c21eca39a4413cbf2ab4438958f37f8ddaa270e34f7f8e73213869bfb0c8bbc1e69bac5499d645743de8f0df30dcb1281a9828a55ad53212e00c0cee23c21af8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7069656c33e0efc80b007234e65d49cdb56a6b3db2b32e05d85a9a1c3fe7df6bfeded07d51c5c5ee544d047966d35a52674f1f8faa81e9e32a0a67fc88c9218d254428e2fc56b870523209423cace302294c522966de0a0ea57057;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78852b243f48fe90a17538b374f99d7d54ee1d4d88696b310ef4077dd32779a5633a3fe08d923d048188143400c28443bcaea51d99f7752451fd34bed7a83e3e9028ae5f91d86b0ff97e7219df178cdf0bc765dccc18a460c969a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e6d606d8190a2caf151e3ce7a912e491dbedefca8fcedfbbc11cba92033d2f844621d6d03732d16152284275d63dbdfed5470044f59d4123362dcca17c3b8364e4cce6d0c36260d1287494e85dcd761e4c9c3efcbb1d1b6a67c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af02802116b50d2e53db1a3780da548772bf0d2b4117dfb08611a6147ce9f8901328f660bbfebcb575073f7cba76c5ca1db1c8553dcbfccdc6fb30ad340506154cb6e1f6c88827fef4dc74cdc3efd8d2e9bcc27d01f18b8342f571;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130afea5fdfd79e9357d8bfb80e70c619e70894f6b8d615422f3b632931020517367c701c3df4a3f081903e295e5df837ffbcd633582ce3f936687d0078b2b9dfa9b7bf672d3963f443c2678a84bf7402392ce431f9007cbafebeaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ca9a0c3d533af08a56e16b198987ec33167eb32ccad6d6182643d1e36fd03e7d400d9e38ea1c9e0b40725090f9af1457b1ef9fe8d5c3e5c2954c1c74e85772f6017a306373297b54c166dbf31ee2d58888750e9e0e12902725604;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b4e0ce94057f0413c6caf59de085a42b3dacce46d248c4264781d7b9e0cbdfa426ce14f1f4dc93c9b154f92b149efe83f2ef12b5b9d0726ec9071562d04d8fe01905390b68cf78f7284592ce215eefcff40960b30be347006ebe2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154b8b942156efbf24aff5664f1fc350c4be34b69a4a795666c803d4c75c209684b53c9f289588fdc1c225eaca9b6832f7fd45a7324910025c7dd818b9ef079519cec0532de87c932ff1dbabf05c21a7ed137c82148e19e68ffa2c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf57b1feeeab5130b0c6d33e1cacb850d3b4203620c59773b387d09a5e41dc2e36a349974e8067fa1c6503541d54faadaf55bded2b8ad3a7e84e68298a53c088d017a933ad9aa946b1f78497449c1d53c460c2da21d1642b5643da6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1271db6846a9c0d2d7bc89260edad541ac03e7467c0df69a51d001ca49a932021dd757d28b3957667ad499fe95de99f0d9af6cd2c29b668ce31df8421af4976ff48c21dd3c7ea170c36ab73f85de6543ccf5badb49a033660f14fd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h969c6b558a5d81e6da1401e3f3ca714428b1d6f69ec15a2ab3236cac80b361133adc3942467fed290d7ab402d35e72ca976bf152dcc00d20e3c843cd26fe6e71dd16b17bffc9a3c0e007bb984e09783cf198acc91b57c061c75a16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h503f9fc85f5fff49bbd4f55c4bf2c2f10c6e41a8295bbad27d81ed59d6de5fc6b7a7e28625512b6c68e3a5ae333dbfc369950e91a4c2f4dc2df194e90fab3eea2586727d9eac7970ab98633bbf7baca2065bb379f2affa2889703;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1100bfa2a08dbae5369f9c8d1f789792d90dedffd79a61d9a90e396f2d23fb42967dd2138d9cd73d19792e0002745b691571698b840eca243d1c6797608ba8729f9ece6f1e70ca199c4783c9b86161986f3f9183dc084395ab753cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb02f7dd992eff438348d598a5939185ba3369011ad46186cd404503f56f17e686f65761552205970fe95fd494bd78e014d080ac713051646497c1071382967834e3924b398263025337a597ee139b5d21dc23de2e66bbfd6f9fa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19894fd6e7b7141bd2cb854c5e03b6afd5ec2351a4da94ccfa0e171f67721fd87ed45ce2a13ac6c2fefade49a28f73e0ade1e1660ef19649ba4477461109eaf0a3661222f1b22ffd4f2e4d8021a48b349103c4c8ea4e565075d160c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b223570c5e8ba6cbfffa67cc3369049b5d0c4b8bf6c2bf60c75f7c62693d5fe664ed54a8b821e5960eb374365fefe5290faf1bac579a3252962d5a569bacd2329289dac17f8637e7c0a843190344e70593c935bb4fbeb658ac21e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5f5f42450a6edbf65822394fc1f72a3e0987088872887d087c3c1137bbe6635c26b49adc27caaf000a4932b31e55b48a2c79091742a421d361186c48ba89820c34d85205f0b0b8136364a6a82fb04a4695c63735b7485fb1d4359;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h505c551fa6480d499e1a61545331abad863a462462f9a7a25280e8e55b972329ae265ce2823bf3e4af589d28d997af38622471af42a475b6f63e624eda419629e70f0026c8309d73c54c603e778b79ec3c28e6c27ddf3dbebf1f33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d6ac21dfda6c09f3f8ddd21e00d6c8181baa584b4cef14d3be971a7849a9c64c81d489569a41ed15b86b439eaa9a22774794d16723a051a0b66ceec563f8bc801da9d1de711800a770d48560ea683642505840cc6096f81cb7b93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc09f55ff0dafa0882e5b216eba82f1aa5780dd9b3229eeb21f6d2ad8e1907f0de7f9d5dca3dfc4cf82321076b572e0f80f4f524a96bcec197c6dd8296aa6e6c6ae9bca311f2712f0c7cc9f299f1dc855da24cb5eb6872909ebcf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef39e2c4061601274ec695d5c9ddac1dbdc0b599644877c404e8e4de102ea79aff013b891a2f89a6dc88372f8944116ae25933f84003d3fa50fc63b731f7ac948d6eb23a49e7fa14b205415b7908000a1fc16d508ec204a6b50ae1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57c9ca18080afd23536f9c4657b0b536945795e4ea051f711e1aa865bb25278de7993c9736c5691fc32f462092a88017b4beac1fa82be02f8ca002c1d86056c8b51d26243c2bca070ac4281e3d367fa7fc53d265d0aadc392a64ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1355e9535f3077653e1a31a9f4dab11639e1727b0c5c244322da0b966d318436053ad8f5f228f006c4e0064b412596a6975d0752d234b531259eb8dabde077306437a55236fefc099ef7c1a57cd538892284efc527db7650b75dfb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5429535d8c724b3c2ddad28f23ebbc30565c2334295ae5cc6308de87fee74e88f735b88e8b6defda642d5c5af75bd6da668b02ea5f96e4fd87970dd78eeb0ef23ec1de3542c30c594c5feb9c0d74eb7521fc012377bf0eef46c56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2bd625c39301f8c55c8d348dce7ae62a0001a5fc3dead7ef630428f3a919bfda2ac36e11f998b9f3fabfe274f6118d509ca3d6aaf36412d65d8b1e326da04fa2a47c8886ac248d7e059ac3f522b8e414708e9a46ec8213ef3a7a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19142c92b80441896ac2269750b0c8b55b6532d3740e6c9353d47e64d47babb7fe42b95858d37216c6e285bd86ac42f6c8da37654b5e10b93248b28bbed58838ed59dbea62e655cc7b4a285805e84078011583a0922c3643940d70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b75c9c2de79125729109b1acf3344860f0d297da4c4dd55573421b37ab8c0f34ea56d2b70fc78606c0d94d09a3a0ddceda43ab94bceca72f18de6b1a535da61b7197bd70d11711a03e0f758923a6b7e455e7befc418d3f53e2aa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baa54de1def7f3dfa05defbe63b0bcb301c856445d5ea7974166c7ca040feb557e8f367a68fe7ce7da5405184bd9c4924e54e28b758944f170235710e8d8ebcc55fa88ce49c7cbd46f957ad8e9bf166f6ddf4cdb3c2c787d442019;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha25cc31a82ffe76a0af94a410881b099190fd7b4912859041eb81aec3108b60462b5f426a225119fa286462c1da04b2917f8bccc8a9c89153126e9c44427b018ce54c9b019cffa127091f09962fc1a6fdccebdf7c2c5b4b01358f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191bbc81aacc6c4b7ee0d183d09ee002c03ca84af5c56a31ddbbc2d1630d694aae2d5d3d0634399233d94cddb53a53ed48d73a232a6b1368b406c322529731de415e2d7096c7fc39522e81dd2367f1e2290331478fa97080b03374f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4bb1563816614b6a15c72e13e0c62d33753cbb0500dc617be16771f98361bfbc7264ba1a354c9a51e2ea068f15ac87cc5f277878e61215ff01b85506626ed3fd35e1d84d3c775bdc3c0b93787f10bb03ac171d2fa4ab4f1b867d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1474a31126245f1bec4693149bdd246aa7fa83c5cabe8fabde47f929a6fdc42ec057c79bce1354838824369d711ec759e58e578b7134d77afa31dc24b56ec204807a554afb1cf34e6c32f054cbf1bedcbd8b345117935e323e71824;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2dff9c77fff9db2c595ffd50fdb26621e47e2f76d6d9dc8435ab4dde56209c00ada75ad70ba22a9d9e966c168c9d630c23ddc98055677ca3cd91032cfdfd7d1c9ebfefdc6d9d7e388e3fb8ba112cc43c8308a2423cb1170b9d7d34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbfd77fa145d6a7acc9013b03d2214ba2614d2acf5f4110983451f3ef16ce2b4c9b112dac4a23ea522e49dd7042c66bd5f73628ce4fe718f6c2d98c9f1e235d8172f37a12ac53e0d48bbccdac760f59a7296bf74e61d04c931f235b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c03b846afec25373977dc2140a56ce22c71b0a79a1d8384eff4fc11b44756408cb248520d528ee0f745cd24e8a0321799c9abe7deebc2825260722d45250f96befa2b4b48f9b86b116328ac8be91c7802470e9dff7eb4b046ca6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7687a2c60329643b565e2f507bdfe21dfba9557dc99f1fb289d37b993d05a21e25c7aa6ad72ec1910609f41c5844203f3fd24851c034587c717bafc2059fb2e812a86c5d5f02ae8bc84a49627759db3b841d102ef4e94ad55c2314;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a4acac3873ef4225f6dae3087f9aead39562eb3a6d07ed5b61b5644dcec49df5714a68b65fbe5303bfd60a929ded6b805650249b8fbe810d6c4d4f23e7acc610858d929c4e8393abad8e4c5375e5444522f390ba084eaa3f55f39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19796e60b7f8a5e8e5a0019a087de6726014356c68e14951371ecc239d582f5342d5bfb3080ae178aed83d16580090afa6e4d9a1f2d9eb10e6c63f2e74e4633efd4151ff840ff76e92fc84bf4f295313f2d6910e6f984b73fd677d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6ab9c669c63c43f339e507f0d22106b5a37036e27dfe5d7a4ae960f91f874e8f736ab5a1458c9f1fd35c560cc24de8a95eb4bf525de51efecbc9d32a200977f7be2181baa471d589d4f4540b9cea965ae11fe6bbceec035f11f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae3d0117534b092ca13d1fec46c6f78471a24c0de6ab9e100e84cae849005b72ee7b00d14aa337c7db1f6154875fe9d01db3808a979f6b3fe4185b518d1e550940aee870cd6dca54fef222e82a2770bed562a3e8c54d1522b84f15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdc9384e111ab6737a2a44df11fc8b8cc0b3c35c89544399c486092dc0064a67a9b7b8aa29fde6b349cb21a6adf2ff28a53c6eb6a112834594ec636b753d42a58a47cd4875d73b6e45d8e05e235eb56c2d6acaed50e30f561f7599;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b73556c61a4e5d91035b43580651ae601ed53b6637782098db857dd7380d045570595e6c59e8b17f19f6daa00267ede30e88e33f5d2a5ebe9dfb51fa79d79b9c431d766d9d384932ee9e8a39db72a7322184daaed51025ae0757f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15885736c30d6034b9923ea312f84a4e045b5b3ffefb0d9351029a231658a36ddc5a686b2b19e29a304114ce4aaf5ff4ebeacab37eb381569ce8415623c17253ee0ee3c9bbdd3016f5892a4307a65d899d1017e45a22ae4ffb084c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb049d653a19de8eaf56edf0ea56b527b01ad531c5dab5030c7bb72a0c47af661843053b46156829befa2f241c6c22766d03a7b722f4a50ed24b6a2ce9fb4c5e246e8b5a3c3718ed497be5bc64519d3739943cb524a24fc87370dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha33cf251e8fa0fa6f40337ca43dfbf36cc9290c5650ff2b2b5d6c8422e74db5aa2b8753f9e73f19c10e8aab8f86c09c7267b4efaf46487d6283e1520c27b7adbc4ed649429191813db4ac0cd90a64684e5ed01020812df1ec598b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1840acd6d72688cdee0491c6f0f4cd590747e1cc3b1da30bf96b823e7777c36d2a038567b84d104cb16ddbe562abdd338d43a9a24c5f19ad52142153473c13bbcaea2201744547f26904a64a6ca36c3051083110d4081287296de41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170a240ca93cede41506c081602fb4320394624911a4ebb12f4a8b1150273daa73a19ecb5a5380a0cd5cd64885e97c96cf1fe0e86cb7fa5094cc9a3cf401e5a9c0b8d9d4f6b6324ec9fbe1ce5e39f7eaf282826b1fac43c4d4996a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ace1771339b71492ec41cdde1ac87802155907d2582f864785eff00ddecfecf992de9944e32e21bbcb596be675ba4c53fb74d9d64b9fc5f4d51e3b9a4e7b7ecb01502db991e817a750437abe003a4fc99394b06d2868b37b5b4d16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140dc7326c95627d428a60ee8aea3b19fd864ef2949dd9ba6b9f45b42c934ec881d66bd5c14e43c8da4bf2efb107f11a70da3a498f7e3ff573a14fe530d16d318e1b6146dbbe10f4337347d238d212b16bf6d7af9c778c8c8004c74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b8eff4f81c8b65a8abd11a332df241addee549c0de710b9689faff13457f14724d10cc2a3fa2cd1ec73d21b68dfa64b282509407a28e554ad65e9260a3a6e9e1cb1e9ea6b768258043d6de2c8d7e99cac5f14f4398453eed28302;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20db3758275de914aaa6f52dd9a367d79c3c56ca8916b299e376a953b70d8ddfce24c542627a6a7e0cb89978e71ae1859b484fa48aa84b7715f3f5411cb8d189072f30ea44efb61e497fe6072f51f5b436de4d04ca396433222c98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8d814c84659762859f241fc4d0401ef5cd71e56a180b645e8ff63d39334455ce86040ae108dc5b0e0ceef5b7eeb24a5f3c8501da83feb7952e592b3017b1211f4885eb6d74d2c4337df5d9be9e3e04e32716f67ecf3fe513fc2e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd14922cd524acea6d1e328b6309875edd07957b82ccfa52b17ebcdf0f8666b0d62b93b6a96c6b318a8123c34263a99248529efb4a469c67fc92d50f6f47424de74929ecf3b8ad2752cc6071a4d1d5959b9eff934a35b92f3d66180;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h687575f0cbf9904876cce4dc4d465b9c5b7daf7775128730b01b089c00828a40b3a42ae06c806a9be44c241bada7367bfc6c8d1638d8008a38c296d338b082e589d0d9f1b4ef8806c9a03cada1cfa97de9976a92609b4a1f3fe7d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b733f3ba221a67269ace8c94cec2101dc7dc9f3193a79dc6a32ffd2c7318770881e04089d22038c720a3e4b43572e43ca0c72ae5a6e48c10d40966e1c65b104393f7541425aebe2b0aa122c28fa80801574ca54e67e7837e4920b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c404d24c312f27e1227ce72d5023c2a84200926700a0178b1b4307bf1ded2aa356f23d8eba79373d039e0bdc29263ff46914b5b5715595d60cabc1def4fe3405ef0d1dd782c82070c9630811defc18c1e36f3a79e7d935d607e5ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8ab727f14f577fe7cc723150b1835f99825a129e536e0f5ab1d1cd2c8cedde3a06f2502cbbac2026f5f97e5623224ae3217c46a566d00b6edcd3dac9e4777aa37fa26de0b161a03c5539cec0228bba1b5572c80954123dae9ef47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4b859c5f62dd9245da67a95eea943c13f9f5ad8d2e84b7d04b33454db173d3eea94f39fd1c5368a6cd3f0a2cc7e544ffc20f8fdce61c8468bc4d3de369961579a87fcfbfac7297445a0dfe5725c58cb97ddfc61432410f9b7df2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb774c56ead0b62a7b7236439ca95ed2e4e211b7baaef6f2d6241eff5158c07a3182ce15b1b618e32946ff14f8b53710566a28fbca15f6f26088e1a0037332813c75dd69a5c603ea11a0d29449270eaf9e960a44fc0c9ceb3f6170c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3e23b8ff39ffb2d2d40dc3bec1117c500c6c7eddb4282e6c614b8319b61b6ae32a527d3438c3b91040e212e7788f9141efae4d9285f77bc18b3762ace60d13c93b33a4230a5d6171d3e973a7ae8fc2b6e7591c4221d77c2b3035a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a13c90ac51a0997985afd479f5b8e6ea8745915db56b53f5137eaf2e7c86326e5175a6713d9a0069fb5970d72a86b686fe876594164f57e1ce409ff7b5a4581ec79e25e1aabdbfe07436ec5cc72f8109f0709cf23bb9f489459db6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e36decb2e25ed8836d81860673d2acd2dcf84eefc72f7d6d0a3f9afec7e94dca881855c8c53810d2b2ec92cddd68e0616ee874447b4791a337d8d8329f5e778ad7e6c893a806061df83565338a356ba0afdd32395eb0fe25146f99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f63862f1fcdedf0862c2b593d7f4573d32350d6bc9ba907b8072b5594ac9d74fbc91abd42824c2833c9181077356acd762d2001844eca2240d50c85f9989a21fc8e998597020fe7b8f636c321475c0d82ab3003a583ba2706cc896;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ab15d70aa7281eb3c59e752a6bf918b3ff74f51475705a70b5192748e0a359bb78050812f6e6e19b62c5423523a9827488df6354fd82b9932798ea2435421b4030fae0f79f1af4dd2736196772a493b49755a397f632cea1f6a26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123ffc1e77063994d3c87a81d1f4e247115682ce931d554e2d332ae5ee50a4d07bdcab5067443f5f59e48983f32ce13d0be196c2469d47911983b37edf2e8fe1ccb376dcd701d77b6f2a57f2831b33d89aefb79d1554397ed746361;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8c6b1741c3b3ae71067d1c2adf4790815eda93bedc1f5a1a8b7497fef472eb02846b5c8243c848b05cca458b60fb79120d4b493ca471e94395bda86ec01d9481498402193b06492ee7eb9a9bec2e5e77979731c7cce6d3c6faead;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h895a83ed242e544f32e0b88b18f44d59de3200b691f28e954e81da33ba875d4883971fecf3e4ed71b695ba9b325cff8d63ed42fd0325fe5919e61a256c6aec6666d7b8593903e3dba94d35e9196041620a30b8ff4c3ec253376fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha906933f89ef4fa32edc2e28f8bf0ab126804232c203dfa352b4f7c7680516b23b13987a321e39266807693d807227408135ea42941e2b7bf8f83aa2fd754854d2a81161f7d88f7105d7cb05fb285f0121ac4aac7274a48a317587;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h829861cd94688c3df6618b733ac3873266ca002721fc787b17136ce57c81b35114a6c0e7b55095163891ec74137773819f127ff5ce311bdae544a59a423313f7c5ab0babca692bf311945c88dbc71fa2dec450283aa9b30e9d1247;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18643911d5f19d2256493ddc360482897a810e7d671b9919675dafb1eea18f51935743af2d89d0dda08e22c3ffa82de33f042dfab9be82a9bccb92a70a7abd0bc3d8992ac85cb724f28502edb5a8184a89e7db997a1d3f977540fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ab247c9b8fad03d4c24eb218f3a90ee9e2e14ca1140b00bb211968925479d762e4fc7a90ecf6d8b9c731cece8addcd55c87d07e42393841a62beee82c9a9de3235dd7f622083c85e1bf1bc49346a78047df70dbcac50d959845e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4070310f1a270064b5327e9ef2465048d8664a96d39376bbe18557d072ac55b523fec4744976f65dc1be4b464abea901561514198c4330bc8acc1b712d7e4be2787b9cd7d759b444313b6e04563768285f7da68d4e68b7cbe2b9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d9c4047c79a069a113f3b3a6c7ae87dea81ef5578fff05589a5c79561123664b4970fa71365f7699c87288225fb2eb8fdbe865fa7d5771e2d6aa59049913e8d8c78823c1bf4c7ce02556a03293c16064eae489bccbcb8a43567e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68e2e81618ae34a89fdbca4a0ea5c2b37b2c0d5a738dd0351a7026d4eef2a68cacc3a59b2ff2f930ce48e9790c219306570eeee5a6fb14635fa137ba86ead5b0c8eb133c68c42c6a87e1913ce50b9974a7e1739cb88f194d9b307c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdf06d120ac96dba469cc997b2282fdf2c7180495ad3b087e478a1b0504edd33619046d1a5b1473365659838fcbb88e00cd89438da930582a72bbc5e30d4de6d1293df9bff28b6e2f612d110bb947c2f94255fdb50a7427ad74e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25d6bdb941e257bcf1aba9c90b5b5684ac2df694636b26a640a186410a94bc94dc14b9d75f6a9f724df68a33d9bb3176f66f992ae2e721d694d1f46b6f319346a58abdb7f6a911f3d26efb9d3a631a4e29c3bc72d2a4f34b28ab35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h877bb4f94f1923a3d3b62327f38bfab51b14b6075748589c9ae1f093e1593c2058e69ae21ce99e2b338e76f2a76f769b7db8a6f882bc3cd9286bf1a7266e707674b1905c91ddc5c9dcf49b0dd23b6aa24d56cb538090432bcb25d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47f53792af4789dc9c2bac71b1d15169c4db8cc9352d972c177a0d108e1aa125d7740aa9eeff954b76ef809dc0d67eb63d0009d1032c9d1cc4b7a854e577958db53e2a87f33c2a0f96dbaecc7a693be3acb127dc42b0f892b7867;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5c161c3e903d40c934ec2e7cb4f4e2208dd9c1305ec41df6a53bfae22eb33534178ace5abd4093dd065ab461289f42887e7d0f01cd8cd0ba4f9899ec5c5167485cefd0342d0e0a75a2f9c74c941992cad16bdeb4b8b000ab7baf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c2eb492be14c4223e63b7b7059e77333cb910a0c64d8270d9f0db7e8284414f5c58bf7705d3d4b43fd680faa20f11ca7d88d00503e2a31787fe9956cc624c1226376b9ebd3b8bb33584d627c573de8095b58146cbd9fae56d1788;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0768963b004632dcb0878db28bcf87d447f3bbea067a06e114079eff13fd643ce208a3fe49db7485e5b906f5e7e4c3339340d14176188729f68d895d3db7dba2716c7b15bb59e7c3f67c68e7becc2b00f8fbd3a86d99757bebaac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b72eac06fefc53320c570b9c440368a13cafec4ddb9c113521744007c657cc209b08ba18f8372b28536baac8b146318ba0c41aaed3246db0bf35b81a825f2bfa2322c12f9d4631d2afff0d1bf06241a792342ba6a4de7e97fa220b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha66764c21832f6ca01ec2e9644952564411de646d646958310fe4f5688764b03c13a79906435c0db971850c816a022103021954f3cc2c27dda3110f0c17547075ae5608ca642df7fab4323650cf74000e93c3f638dd3363f8b91ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f90ae03f64a98b5f46ea462f4b0634f28645c1fa09290aad44b532ec9463e21ae2db4a418529361267e07aa8e881dd53c8d81fcfaf77b5c3df4d3920e245e2e107471fc419cb72a28a19abdef751667a846b192d12a0a2ac7b07e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eaea36b17b7b13d25428409e46413db28bbd425b992c26f6522297a947a0a7d4daac592eacd0ce7dd6cfb76b52a391505ac5e8a60972e815aa7d90ab50962f4b0c10d7eb3c0001fc1da5b36fbecc33e09c6988e46edc497e8ab4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101817269d793b795ba2b585087bab01a24f9ec87f9b775431dc2531eeed7352baed07cd87ad551be5c0b77116a7926618f4625f60ed3441ff7fff462dc7769ce7e4e566e59932fcca63b9b24a59f5c8a1e5f84302ad7885bfc7403;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfc03956159f6f1f07e08bc54fbf1ddd08f27b188950d4f1d3815187a3014ae89a3caac385e59ee375540d50ad53679fa5d78777e311235ca8b48f7512b7d047422d4ca02a889eea89b208b6745e2572d81d47b2d875a78301850f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13de1818da5b075fc93f08e00232ab75c8e236ddae61ac31b9ff568a95bfce7e5898d67a4677406975849073ad81345dd912d2b697a7c961c2416ab2bae67f48111bfbc69e7ab81a8f614dbfdd1e23df42a6af01fc93c2639a0fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55fbeee8f9ca298509da6dfe03706c1198b5efae7406f4e4cc0d09f82adc65425d515a49a0a70b16e248659320977679c67e11df696655745284e3ed7b36dcba569b49a090ac1265fb6fed8679bcf343a7a412d6e5d48fea284cb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f807ebed4d66229692da6b85600a848ebea9cba7fe550005a3b25e1717b63e094ad17def5d73631e316b048b96a91c6b1742166d719e8e059c7e521686fe605065dd7f90b625cda9d4286464145e0129478c47d66c29c0db56059;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ee8f4c17207f33409ae47d347e7ebedfa519b89a86c1c04bc7c311af16702e481ad02c1e6cbd6e27b40e603bc19aae54e333b671bf35c814e4db63217de84fd85bf0a722a5c8524effb0d9d56ffee0ab949b6acd2441c3bd7ecb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc244a6b2bd403975f7609efe3b839dcb85e308f0da6b8eaf20c359641c6b0240778f466395fc2cdd15d6a3d4caee8adb002ff4df0a74180d948511f8388734765fb97fabb45373c4ed162262d0b7a23ef556eb3161d09e65f115e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184a85efd56807b2b4733d3fdd8b94db6e8138347b4a1856788852f1fbd220a37d8e2af26cf179dcdd06f9abc72b0573363c3be4ac8becf432610c6cfd4e68b393f50d1faa88b6a6cb64927e0d7a7510ea4405601508cf93e2c7a0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10dff769db3e91d96e78b3b591602a31d123bc7c982d21c7fc53531697273c2a95a6528b92e5d940396c08dedb58ca195d07a5b7b3b83ebaca6deb958c29413eb9cfa1c50f801593219d13ec4fe634066b2fc21371d912f09736f0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35e217b933f4cbdcc83d5f3072a2296b68d4a3c87c75d384a1b6fe85b7ee6bf63700f2fdf970df4f43893b53664669ee37614e8c8d0d80570e10d297fba7b995e19e36b1efc29018e0d6cd884ff71f89bfe6a62777d562fb9d0506;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7871967a25aa35cee6d02ce2755a08d702d51d64925e9a75062c8aebdb8702dd90beff96f246c7bbf8d5db56820acf1c8c029b80bbfae414325ef2917b3723e1ca088a882f988d5ef05b036aa34c35b7dec66ca64ca95007ece21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb9b7c7e256d05aa8765cb5d5ac73efe603c896c6b3554faf027a13f35e25b29f8b030ddc39f28d5faf60643b64dc33ff0acf99844942723bf4b1f7e41e3b2e4688fafe593caa1135503c76e8e82d60c942e4c39d49c15a4daa7f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h908a64fd2ffc812022442b60c3d5043945d6ebb2fc766b0c3bbf020b0685e6a7683781f94620940631e110b6f618684e3f960d46f69a194287d58cce1781469f6f435875dffdf2c496d06f00d22c2279eb2f2f0fd3c2bce909cd5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182afe557ec5895ebad79c883384594a03f0133bb6bcae892252dc7d518fc1a4b50923314ec78b0b0fc9ea445e68b8a0a2129e08d70d52d763fa9d8d4fb16c018ff6500c711c35ba6097bcdd361397008e35e24f842d86166e0b5c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f1ff33a837e56e5e6d373b8aa46d56b21b08a9a1c17b1c82090f28ee90848757803e488c474827db65e340db1b3d2fc98f6e97794f40c856dd2df0ee51662954c07d4c9905835a89f241faadf2dbf03e9b58c15b82016e5e660bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12be8ee344d332aa4f4d8543eeaac8a398a6517d4188955c2db8903d2112dc9329a261866a8908399a14309ddd651944e5a21fbdee595f7e95d6ddb2f240ff0a714257d95aae1f6ee8bead9ecf81a5b4b9d5e4ac9c6b9c36018993f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c68ce09828864f5f575b847eab0237cab8633e2357a899253cee9662b028a4c30ca2ab68b8f8ce3be9d42ddc1db1125406aed8cc5e18efdbe2125ffd566957e26cb497c70b0f977c9c1903ce73c1fee5e3d7646acbc8ed9dce5b1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61591788da766801471d15060e3ee060b6deb28fae71cac861945f4986702977c69a71b4be7a4ecb879d01c145062488f82a2cdc622c3b7ec29435ab6117869d43d4b3516fe27b80058d474ecb2412024f6b0c7b57f8901c0af1d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha572f8d374be42d083532bb824cc290810e402b39d557fef7a5cb7820877f0036a9ec3b888d0a40ac3a007962c8ca5374d784255957ce60bc0d01ac6b9967e2826090b06f5632ab1355c869a03b704b73bbab3e9e96a2972fca11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc25379e8b6b0f5bf7c0490a2f593ddaa2d1921d39c9363660ed2d365f61cf3d67099f7ea6c81fbc13036a43acc9225a633085eaeb84909a28c6696ed878020cca7c539881724e6453ae14cc4803f020408a26517ea6827be63e9d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3e2aef94697b370050e0a650d1b20afc6a5d86f92f0868f3ffcfb9ad3abad62f27a1b88e79589bc16c34a8f67dd8f13351a5fe3aa46cb90d2dca321e13707799d7d104181c493090b68645a6ab47cf2b67c72f9136df9d0f1fc82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb20189b82864af5813a9d5c351918646b4d6ac15528dc5466da264a093878f3f7729510879e17ce35a4fb9469c2f770b398bcb87f47110da9e269bfdf2ebbd6df3c488beff0d5affdc60365a5c3abe8bb15ef81c322ca60348864e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f01ef7a00809c8a91948c601e4525142f5ed1d4e2908373f35e98252d517de95a2f86303a60141582e29c64de000263b305e155b0e479bf2676ef306bd7e2a44d71866cc9bded05506e213df841e0e75bba134e1fc452e699f0b78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e4d464187267716226467024111a60c483c6e0df86d705acacaaeab7803d1a0c5afa5f27e9f808ef0291c5775d885c03ad4ee5e8348a379dea42585d5c6d2b498967664c3ec7ae52ef631d92f2637641cffdef73ab227e75a5183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb9931a1ed4bd01c6d0892bce72e01650f13d2b27508d6d5dff38e2f2343be8f2340194d678a51be42fb8c6489c22e8556ffe27f8d573048511ec534ff5f802f7ad68ae30ed42eca03b674e93b44122c8c6b69bd456ba177041cae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h947600c389bf1e491c926e3ab866b3be14ba0a91e8ae55ac31312bb2aaa30604b1f6e007d40a3b4b3e010cb0d7852ad7b37e65dd5aa59af220cd4fa31d1c9c51397ba31c0b40ec33544cec5623eb8d99a5e04fa5d1a5b58d1de1cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22066204e2619b6573f09923b33c5104c4a35ac09b55deda93b96dd9da6a23a5d500f8a24330c727264561b4fede86f245c11495efaeed9a2e47e801cd3db3351718a452738ed5ea7d63b003ac6c441ab53f538757d2de9bd3be1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h103bc2f409c6dcc4ada96ffbee79c692420de752f92648f475d38ae05409e9c90d0f754dfb984ca1f3a132e46c06f6d5e7d4bf431829e96ce3874a5932a41f0fccb47d8fa88d300109b20cabebbe744fdf2e0471179d84b9fe9163e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c6620ce7e6421c6ac8491ac231cf884dd432cf97eea87e6b2ae2616bdfdce4cf45ab4a7788eb581711e1f4b932934ece9c1b17750281db03f0d7387b39f7137190c072113a8065dbe8e96b5f2a0209d6647ddaa11244dd1acefa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c06b42a8b000b86a7e17026e00f000771ceb8cd8f3f0e22a6a7a83d7b2d6eca8c008136bcc9f9023a04374b7021118aefb8b76a8acee8cb30e78348a6dc4e5846c695be9bd1ba050cd89133387bc651b172a229a60c7cf6f511d57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad7dd16c9bf44c867f356415c246558354b5988f6e2570439081e50e8015a5b2998efed2949d21682632f3e2d26ea69cd64dee48fedd4dbfed954d95b28099a86b914f12b9f7f0124afebce11f5ede96c3ebe63f2f94b68e98469e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105d830b3fad7851d3b9a86456529518eea2b6f643d35c280d58d50188335dfc4a6ea0930b5deaf6891f109ad3d6be7259a9eb58da59d76bb2343042f226dfc2202fc9ec150bdeb0dac45fade7f33636830bc4d98fbe35983fb1a8e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fea90108b5173068ba17774ccbb1b21d4f88c121386c80efc6df160d18e8cc39450cba040c4a9deb2fad9ac42581bdc1a1010402b6ff11966d50dbb96e995d2d80d4020335ca9727fb96ab6dbc3bfa7f1d1294212ac11e8ec52dc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h421742177041492988377420cb4482ab9dbc59acc2059cd266d5467dcda38592c93b48ceb313c6f31d4d6c181aa163319b8521e7fb4a50201f26f65cea518ae4008fec84d2e5efcb12936a9a891540f7e89cf51e036f21869f985a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h985d05020bc161fbb5582d7f7a1064f21e66c0b482b16d5141f6b4eeeb70fe69318d8cd6f12fc624524a3debde552202367d73dcd6dd1de4d500ee3e67f9980acd9a57536e67086b648ded024ba49773f4d669882d5bf4c31c9e38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d1a9b4bc47b49672aa48c070bcf5cde48b375312b3e8415eac6650992e187f17500c619a068617231c41340863f78c0932158ae19d8e01cf0225f1870138c2b0d96180204f831c0d16025703779960b53ab47451a0cfd083ac41c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d82b9cdd71ef9a9e8c7959c204c4b46fe29cfd15cb8133e02dd6029e96a9039472cc11cecfebf0d12bd9c732e91b36f167d825c6f1eb8193d3ea75c5c38be6a2dd36b1abeb5f0aa962e8f7cced1f38cf4210ffae39e79fc0d5578f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e5fd9a7f38529f6966fee38c60b72d6e79100490ab0a99f3c8088465cc9264c12574038e0216bc19e3b1eeb1440ba0a1ae9e49b251b6d76977a49d708b2feb644f593c39aa00c20e28d30e6acdcf04384c6442c8ea35380a33c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53e3eb735025156e7a74eab28d332cb551693fbca6682c1fc11736c794c20f775c3b6e9eb6e8222bb744a59819c092edc675f171d1244cb3ccdbf4a5e0456f0162804458ce886e9b3eff8ad96b946dc3849cf5dede91b50d5adafb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37b3ef948f375731a63dcdb929ef2d26145abebabaeacd1cf045c9266122bb8fe996b9f3445468ed69bb8085da422001cf44e5e2e762d93e308dc9b4112f38bc8473a686219707de466ec588670b546857e6c8281de2d2bd39e5f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ea94b27cbd5b1b6f608b96fe9925b201e0ab1b25231dc747c754b5f8aa74a4ff6d92a556664ea9798593c6df6e8a7f7a11a48f51d8a828773d2646f9d75f719e71b6b3ce2bf65ae6a5926528542870ab92e3d57f2cff775f5b9c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6198ed43585bbcdf83acddeb5465999897f02a4c1211a1c7cc32a85e4954a6b038387993c14b782c93273ab77d28da5213fd0d0f8159b17cf1657a528b30856da9b55386e8f86b6ec7b1fd12f8d465d15906f56c33cfb61c6d332e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e48acd100528e8bfba9797b1b4e232446ed328aa1535870a451a44af0a7bd1a52e1be134d7ed5cadfec3f946c321e0bc6e69b094fedcd74cb89ef6732f1073df6fefa96eeb9ef2b6e83221b27e0b45cd92c3f5035d6ca72d31bb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168a5e6cdf0fcb7e48c033b6bc90a047f3178adc833c841ed631a92d1a139244e25dda821c633a2d042664f8dac156722790a5a5302f61cc996e9cc7c75611a9b4abac8ca44a338c8f2f6973b403bce70cb9348681c7046221b3a3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h337c1eee13c6a276a2a2b49df13818b7a89252fc9ca1284036f7362762a151b24dca463c4fb13572a8922ac26c1c8c84df1aef22018b2619b72ac31ade2f91fa1ee552ef749a1e1d1ff12794da6230ea6158bca96be2bdd9ea5016;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eab10a0d17eaa3e97e4bb7a69d1bba6b08e81ca0e8233b730912def21731f23c2bff3de46575212e2326029c300fdd86698c77c4361d4ead25ae5ff1fcad3958ce208274acb4584ea4c913b2389fbd47077ec773dbdcdde922cdf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6940f2f742023a500892d04678e041ec53b65bb675d031c1ecee49ec49aedb4df7de722d1292989250b31276c5c099ff9acd238de4486f7e35b8bd92a9cd59e1fedbf9d59d710d28a2cffa09447020ac0d9f0776704cf1325bfca2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95f6c736acfb2a7789637a4f3eece27aab6c6ef78676539dc9a15a49bccfa6cc93028449205a6aa9915b9e773d80b2a48898a23522d44e54d94489a4a2cc797868c707612702ae1a7e2759ce60a1e29706001893dbb8530f55c1f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbae0028a4e27b6153082fd55a27bcbc984be492c7789876d1ae58ac7a8349b571d35da4696ea97a4116118031b4e9ad7d9e39b3989d6e01e851100481d24cd46b4fc542b98d8123dbfd5bd33e32ff3e903a6ee88b138d107b4aea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hddfd08afc44cf26011a087b140426808baca4facfed403d52688d19df357a36ea8799963a9f34be04e51976fd1781fc3372e0b4b897dc0e47b3c034b6fe06900dfc5508da72493678ec2144f03a8f687fb0b7e0079ec51f2ac11be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acfad944ddc7e523ec8cd1e2ef0248c1b344c91f221b4349a76e7086b5a2bd244d5071e87ef2056904c330a6056e017c5946ddf27a46d7da82084ab3aec795d3f66e11a5ccabe65485b46205c8835e9f4755fad0a6f27709078981;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c82b4ebd8532317a86c96ffbd90627945832e14347a708ca1fc04d828287b1294de88065185147f8cab1ea84f07092c2f8ca2f6451a6c133ff7ce8371e5692c6811f252ebfe73480219ccaf366ecf1b04d4c3983c99c9a0e516d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d0432c33ea2d13c4e542ce7257245dc438cd6234becb1045cb882c1cb47e82e4f900733420322c868978fa8ede692d0424cc68ec76d56745b4ca811ed2db0c8098a316b0216f7eea08c2785b05828e52d9a56f91fc38d60934ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1bba5bc42743920b47dfffc026ba962ad22c679b0b049d3918a45f3b3904c55c9c9d2693bd50a1a24f3e9cbd81d099056fb701bf1b5407a67e65dcfead3efe070b59952962deab063f7c8a7e99054d13c14bbb6e30be2227b5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195cba6893450f8abca70b08277001773d25dae2ee17df13864fe8dcd25090a256e5eb3d5197a10f5dc1c4c68bb310aded4595555ad86f3aa72b13f2b8f63e209905c92becf5896f8986e62b5cff0a711637a113c1bb8d84b5f6e4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cad6dc8ff4f4a7d0640a5dddc8eab49c15482ef625deebf472e85c0c410228970d9906b5ec447f4a3dfdbe27e235bdccd607a7076faf98ae1b7d671d700fca21e1fcf3592bf6746af2ab09f2d40c5eff31339fd31c449875466be5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196209e568452455db081a78d2582766105b1c50e939e496a25b08fcb9884664f4c6d4bce2b788140c31c97addccd1610850e66f344443c5eda651e03a8ce93254ff19470bbe3aa3b0ead8f8d85fa735bfae04f41e9426becef6df1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc36f9684feb81f3103548b4e0542e3b1ef8e03ce518f6616cabe369596e8ad8ff850fd2578b8cb45b0148d8a589caae23045f6db463e212c4054dc7e2cc4a61130d6238f65af99f94272d8f6fd5dd85e0d064e9c3269a15073c090;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162d0b41893e20e6a6ec2763bf0dd359666becd32f41b53fb67c2b06223a085255c36b2d56628070852354d221d5041b286ccaf668ffd2e0887ba84810346318f07a33c55b89a2da328c54e5f51bc56809cd09d000afa2372b3af5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d324bf923f9383b79a102c8f412c75f8cbbe007198f9849e2240ec10823df02f32c6ae12c14059ff2f6b398f2d8dc7fe445b364577a438fdd750488dc820f0cce012a545452a8fb36e454affd06d087eccfb841458d46a5eb274f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1e1f2b4915ceddc0f90ef46aa8580e6b5dcca32dfc4dfd6ddaa1985213b4f0a31c612bce1b3c3c86b354f2bc0c7cd8c4a5a9058c1b6b3a7cda4e9d695242e21470b4e4aaba994d54bd8ef6f17ca77d4bbbb119e0b736ef32fb698;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acef98c345d8f742889729f4376ab32f72f13ec7c3a30876a38da7c1f767800f05ea5614c105d39d523c8964876103bc5e1680788c3b9c9206318329d18f478d80c6214e012a39eaabeae52e61f9f446051948c04bdd8e51fe4892;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe55c2319b77fe9adb2652e51fd70283e3fa560c8db3fc9f51d5eee5f10793a2359f433d940b6796ced8c187c1b6666d0fda2c1e9421ca605bf5b9c2f3ff7151c5ec3dde623b7b4f9bff8e096c215a7dd88991bfee1048d64017fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e14a3b07d0191ca16f2b65a160979467b2eccb6cd94e63918f7bd1564d41dd37679dd68e1bc704bc32b604c425235bc6472647605c52848c99d8896927703a3d9ee4aac4f0155bf9190ef342924e84e8294df0ae56eee2734cf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ba38c68056c7787798eafab3ffc48461f757bc849be327a981ec00fee790e65793725ccf290e65036845fd971c034136f4f912b675291576f337364d441de1831e7af6ad871c67ac43a98269c5819d058a30fbbeafa4eaf26674c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd77872fc8b49ae2f4a447fce5458442b4a051a37f30e79f13c1231357afd9735c3b6a3608e3ad7726675fe1b9b42fefff002eb44ab55059c3e50385ac858767eed4e159318aa31c0cb2fab27dcdb08c56f3d2c9502bd4923e51ab0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78e8cb8d807e39bd54d2dc6808f3e635a621eafccf353e2abdcd714ff1d1f9366db9ae719c8a1206fec181ec648702cc1aaaece726ea5c606fc7ddf8ac957bb894b784bd32ecf562395328760865bb0a3df6b425cea2e581744e49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2166e39b5f6211811d2bd48f5bd91f8f326f4e336caea6a7d2a1ff4757fd5e4e6987f1467a0ec91c755ce60b4be7997b1efb4fde3ae85ec95b6058af91f17b11eb5f5463e34278c774fcf9a01a7286353650d6305460b0a5c6ef07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115ef2da9bbff92c5988728e315eec0cba5bc22133bc8fc06dd82240e8b4851959b4a0b3adf5a576c650f7de9172417f2f8aece56c3b983d7f333c473fe64127a046f1084f0856c7c9dcae3ac0e2b935834a3b2a269d25502c48b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82f8e3dcf1d991b1b644533891d5ad99eea2434322150ee077ca892fb851fd8e709722e623695f45993dc4440aea49fdfc123c13877d38256037b505d44c7adfb0085cb06305eed02d349fa6fc9b2d140eadde1877166ae7078ec9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8258d7e772513b29f1b63961ae7da30d7e72afd6cbf01f1e1917322573729da2c2a247521fdafe7d5b071d9a8938ec533bdec629a3005efc241c3f9b9a1e47fed34ff2e9085ab69d0abdcc3848ed998531e437893b3bc295cd5eba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125bf29d36189f7dd904884db5aa2b94beb7f5e33206c475499533b09e84b3e7d8a57715c9632fce5735d5110064abbb5b7c8d1e2a0a11425472ddba0764a3fdd6f191a4b088c1fbc807c4e8d75895dc73160dd69f450e17529ec1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27d426b253ae9db185887e3892d8db94dcd8f99e3a2dd53427fdff0cf9feb69851eba2ddef19fca532e83e75c4688672babf8f58b4de85b10d6504364fc14147c530750e3175038f7f6971ec1a1f2a2916eba928c8c3187053ed02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c12ceaf04af53ec82d8c6823b38a9a8a6246e1666a2cfb29922985a55838a3a8453e27b34725b8c53fcda643fefe29e47e858c1289c94624a7a1d28350d381039b0b0fa8bf8016a0858bb9dca124ee8f3070739371ff3d558206b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8c5316a97219ea71df8aac7c9f094fd7d407bd0250e5f811a6b29e1fd417106b2b4ac51a1a1c536d388c88b615e2f4ab54d60f71cd90ac89b483d6e50b517a9c1a115fdc95259930664658562b8b004ddc6dc05e3b3be9ade134c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6ee14be0ae9aedaf870f5fd6d6d743f0ae31099fd2457496ed26a11721a5d7f486a5fcc6ce8d3b7beb91f154104a59f86f0489c3dc06b26cc61f5ff5493fb62063155fff22f75952aa41b1d192425d53e870d3ad7ef1722d56084;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de81fa394a960fa19592f9efaad33f076c085da8b956a8d208b8dd3974bcc237ad336a46f24c2abfa96fcf65914e49fbed727fda173ceed6109e65c7b722af19d2fb5e27fefb91bdac4d8dd2b4dda6f8947f2e7833dde5f45cb6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1238dbb74cb5ca0ae1052b18e93f90d978281a5c58252b706d1ecb304d44df9bdb1bb66ee782a68a712298da7472f099af55db8de480cd001864424dfff936e5fa991841bb19cfa0d01a54260351ac2010e568cffbf46ff9659bd29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98629bbe1a5899344e146544dcd8af3168202374d7bcbd46aee1ffe1eae7fad911ad90358398f5535c684f4aa461a6d6ad79b132ee3d1adcd2a0b458cb5665f6997edec7c9e56e2b945db8feff14537e68f6d9aac627ece637facf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3880a6bb9ce0af5a06ade7cd68bca39eb734c17716388a17ff0bb6d614f11209d0bf25a35f63a3541b7041924e34a249fd6a73d546d6bd6d77afd4b58a3352f53c3c2a19585e48e4e49d7e8858ac72e0e42f4fabd4b3c7e479002b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h616c802f8857516d5cd10582c910a2372cfd284e53e39bdd731dfc5b17e9c673ff81b0b776ef68992adddb63d58768c8e218cfa16b27f25dca3d93b5480712d276e4932b9cea1293f1a1198c31031eec05eb9922eb3c9952955629;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3db796b7735f979b9d798bf01948e5224bc1f32c5f073867b2de9c9c6876aad597e08ceab9dc65339fc6cccf174cd1f4c435b9273287e9727891d13e4603fdbac21e2a1b2621a8f98e14532bce878992addf37bd8ec04e7789dbb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10449e70c627e81f3b3e172cde43ecd062eb90b1355761f80d09b046238b3d442081767f3f3bb87eae2ffa4843d4852b855c88c608a24a2d8604580febdafdbc08e6bd84af15c692373bedd5b355a674fab45f459b993ad1f5a506;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf25aa65874ed0ed071f881d5b3cabf134b818219cddbee6a060e18eaeabb1b526fea2c998ee723fd47136fa5bd3db8bf186119e2d209053e175b8505bd1b059d74709c73c939ee6fd8888e4d0196a38fde5b0d444c8b3f23badd24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8eaf9afaa180b9c73218de2017d51149b4a19d9fca56e7a53915c4c7cb967586b3db1eaae077f8df30c92ab0d9d87bc910ae6c624547ef6c8d228d832a94117f0a22febed8a29b3d61a58356c75a8e3b6d674b16c497259c1aca5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1427f4586ad58907db684f400254296205a71c5bae5d54ff56ebf058f23893b15bb9b6f2512899bdfc5a4cf9e46face1ce2e564664a2a82aaf6369fdda57cc248e05271c1f5afe3879dc24743d6f48b8bc4d78346cad54311621105;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c1dc6203cfec6f0b0aeae26e497d85fb7e1de9ce506c31327e2a9675c5bd35239ca7b678801abce4c3b0733e9167c0b6fecb7ae025ed5762020db4641ecd92d41a3728c2ba1215e483f84178941bf1b2f44b01a9221c2f9930ba6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d2b17cf19767c97cbc9bb6a51c35b2becc9c97fcac9e5801d7aa9e34cb46643ae800fdfde2dff9aa15703d92a771831fc31ddf4774b5e0e8828eda9d44b704251f9f3b38ba968a6c9f7002ad518f0dae72eb099c39e50618728e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1821b86886250753419ac7d279303a66cd7a78711ad4c2e0addac9c036d6775026dc56d76708f2e8094a029ec6d54db5c70a65ad0d2ee583ff8b8230ee411a13d84d7aad09bf5d054f789cf6273ba3a9a93dd5a722eac2655c4ef3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e881c95583c904ca2b5031b382cac04336e6c73d6c5c24583efa2ce3d74ebd03b2b25ea9b9f1f347d12c97c31690afb78843351ba6153649825066238251664c72ad88f3a65385525ca3c636a4f36d158083a13ae99d9ec78483a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he91810a0ef743a2dbd6ff5772fab24185d7d3888dc86da05cbd9a0455f4723935ff510585615090f72152b6aa67419f5db1f7186e43f77cdef22d342d5672dc5696322315bc39f78a57c4bd8be8cf02858ec8e1bce2d1ac3d1b15a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4db595e4e6bcee3f8b7399ccd7c701af42bd9fb4bea8730cdd10d19de284da657c0c6109822153da231de2af2a676c42ff42ad32927ed0b3e965a257162ada47e0eae52ae6a7e7840a6388643b3a09a4cb0d09e92f86fab73d69f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147966c62965ab42afeb652c296407bced8be63b71dd4c1ee36eec6a9dfdd3d919c4f30907423dfa06c0869d03393a566b6ad00f2882800e87e08375f13f593fa94a80497a2b6594b9eaac05228705db35bc8dbdddbd90e0ff8ce46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d606cbc3cda7974eb91f2e1d17b75aa480de0c84ff56a36226a95cd98ddf403843bbbe6353a278ff7846a073516387a9606425640b003ada34ca17da9b2ba265f4c22a9458e9ae9f092e21960dfe9ca97c32e3ead54243d6f847b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16235421db434a9ee4bf28a421804e07d4ca4733fb759bd288e62046003bb386ad37e7067ba869fde31b69a8f5537c22ecf3cf09e0e2ae2db34563e915362aa95c0a755efde1c200e847d435facdd47a92fc78b3ddb6248e148bcf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1838d55277efdaa1b58990980da3f2b482bff05c2947c08e34beb958aeb0c823e7eee7ed85c216b0493f10b2ff23a33485d377f9df5491bc30644bb6c545769e4ff3ac16649dfdd9965be49fd4640e4b68d8fad86ef4f8d0e6879f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf5872374f5c6b5bbab1a02ad4177c8b304247942f6c50649616a497673776b4704880f5b2bb775d0beae93cc2bd701669eec71494e880f40b26f8ba1a3ecbc1aae021ab630bae0a764c575a46a0e02046fb7934b44b7f18d741e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2637301d4f6a9c4f2486566017b979c503fbe1bf1fca60d28fc70f034ee9558a505402136c279959b895bf1a313f36856ad5786c1603ec4d8a95f01b85a2d93e233415aeaefaad71618d9df71d67c527243be224aca1cb8e6e522;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9de9d0fe5863392d018bcda1e6f4143a70c602fa953c9ed90fa30286f630a493db45ec883831e53286fbaed3fb65fedf0c0c8f521489ce854ba2f7a3fb9386e5ce60aa45da3223f82ce83c1eb7c2f770e40cd5c7bdb58e5bc239e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6236b5b94b350d142bb83eb2a6efe36d736a62b0e4dd0f5719d7d143d6b92ab5dabc2a32a928f5da2d9dfa7851e5d23cc63b98f9f3a86ac1ca4fe619834ebe2802d8f6eb491be5940f2563da3b4517e6380a50fed869f36479bf1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca18988244901ea858cc84e1cc98fe665f3d23105ae68ef4f0bf44a11c942669a07bebe1e8b3240216e6df3293d0198d1f5dcfa414acbb0eb9884dec0316c29f921fbd326ae3cae7d8b8da58d9e85a10312965e2ea28af0dbee045;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196a9756d3164e5f4f30e774ed65d27b42af865ac1bc7526e0da271b55d40d8300fb54db0d7579ddb7c8768cd83dd1d94a5c755e4e095518416cb7f46e38de9ec21c03dfa709d043e6466d910e100637ac6534d47ef0606ce48eec7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85c7ea140289f33301c3430b4e85030250c4b275dc66e287896950ed17a190500e66dd9acc8d09b67c4fbaa66aef76728b8d3aa682fa8dc1a8246558813f752e4828f85a32a3af4d35fb5cc15f45059e6c34624ddd89b56506e3f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96236414e845fc3229746ab61666d1d3cedf7f2e0ff7ad364dc1f0db41a93625c40fa1f3d1b16d2fed91b0b807c7b324a41351774ab74fdca003a1ef10c36e0cc6c9e9b64ba314cfe64837c985cca040f20eaec2dab2905044dac4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c026c05f02bf28f3d571a84e10bd411836f546f87a96b8adf325384702350368ee08b302d56fb1e3ecb26d14cf2e55bea20f7c958b80629149d5b3dbc1aebe3bced531bfe313754492560bc31499dcc5a9bc8e9674d8ed235f376;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d071cfcfb4e14f1444e725a2751dacdeff21404586cf26fc4f90338942c2a9472f230feee4e2f667ea00e6c7444b23f2eef830836b5467e966a1ea5ef994b392f91b1944c5f343d4a32aba04479e53e9f8b21e28780185d3de6515;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0e8071cd6c86e4023def72db32cc6f60f16c498ff1d167af8d42bcc160cd285a86a3d33536dce6c90876591b3e50b19c5cbd4c59be27bf478d02340477066fa165f5261b0b7099f6be4475557e18f0d6a4e9afae6077efe00a699;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4070d31d355c4fb8f94efa6b21c13bf33ac0e05f79775c54c5c7c78bdfcb843ebaa0b892b24be4ea6297ed8bfc58f1c3b6a8e150be0770178ed14dfed8ca26e4d031dbffb0f50e49703608689bd85d546d3b13ecfccd4eccb9e774;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c801e2ce379f4088cdf5866e76e0412f0bc8b64ddfda24d0f1100798ed4975b59e1d1404058584c4e1e1efb74bd4baa3dbe1e57311e060b860cb411d758ded329a86b8280b4c8993b233be511628f8ffadc9d77e0859eea3c68e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9fb8e788e9c548f9f5549a179336eb83535d19c56dfb2ec711a89d63f69b3d6725fec8ffcb6b4d159ef25b050cc9eb6a7e419319b1b391366b53fd4797531cc2aea692329df8d36dc90bd8c738312e1bd0a967b7e8c2ebf45f4eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h938d2e0ac03a954a67836b120803f6719c40c2f506f6c0872b4817a4a0b16317469dd2f5344181b93aa03295b9752e2c132583d7af57e1cabc20fa11909364e1c5e20c21eaf37780edbbd5b41bf806103ebd013d42935d2e0aea81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d4ad2835dfed23a5b9b7683c59e7133ca4c992581be8a836042275d4db328ff4682caca1901cf5ccea26d99e1fe676c1f33354de1e64bc0e6c767e90de6bae1258e5853f9e83550fd63cf17ff0df14d8cd2f267f760a774253008;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd40b742d3c730a4acd7a364683d080b962d2add44509b97ea9060ed1e0c9d78c03079de5080ddd898170ac97171e66644f358564bec06fb2befbc316c146cafed12566166b8c70d8fdfdc01d8a1697a9e85097c2c597c26217e351;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17253cb7af54501fcf8727aec6494375182d02168037888df347694c7b8a3969420c5d718b046aaddcd001efcbdf5883d20478a900df2f1cb881dc38204927c6da4c8bcdd7bc14903ac0e02c1b92c445ccd1b49e5051517fd643615;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ecf4d91e339af68b65d9f213bf1ed25d32cf2f80c46886aac956e9fd84596bc5141e4d0cc328a96a06686555732a797aba92375c22cefea14ea57a05763548c40e48d69f820236f72cc33627c64e6e23ae059a39bcd9af14d9924;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hacf862f60b696ece77c00e61134f08d8f587969eb2717c056d0090a0c759213bfc7ca863810f6b5dd4e409dd56a454c1946c07cff6f465d74813e15a321128c2275288986ae53249ae191a4a8f3d6ea9417bb1ffde69cb41e749b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181262ecdd742863d7c32b5727f9d9c440d6f7f1f86650600b6e6c36c945bd3dfed4043710eb4c2c72a798fe59b3f40a773a661589e8c5850de5cf2fa3b2370b6c1bc2317ca44415356469b54e8a0dc65652b314d286e0336aacf51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bba6dfdac702e078761a73f5d3959bed96cbf99e5e427196f63d3ba1c53890c67a1564701d5fd565a69d43907cd51d3e12c59502d6b3938bec85241f31cc42180a0f0a0f5aefda0f4cc05c6af228c66e6fc22bc77e2cae3db73c45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a65f9dd4fab107e8c9707cf18fa86f423d7c6d956be7eb00668f241ba45571811dfd1e0d737b7b7dc85c9e9aa8b9d2857449c48bd9bc9d7f12dccd067173f50f2933e5fac8fc25e6911c11275ec2a9c3d6e25ca114dda11ac09a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173370e6420bc64ff13c9ac7d2d6d9ae2dd51723eba6aff746c21bcfa8415cce05e98812e21176f9a512dc9588db8e54d9385b0af97f7e66dc51ef54e02397ae6b256063dd6449b387824b28e40db02e3c30908b59387a2553ae0a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1623d938b44f335f7555e0708c40d8dca96e8a52216bf34cd42721e4893ac2719f395b93883cc12520dc52495da48a47d811ecd079206a5eaefc52b14efc2c24a8e64c78b3010924c8962c9a9a4ccf387558c91209bfd878cbd5cb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcd0019e9674f0eb7e1c47264c3b7dda60027ea60445709e882085501f84e867c03140cdc27e81de3ee90d94030ed0cd0dea5f783a608903a0f6c2d27f460f8b49948da927c297ddbab3631dbf284d0354eb31af9c60d91c357899;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16be1fde6d344a4d1b603a8fb0db0efc90762b84a364e9930163ea9c5a4f5d1f57dea3688191ecba3d7f61c1198d5f93b417f6878bf3c90507df644727284b91a419f052d8184d341b109da3e99531d1edb2f872ae83116a8ad2019;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196e793edf5958f5febec8dd944027178ff6e42d3b0e4c10f4ab6cf67d406dc5b56569006b2f6dfae464540564a684ff006f03ba03c6f955dbec8d2243dc732dfe29d55d3569fe39912afd2ae6f5b4225d57e51f66b814969459d20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf16831766241a77f733882e26b303c36091c628c384a963bd4aa2622b74ca94972e647f206510eca85b948f35e6daf4c34c47adff755e8108ff5404644ea2928ddd865fffd2caaf8e1726fafb08ae098b51abe1e04ea2c0b6e5554;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a732be9605a8ae6f863344588158f611e30554b879fce300eecbbf41ddbaa400b7dd5ff4262184ec5e062d16f31c7029239f05102e29292e3636b0427ee01dac0f60976db67a1533df7be58ab88635d30d3d24815e7254b401451;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f02507fa6ddd35971b39688b369e6e920e38e8bb48dd75be98e94e6d6b113ac30419ac8b2c44cccbac6b5734000599748470b174e31261bedea125f0eba3a08c0ebcfa7f1f40e16126e230a8ac8cff9cb3d5eca559f807e9e07741;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1938b22fbc663bbd231a1db3a05119461f5311f6376c89e04488cae955504b5fdf8bd79ebe4a1df3bb4a7f29a73537b516bf7ed84bf2c504498bbe0ff1fdec161a9a5f5cf7cc266904a10518a800c2a54e48dbd210508779b2a048a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ef13127b92c552253858fe70c251cc826caad4eb6d7671cd061d20e567217b815ac29bac8512914abdd5a9e42b97444cdb48a237c9458f83fdc3b26cfe967602984fa45915929e6c971431ee61947c2512543de2b8d2d0270c3d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d54090733d63d519eef0a8951ba57bd3198a3de4d5f289ca94e2b8dddabdda723f288c7f41c205ae6cec4e58e64916cec886dfe1e1e6389a3a04d6673d95508c40e6d1ded202da762f294c783928252652295cf165f3408e5b6aba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h876f96fe589929e5fa1ca9b24917543c9f5546664f20a2bf2a6c4c4ec9dfc7f263d4d6b33224e2aacc3c5c38a12b262253bcf3748f897a6f32153c69692288a797ee411c1ccb122e7fbb78d2b28d1eba0a8389ea5517b166d91d8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1320515592fdbca1ff3adbb06cf1426cd722878304655c62ff799a33df31337cb738bee654132f025cc425b8519cd71d0008161e07fe5e424109050399214f2bb8bd4f562fc46d909c5c87ae9b802268d4cade130125fb9c324a76d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h243d3fd7441b21b481a0eb0e7ae591324e1791c99d2ce9fc844f1d2220c2244e3f8eda58c075ed4fc7c5772410365b0636fe0eb9cefb593c4447bde821fbe5551c3e2dad5a30f9a314f14d0fe1a06e48f2d99cf756b1a16ffdd9d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbec3fd53088ee798ba85c5b25f12d0e08045fdc4f61f4b39402a0a1c0e8a8fece962cd821f2b453d43ca2ff661ce40fc0afcd5372e17674840066bdae4f1dab98e19004d6c36a2d523db55edf7efb338a5287c8456f36cb4f330bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1deccce54e6adfc6145abbf309d72448a0593adbfa366c98fb36de1087b1a85abef366d813785284a0af5d473423a5fe0e9d3d6dd3b085ca11a521dfdcc022a5e176ac30bc381803f34d3e3ec851866efde20de1dc4d7a2b19adec0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19619c0abf12ad144575e6ffe9c5dc52b19dd233abb0810a19bcf57533a1512c308cb60cf93c48368d5567f3e20e3bdea1d47b5b95580cba8c7b660d9975a85386d3dcafcb6db1443717436a9cd4819520edee55ff6cc2c05d94901;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c2fc9ddb4a8ea319c2aed2f0b70a8752bdf86530f799dcf9d172563afd13b4c30bb32579f006248cf86ee114b51b30bb7d273a73d37586b08beac6692d5d809ec00dcccbb04fbe29ea8d08ca9ffb9d62e5bef0fb4992e4e4601f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f47d25d4fa7c640e35114adde4bf16b18bf2d24dd1841127d2bbaefaa940745631c0620da47c2cf6c0183a204e372b3c8d0e7387a013f171baa086d46c09d4c7828f9f75450cb1f88e75a0175fd9780f2ba3d651f86dee18e2c27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164d478539dbcaeea39ed91de543f2812d0fae6917cd605a93b2a33320aabf3b94e2200b046e16dee679dcd55d7ed8a2ea260b572e081615135eabed445c49bc4554fea73ed9c155e57b8aaeb71d2e956046dd2c6c1dca3b880e77c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ee0b42782a85c30fb2d62eeb30488abaed68b8b147ff35df240c50d18f1e9a12cdcf9974f8797c200a3f94a929b1c4b523e095ffe7e8de36bad8b187afb702d8ae82a2a98d36f72c15f1ac400ede884aaa3b6610a4c9d6becef2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e1c446013d8e3430f9d74e2bd8d9ffb00197aaaf3da6e15b22e67d98a86371be491c803768abd4681e5e90a2b9cf2aa476d7366ebefc67c2097931d07e55e5a03f16047c42b34a6313ee04301ee9994f1cf6e3c54e3c059660c93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16aad6c61a2204e05aebb62e601362e44109ca148a19fe989cae5c321b59b595706c770e5762c22b79f4f5a47fd403cc8ff88428331fe9da966e81da924527a192776d9e4ed3a1a9b88edb752d37e91660b1a946cc9d2f556eb902f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5d0425909e1d4d91d5c44c486c9837070d062a2504f64baa04887e66d8f6fe967adb8f10e92ae94b390d8ffd5495d79ce589144cbde9296c14863135612cb095881d0793ead76693d0892d9fb385bca924f1f82c9813f61d72852;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa593f641582053b06c655e286e3d40417281fdf2aca468816a58af794f1e1d006f6ead201d3e82c7ff82afd20352345ee96fce63ae1f56f41be0b1e9ef31d637ec2e5fd391e7f96d09ea1f42b9f54aba5ec66c208f9ad27dc967f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc1de131a2d64f8f3fad0fa8176d2b14d1eef6fc32a2c3290af4d73fed773fffed2d4547fe5ba23765aac6db22c02f5e023402b58d54afc67dd664b2fa0d36370701de055c18f448fc192fd5a81086dd76fa7dbee926a287d0b5e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf1ecdb033f9575dff0c13718d8048c934c37f589578ccc1f0a4ef8fead8cae0dcb165c3522e393011982ad11d03d38ea4ddd668aa702d3604f9d5e385474ea7e6b53da107a32a5fadc8481100f318fcaf075290463664e8090d01e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccd7bc86912cff95168beba7420a31d8f791df489a5af57a75b84d2c1f876509e7405d67e50b17760d7d6cf285c76f5fc0bc2102587e98ffe629bd98420fc704f5d5a8284a1753f05ce798dbb6909776bce90f61fd306a33f0ad41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd5d8c30e78b2ac86d675b95d098666166219a558cb50e75198f39b71058b2654fb8b399f35459db370436bc3ef4c6ec6bfc1ed5be907621b34a00bf13f843aed801116ebc7da64db37fa1f795d81c66ae761baa186e958c75cac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188f5877ef762afb3804ca266b36d507a10ef3876fe48803469991b058c6512b317696f2ec1195557b9e3296cddb3103aa0e292c4d25f841e7db54b8ef77330cfdac32f8f129f13dbaeaf6a889970fcf8123c8502edf7a737a6f34f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h765d40e0265c84bd6a6c19c0f47120efeebd4fab75bdc0e76b7ef9d61c00199333cdc0466592cfe0e44f213f99694dd31fd32cc0c054aa2c2e8e4f3f0618049f187b158b19cdc3d735e2c64e9c77ab4e6fd72a0ebd9501ce817449;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d75988f4d1ea9a9d266bf7a23c8c751631533ccfb58a40931f5d7706a5bfcac42ee4155a2077fc6e7262591cdb1a93e9332573856f79a9405436a2aafcc8cbcc17c3c01408538c2ac613b7016b80946a1342971956f1cc8de2e31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1243ee73bda48e0f35bac9014f8a5094a77e51726e1238c8f5d652e5499c5bb9de8d3b71a648d21a740908515519c188078979b38d97e00892d90841cae452a36bb634ae79366bb4b82ff3c8dca42c4992569cbe9bee2f0d8919f5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b258c63071f07392768d2663921a4bb88a90d1ea51c875ef976963185ec82a70bb977c09b0255fa76063b8b2c8a4c4181c96b3e4283798d3ef6b0047a45fb03e04e8765e24e453ad9949aaa1fe0e23fd17c4796ae3da49cf4bdb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a150b09c35fe8b92a54ea38d53d85844ac650f2e2a40adb80bdac706bda109729152e013472a3ce150e6a9b39d8dbda025a0267d824d78c4e57056749879f461d48d0ddfeb65da61a76eba011f41ed413494e1297ec43b82f37db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h902215809afa0a6e4aee5a63a68a109706e344b1df27a397b8f140c3284bcd8375cc6c6cf1a16421035a4caa567b7d2e41116047d86cb56443e02c3f0ca3a8ab3828eff06794419ede45efee4523c9f5423f890959f26fae257383;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha31f4809444799a9d60a9d295729a9e48c756e5739aa90acdccbd8e7e125a5a8de928f164f9ce66adb920a6b56544d24b505d8bd4c057e8571cdc603c5813040e58771e6c64f8046d44df010c056997dd759d98e80c5258c554276;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a439665ad1f3cfc39fccf871ac5e357f003fff474a16b4acc55ea74d9b92fa2a2527624b3c94f1452a35c826526b47632702433af9a15ce03403ba642a62f314ad53e5d3c7cce3a2a9ab0defaf3d1062e1d6cd91740101048954;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf07244a968c054742c4e07df0d8fb3ccc67ee2e9d93d572ff0cc67887b522455ce173ddbd565305be3071156fcbb5b603ff96442ecbabf7bda6ebfe12cde7a27e745ac8ea03e39be2f923073c871c74f9dc4e9d0f2c714e25f141;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13004208a8c77279fa8f631b3ed2b3218aa3a6e69f52a92ca77824d26619f0165e123c7e2571923fc17934420903c6c67ad08bf330635bf7c6c2fcfa6cb7c1dfacbcc37e48b7430189913ca0adcb9df785ea85d696e124bebe1c0da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he441bc91bf9e493f6d68f09c9598d3320272bd5dff6e0fb791c9dab4546dcec69a5be90fb118045774e43324e8b9ff654f1acda84171a2a70430ce86e0abe6ea4dd11504bcbffd905383493c8d07b790689d303fc3849372eea885;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c32e35d4791c40bbf4ccef96efdd7fa7826c6321c1d1b72be6262bf8183cee99418ab7ff1338ea529b433027652f7ea36f2add2a23c72ece3bb761940697e36471dc9f8b24c0b081df0937d7545243f4f5570d5207046b2c19223;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c9a2d3400f5b885baa055924e4e8899eb738b6cae641d3245abd99e040e3e0c6c31ac604bb3fef5d03d42fa58d87f600b6a9c219c63dbab0a0bcc4cac57ffa74bad7e4ee2bbbab42ee439cde658228492eb495fe5e5b7eccf7622;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd49ff9930e9c6475889b1e0d1347c98fb3020823035a0cca738d4aec860a3e8e1292fd525462173473707ba6d2c323521e367c068af43426aff488b7027e678b18485eb61c857a83b6b2021b5a390075f915c967c9f1634de9113f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd35bad7acd933aea5c1fdfe3d4a4b461a84052aa777813c94b8314926fc80aa1f9bb2e51a318a246dd5e453c1f4f95f7e9e8aadb2c85585e1ba203c431a5651f7447daf6bef2b3727c49a98f22d03cb16c988a2a551bd22a8ffb68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17937510c707c2d329e8442dab8746504c773db8b26ec2f22851ca4fa8f7b8f24525e131ebd12ec4995ad3fdc5b5e06ddf7732f9229f84109793213248b20f8fe577f6c34c9e9d777b8e2d19ac8c80e7c37a5cfe91952b0673b01ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e16cdbd6f5a9074127c6391f6a561132db17abc6492ea1c55d8c07c2074d127dc4b0b02f981c38346bde3c6a7c5156c0e919b8c7b0fcca97feb693a69f4da7d9357775d0943ae614c5df3b90e74732f748081051dba8b0d8a474b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cfe115e4bea2b03cae65f0243acd9efae3fb260f8f0652e7dea07c6b474fa6e6e754096e14c6b5c6c6877b73075aa703d6d092206300fc61f95fdaef11e1f11743be0856828241f48de2300491888d77e5553aa16a21b93ba0cac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e949ca49a5d92065517dcfa453b9c236c041e71a5db2e2e6848ec0a2ecf0d81eb43e8f62141096e881399d76b47cc7dfa9c246bb24a553a8f60c4ac79b05d85c68341bfcef6ae14117fb36580bb380b5fd033ec10da0a898db48d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50e955ddd280502bb79074e888c79b80091649f0005d85eb91e9f0d1bc004f141a8c9b914e18e75ccafdf3f12466394d917b7ae6544d3b6a138b960f07418673972d06dd65c0b7d97b1ce35c015842d274f1b26c08c0b5248c40d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd34c64da0d44375b4b9da0e559ff8526124e017549d3db6ec257bd57359c38ead0d1e5884804e76ba868e94fd079459ec668a87640406e38b8fe41ae3aece52fe90659fdc3fa0707b5a767b4c0a2b8aa91e1d9944dd3df21c2ba05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102ad405f80c4d14a9a120d790f333020fe5443137fdc58c2bb89798b7ad35d59c9380ac7d7cb33467f109a48696e60b335932e38e931731bdb5e469cbc1cf6550c582009aea7121841734d8f5296d35f8e2a57cc611f9f8c0af721;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dbd392e149e50813cd976f41a1605fc435a9d1aaf626b106da9424bbb2df720b1c23e0f920771a12fd14938130d7a84f224223b08312458c007c5dc4f68527a2505e928cc348e37e291a2521f7aa4547443d1de00d5afe1493b99e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed4b3a0960b0f98db0f20574fbb1c6732d7ec04c0b6fc2288cf4d8929757c0fedebaedb3fed43a7cf939b4ab40d9b5e4ca2ec9a611ce47d84a5476973d774acbc1deae831cb86d1f92b44c68da1236a7400f6aca397d149bbd5f5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0a0d797ce6c5f04c081958df87c167c3520def00ed487f80bb5d32dbc767aec001e687c83d1d77b7fd10e6dcc4f45e800ab74567e90b4c7a0f4e0bad31d8a93b71b1f02d562651d7033e52047d413cb051b47381ff00ffe8f99d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14db0262a47d062d307c7d425c1ad4cd2fbda1d7635a98e5859bc60aebbb59bce05fb3879976567eb47a6ebe9458798396974a5974b157c4020a0552a958f9e6662208972052acf3da3c623d6881d140c77804d478a27df913617ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdf1339bfd516da4dba5da2cb4635338f0f386b8b0a6ca12c2f4b41be302a906b36087db9044ba4f9c697d7742116ab6b364813af5d5d43b2e5f9bd41eee76078d8df0bcd5cf49dc9c12fcd18e97f1f4030f4fb5f9dd81b12fb11f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ecec2663c7a890556e081206342a428a83b7a5668c0cec61ba03252ea8b72ebf9ee0ea4239474d56613ba50d309e633cc9edba3d5f33035a74746f1923b7bb05c57692525bc49fec793dbfa69989af5b2a222d62238000d5ee75a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h251d6f23f67885c1f99770a3074c05ca4895d23439030ec2f964f82e945ba3ea61de74675ad1009b7a168a454296f31bd8c4aa98c1e99920317e40538b974523f83177d42f644b1a1e6155f9a1d2886b9c4e56ddd704bcfc5a4498;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaff26f054ecacdccfdb4411f5049afc47fe1708bd0ec323c9e613d6ef65c777b7b386a2ce2ee7403fa328c4676ac8b8a41bab73268aa35b86742c85f733c899bb9ba7b42b188802cd205f6265d1a5b82dce8245d84af4723ab43f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcff1414047ed56d8db62a4ffcdf4ee917108e94f1f6098c936288c963954a64f6a7f33b801a85b18cd772ccb3b2b964a02935a54cf053af8758bd844f0f41222f2f4be7d0a476a4a96a2e3e05a6aca6e7da1a019cd94ab5f1b6170;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1496865b2eaec6bb8ab87234fe87c311d2bb3c59e21b979699b1edba8931f1aa308dc626bc90b1b8f960923d8425963b3dab955fd40c23713e24e3256601bbc3e29639f0180ca6035b0c31e16ec652b0ec04f0907d42072bff5596a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he77f0f8db032458fe23af41d21f0b66a831a1a5ad747418c0323e0c9a2acf02614fc8e61c1630adf79fc8b7fb986c6cb90e10ec68a251319933cb287aec3f2ff89e416a5b69432fd42927b2ccd83ca56743a65b8e0008c44472abe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8892faff44630e6bec8a2105bd6ce6fc85041de86768886d129cd18154792ba1bee1cbcb7351e372ffe973832c1c42a2271a8566acc872ca4f1de98d6c33ad809c2961f9ab6231a2cdc78278836ad223d75f7249241fd47f07945;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0db77ab327cffcb1e5a30acc0e2b3851afb2738d66f1cc06cd08d4bd2938caf91da3a9967204372c364a35df28bf901e964acc91b078e227cf6c79b5fd8b912cc11eb8e22592dfecc33523b1d1c5d228841bc3e108c8212c5dfa0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf08346d63807ff06165bd05e7cba2a2f4e842a54ceac8f984168bba664b3ecb2ccdc04c5b25ea0eca8538069c20864481d550d987e04a578ec99c5f527de04ce445cec814d85ac07d281c48c24ec373866b526c88ea5691b1b545a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e10e83588689448a513814e19dcba0e3b2b790e8fefb0c31abdeaeace1a2e72507e10f97fb6960424a86d9dec21fe4ffcd6f4070bde15036f52d8e161820dcb5d4ecc9de0077c99fe5873aaa142bf78b91e7f09af2c59545e14b7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5699d962d5c1d3e42f982f42d05d9cf9a3ea14ef951000442009df2e4c368a85e10c575406f6dbdb8dc40c18f03153496f0e480e143f732e213586255c37362656454741258f54310a60f7ee8e671dd11cb05617367ef412109a45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9c6fcf58ae6d2ba5e0841e5585f3f383a2d651a7fb02d833a66859c84ab0d8c75c31ccbfb1216bf417141d26a7dc7e4a364130eba22863f721a69f51b26249cd854d373cac7ef1a09569c10e2eecd85605a0f6fa3322c82966cbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd2b10a810d08a94a0300ed592b4c288bfe57ab142f01978392275f80f9ed0caa8d017ef87cd956be0b81246f9e7eccaa87873924b75eb8f078a6ac4ef791f8d34558aa57d0e5d306c3acabbc8d6c32d88faf553dd1e391b602c84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3295c123574cc0614ab1b3e2eb717cafe2488893e02975b3228070c76b61ec3e78c2830733557923d905f9b0d052679e5b73ade4e7135487379379c2788baf9aa1da331e7bceb170c4eb0cfc40030998bad7c2d4a1b9ce785f0fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1569734e27277dec2267513623b1f4a3428676f6a15bdb78bbde54bddedc921bd3e6946931228ab41e3b9d92bcd615a539f536cdbc7610e90c961c3f59df2153019360e4388e0f8c57d243b303888bd37eb081f0e8c163e2be0f2b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f44dd76b5239ea1cd074c534a96b5212f5d4ae5945d712d0cc2a5d2660c4c47803a55128ee5feebad9a7ed74d17dbd7bc6f2a9b9624ff16ad711d845d7b36feef2832281a5591bd2c4af672a31d21b2e8233a2daa7cbcd64b6eca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fece002b81cb28144651731f9170531cfed575738468ce6dea785b7f442f7c7d1be464adb61aa00c1cf857bbbc70058918a2c9ea05c21071c2a8b8dc5d945df16f85d5dda58f716cc032151a4e100821e9346a143143a687a97e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141298db5dd27237badc078adf7a635a88675a344120d5e613e1d852e11d4e032be042d8b937f71f574a9f471aaaa717f933943ddbb868cf44452b86a06a4b3e8130f7a3004ceccd7447ecbc5318e2966f976e67e57946ef94f827b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1602230d3ec44d97526a0c5e878074bf41aff5642978b54a5486d8d59da3d7ab2a7d4e79a36ecf6bc49c9bf63aa0b2665a00b2ba09bfb6d55e9ea34af6560c67508e52edffbc904dbd445347d4214c99e796c5c5ae1e2e1ac6245d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7ad5fb2b109f746de619cbb77e54d0fee028dff7061d5dcd8785426f37e5ba554ba9fbe5b859d298035427ed3664200616d58de4d2e1b54790fb7250c48585f25b661ffda476c459bc3d5ee4a22f09dce24b6526674779640021c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184daaf32d127d9403b618e0c1ab5949aa64f10bc579c4aee2c9f20cd8596d39a8855c4e0e3655c3626e03e42275dbe350a56084b8d5b2c1984dbb832a589d6c745aa1aabae7a2873f3be0e9924d09cbf916522c3b8659c494651ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h944de7fb399f8003253ded8205180ae26ff230812eca735541f73a4151c852f4d550c9e9266fba8f63e085d5fdce858d785560a38b122510335a1e92d4fe8828d1a9a5823037a52f4454b818a6c198ae9078aad368316548a2e5e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fc48731d38b32365cf3666592dab5c6b9111296b1892f9c43891f85b3cecf8a4df52c3c027757ec9703d3d15b8724fe532040ec2e20338a608a01e3cd0b316a2bca6959c6ce017888c8e0f1384811cf2aa18c7b889dc82c6e2ce2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6283149e86e7978021e6d5c8a8a41f551bb5d583395cd39a6495e4b6027d5a115fb41fedfc64677104cc5b9b1d390bcf57262a7af7d8a68a3278a237d8eaba93f8abbd70c33231c9e2706a5d6ccd550cd9dbbd6bc38aead6744c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7dd110562842e8aaf0345e4c23d3ac1ccfbe20933aa5ebd5e327f3dc242893d931b51c5b6dbcd280eca7bd35ab19eda43cb8e135df04d35fe739da09d12d86bfd54d41d08848d3412821454896fe27f26c2f969657a17d856c756;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91fe4e3fdf3eee37069cd078ffc4cbbbe348a08476bcd9d070c8422d1500fa809ee484594de1968d871d363f543893c316253ea91adbe5b9e0c4f2d9397dcd4b2348690d506086760df022016e001e9a7d5ca4d23066470a5e24a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a1e94429b5a19fa9bc43aa56e9bd275b74c75c75056ff93e4c0b9a2786d810d1b050a9b7b433a9153788fe9603e857dd30c99f323d04d2101b7ac80d5ba5070c37ee0030035fe5bf7c93f277e835609abdab56c9f89ca9c9f859e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c9278ed1239ab854bb90b871ae737551954acc1aa54c42a801931a6fca1779c2f2080a366027181240db7e098b70dbb89c466874f195d9391226d9b86e4b2f6778b2a9386e442bea58149e8490f13f5cd13c5469599b6209b9122;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a23ef48f1bdbca8d1f983216a13d42006abdd97163af3ab53fab0660fb8b8eb551b3f1a78f31432ef38e7e57686ebea3503876c95e90bdc8a89ed4eb62aa5ad8b47f6af3f84052c5992b0f688a40f3ac1d18601be94ca633cd5d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c078ad3921d8782454dcf117083b331694d5cbf45efbd63933b9e1a0030c145768e15ccf8dd4e664d392342e3ef943ca9521305a4af68a68ba5c3a0619c6f26c0c5332f21f26e7b46b33bbe42e408a0fdec9d87c016604728211b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf86484c7f908c90d591428ea098d33315c0eb765880ada5c3b610aff687befe47bbc694bff3bb606caaf2f2648090e183e832c024f52827b254447b4922930aa0f6d357c385b2035b2529fb496e513e23594fe51624ecee7b8cddf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6b4476387324b22786b73c3864b1faf1c78cf3e766377b9605097c76e5b17e4c50b6a21cd1b4813c41ffc1927d156d0bf94ffb773bdeeb3e49151195026e04c4de5fd8173c8273c4317f9ff94030f2d385834fd5a6218981b26bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34677c4c0565fe81976a8bbe33089de2ebfe55bc0779ea5ceb6d20b5a3cf3e784c1c9b2a4882cd29375cf92266b4615ba46da6e4db09541b5f8053871cbb59594fc5001793acbb9412165b6b9ed279fd7c53a40b41cc916585d078;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c348316dc405c6563ac3cbb6d75ee4f26bd109ae37b2eaeec3adf8eb56550ec375c0ab1e5a4952c750ee582b8979961e631de8d429ef013aa4cd4ba9c849b93bd7837d62aa01b497bf5c262626f2642405ea2bf64c1407f9359335;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189e709adab06ef7427986385ad103ccbcfe24275cef9be1d98258d9b46a5819403b86edd42f306832d6750dbd62e92326e7c05eab29ff48e63f1b335a9f9e48a8c35149065cee7916f98b8565970f5092edf4778e916c3eab946db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1559aa38b645925b53f2b340235c915a4ead49af1be6f9a68a3594bbd09f304cf51f6db61763c77440928d2a9480fcf3a57fb2efccb925afb69c52d0be03570ad2c81055208770153cc970e9bb3fca6414097b50262b76b217af9d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12adc670dd9b67e5dd06860081bb4dfb0c83a6481a3ae06325469dcb073092dd262cc9c18472cea3218859c9e744c2cc6955c5ee716b7df99d4b1ab0a2014c573440e5ede2ba5ba7d4957e17c0b73ba02b3c2713648c72ea4cf8d31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1383d9b0a57c1a68b5b777ab3dcc87de62ca91f1203eda1d62f584c5790df793e43ac9fc1a5ca45c4572f22a069cd3e7a444d280ec5a80d28295ce2c415e20ac509ea347ef607a7749410311064980ba32a711ba75a91370bf7bdac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1631cf7c79fb18dba5c9882e594e6fc24485c63160b2534b1d77832ed25f44d98bbd13e3e3d25e55daada9f554a830fa17ef00cf9a981bf59a35a21bdf92409ee4885588e197fa42c60c925c1ebea3cd99f05cd023b2dc10e6faab9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135226334e43021707884eb03d3f7b214cdf97f1f2e9f7c1c10eb4d4cfc43883d25256283180d15de44a09dcf951ebbd5529d2128d9acefb6c47b1289e6280009561a8de299ba1f431e1ac27e2450ef0cfdbdc2dcc66ca8202d8396;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a624d1cdbf1b12c78d2af7afb56a879eb182194e85c5475c1bb1a685e323fb31aa7aabca07b387027484cea9c7a83b490d7ca3da5477ba1af05f740eca506af56a0e536879440ac98e582663092473ca6e10c4a8bfd4224a9d406;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f710299148cc0c4b836d8cd491436c550cded3127537ef64cf7baf7d1999f9cec29e4ff77e15a7d5282d1d7ad2c05b8247e2bb315366fd8c294faaccdd56f77680002e48c151c4e510fbbcaea50a608085d18248d85d2cc9222e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e2ae67d3da29d6b0dd7f7a41ee7ae9edd96f6787a09d93154804edb65e2d5fef271c9d3b4c248c8e43fbc79556a05e5e91e5f1d22423964884790e3ff1f6081a4c7a5244c050ded3c08d98b968cfb141ecd530cf8e4779f2660bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha95785229ba9a4842064a646e73f9bfc0a4b587f2a0d293ed079189b307daa06545219572dba6bba4fe1f1b4d6ac71a53e7595a29117a84eac73e7d48931846363f94c3c1c1ceb7480e2c9adc72031ae35ee8b9ca71336711f7c99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde86d7b267f8fa7895b59e4f64f68222fbc55cd8af211399633ac480de9d5b27ee423261e1636afbea25bca878b58066d5b0dbf11271119f2bb245ef6d8b19b4e97d9fd19782ec77f779184f744dde416014b1bb33eaa29cce80a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h415f2e561ff710bc2455333ef04d0e4781c89ba2b4d9baf5d7e6cf6a722394562af7a7ffa78c1ce71448b879bf6f2b1d248dfd02634df2073fec5605348d24e29473bb268ef07e045c7ee2021e1f80b865fec6fd4fde84632e91f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h971dc8643ef7a23d10eee8d260194bd1fc9bf1aaf42542f426918c76b5a66a9ce53a0e71196d205c9b8b1ba72ba2a467d0122d2775206bef951ee35c48ff1e754e3c9ad2fecbd5f57daeb876d22da7c7c9248e28bbf44f4dd13e9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b8d89d3a499fb48da473378d6545d5618cda622f3002258c5f3ca5d59f450108ec4c23720f0a46b0203c900d09a8876dfaa3ab4ba44319efba56d8e50c4ceef26e7ef8b1f29ae6b24dac93928fa5d6d2f0fb4156d8d3bc6049e58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd71361a66d4642a429765d4a7bf226b39ea65f4bfb6031b8e4240e1de239a446988766a3bec024b27d8a3a32e9214413746437ef626c260a0e1d576f8024474fbd7b25203b3de1fbc2c171843b624384279d30e0bcced04412c7f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5581aedf97d81c1ac7be3a9a071e9ef36e3582abf9a77b864eccae96e0788c5f7ee3a331b06d8274b24f201f40a8d122459cc4ddd40103def103bd107d12993fe1162106271dd320d6ceeaf948dbe87673928115840b97aacd7e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cd90943e2d530091d6acb9a273dc42af54a6aab078fbe45413eac933873f4122e523006ea7245060806e31122a3e210f044dae574cfac02cbbb1207fb58d2dced52f1e05f48f59a9071c596337f7ef756a7a750e385371b9c34d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ffb92069baa616ed6b267f5936668faaf12765eabfbb92ed98b3980eea771d56b6f27d0771a64de4e22f88f12136165d8d10a180f299af9d28d4974d9524f68f1a98ee2be1ae235b393cd2c9dc68ad7788308749ef4d9efe13359;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf40b71f0c340a6728c0b44dff8dad56961b0970ab4b13a6cd6019d22d2bf616dd6df6000525c729f8a1dc9f689926032de43a66552582499b2342ca000c655751857c0a5feafcb5ca603e8faf0c47352854dfebc49ee63ff15364;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166dc58f8b5da93ba944a14bfe16396fc5a4e5a3e1e88c50c176b16aff7d2c1a833ffcf7c0be1f30ef35142fd364a28d3c02a2260d609db183e53d1069646aa2bd54f48e6c2d6fb0dcef76490fe4fa1fc08b933a298bff561332a94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h717b2e10f59317a6c96cc2d572b7be32fe0641cb4aac59ad6c0cca28ef4e5e3452a9076e07cb4a6a097decf2384904e8849154cddbbb9bd849c9b8c857287815bf11b051d28d20e12bfc0e51e19b3066d85c3e4980e114c1603cd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45af331ddd104c15c95b2b30593027d0c86a19b523360fecc69ff44a3e0aa4d0da7fbab0597d84b7f6f767e362318032b9e9351d3c2d1cd8cb2b34be391cb07661a7372fc54cf26b5b67e6bb23ac65df8adb1176cd58e0b6fcfa14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fa79d12ff8396c99e8cdae6031c92bfe2cd9c837d536e6a9430e860db8b9fb078751f17b4736cb61b5675ccb6fe7cc20a08ae5b77f91a87e480b1b84fe7d84c01d55e5eb8d95ed60136f225eb30bc8229f1654bafa3b368db6f16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195cd716f0a96a32f1b1b88f03cc521bd1d44719b280a96d7ba34774c7484b9ad59975d2fb83fa0d64e7da68e5ea93bb97f43ead6e6776c3f0ab403fa3ddd53904312b1978bbca9d03beaba3374af2326a2ecb116f5faa07684dddb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a59b0ae53632580447a5d36154e5f61b638c3b7dd56c8191b4b97963d5d63cf1beacfea456661620aa635bcd80094dd2de459cd8c574b687cb83aefed9301faa71f462cf273506070a612b4e33a03a79dcf8a1ac47fc0113ca32a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101918b8f7cf91ddf2dcecda42f611ed104e5dd0b54299a3afed2544d0ed806a7316832962d0aa6b139cf692108e4c70fb18ec25845e58d9e2900900c18ea9a6d72998fcef1899e9efad17597168ae767461cbe66da15170b19d902;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12213ef78ad424515925b441db0086c6f4c72efe20d616c581c5f92c966957b71155b21203253cf0e3f969317dc1d918e0df9160118323d91b0596f44f22fa38fe977d247acd665af3ed78c74095c1a483e62c4f2e51832c086228d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7216d481265eacbf7d74358ed05f77c3397577080c58116963c6969345d43f42a2f25a7a9fc39880a9f9255412d471f4b9bd8dcbecfd8d552d32326fc2d4df425cd209715df9a3982a67331240b8d676f51b151bfa182b60f08aa5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heebad17bf13f7cbe7cda92f633efa3789b538a7a58fee9fac2acfe35842721798b720c31e709516a8690444b23b777fbfc17c15d8ada68acb2fa2c3b0d3bf9514167491bbc6174ce5297f20fc5ee6016c22466d92f283b6115691b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2f277cb8a5d6b45699574cdb260b46b2472630065f194699ef8da0363a9c5756c45ff50c50a970e5e59b04ac17eb995bc3d8a6d2e2dbe5c1ce564274ed6b82cf8542515ffda62392ce150934ff29e66b21291c78ba09be811b70f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1955ae6db8871363f1f73fe6fe5954ff99b5a725bc54f641f28f0f0903fe17897d37dd11df0600ba9fcef5ed8da27718ad72e008ef083a85987f878cf257b20bd3618d7ece1e026b118eb1c1d0301e326b7929214c4fe6f3fd909a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0e1e4f84cbb84e5acfeecee9204b9930a961417db72a539d7d0c6b502f7000aab804f5e64f81c9a6da8ccb66823e0bbd87a213320a16b16484d5b5ab0fbe81939c2227bf534c59b7894bb8bc3bd16d708b8128137e7c7e46af112;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e108a334bec872ed4f80b736da09f048192dc137a43f10962e50fcf7e5b79cc0baa47d4f4b0aa2e3d26517c5cd513b45b30b714e443dbef510605838687f671cc7651905863f777442fdd6bfb379770c062f3450bad92170b53c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a2c808e5182f685db0f003dd80127dd3454f569a53dd906c7e900ef4054971fbe79c41eb3b8150b2a42bba7d95e9499f90664ea6bc437bffbc077173a0c57fa8f1f2cd676fe7f63a6e10342b2999d33af3b6b7eb98439bf0bb156;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdacfa074f039e0e192cf66b973e02651ec8285a7e68cec416068825b4624c1c359ee409e21e8938e21e82eabddc345c4d20102c007fa8d50435bcc95b6d37c9e04f6d89fc9ed341761c4ca8d9fd48bc0f26e3d532e4c801f8e571c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc5f91dcc65de874dcf64fdf6c41da6b6720b43d7ee0b33c6b6dd560dc664515ff9dd176be516ef1b9a3277c5408c1246522562819f7395982c9294e24c2a087c7baaf30f5cc251e1a7598f21df5f64fbeb7e3cfb3e96e0e6b65ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae135faed78dd4f39f16a5032fc80ca5a6e9aa354c81b17f2ab0bf3d8828b8a695a8bd67a03bd28abd1fee476a6553f1247e5b090962308643ee4d601392fcefde98f41e69909e648dac26a7730ca5c7ef81d0b7737484d634b330;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d259562e29ea4641a3fee0b8799278acd379918eee0edc44a6ab14cecb50d98e1129f8c690421fb099fe2650fd3e55f183cef7a39a19c112317d3bf5d1f03c13f22ed6fa4e1852f7b0a228fb421387992b7e5f3bb9e10028473b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5f9533710fc4f4b3716127b0282658fc2bd17ecff3de021e6dd21028a2c75cfe3a9535632bbac31d8a07d8ad784305a79818bc539dcc69e39d9b3d04d684f96e032950f7cec1bd6937eda335d15fa5c558545639b9df7ac23b3c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f2dc718df5e588f3b9faf6d66ae812f09ae8c1bf3686c86fc73151b1cacbe0aca9a3c84eeae320f1d3ec13ae62f172a721f7fd9298a1994b8698b2ede723ba72a4c55f75e292cf98a2012d6f965d81bf69c81327b5b64203a4d5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dad11275a7296839cc0abcd57b91f2556efcfdb6dc8d3919c80af3e954d2b98cc66ce060e289046a695457765785b87936086022c260a937431f7ec0fa17a43d5d6f4fbd966bd8c4bb572cc3d479f3466af54fdfa5fe8f007c34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29c6eb69a5375d41fdec8c398f74b9c5c0677c81c26e660ae49993d566ec36b56caf5b192d0c5d559343ddb44af793464754e86a627dfd5aaf9e386095c9cc4d355cd0a58712ffdbd8c26af24dcb635ab6fa2a126473c2b17d79cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c0c36dcd1364bae03ac57ae9b219732ecd0c89304f0481f06e7e5fd6d45667d996c9c5fb8c638ab62103e6cebf88c646e73de1fbada31fda469ab7e9bbc91084c7674512d6e28611ab98c9f6934dac0cac48ea149e4beadd2825a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8d365f3fdaf3148ecd627fbc1a7b3b572d7c7736a88bf9e7609bf5c87d2166583bd1a373c74962553eae622e0d6ea08a593015a03bee7e47f98ac2a2771edbc301dfdcb6fbfde8cc6f55a02a8dfda83029d822c8e7c55ef22aa00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4db77a96d97394cfe129dfd579b77b993eda52f25504839b97661b7061e0944df1171f28849ec50ed8724d6e43d3a08045d15c4ced1ea10d803f3b70d0771d82452a433775553fa60ab4f53fc70dbb98cf871bc43bef880706be8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h523f4a022b8c6c91d6071e8595b0df7d58040aafc9a1d428dfa7aa7c865afa2209ca3c5ec8961c234c189d7ca1d7611d43accceaae17672590da29cb6f4e1d34b4b91b08fe59011112e1571494c365056a4149b118b9a295e6d2ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c68cab937741d0fd5bb5f4cc5299d983fbb141b5dfa4525ef88da1e426cb117945c4896b7e447050d3a6d67ee73ac3ed60644e763ab0eb0c1264b33a39edafd025ee9346590b3d89306e5e5672b94e19af35b3aff8d4b77f9dc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha63b45d5540c93421ec613f68bd0dc4fb1abbff2c0a385ff599408c70e2f2f64007f91f94088cd2a36b1c6b49c591660e7afb43f5d36724f4dbca61e42d77ba529dc01b81bede039453073f6b8311ea3a0ef3f616058562b42a81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2e0e989d16e53e224e62734b17ed019e7ea7243896710630c5f15c7e654beb2f954ab7676021b7f5e1ad703d7ecc0212b44a58eae82efdaf55123313d1d3bca71dd6e7c4a0110dc288edcbe37d8ae45130d0ba3e534fada7ad97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17eb8c98cdce57347ec2003812610b1024a4b272695c7b58a7bbca6d21fdfaabee4bd2bdfa9986a678f508f9df5b0a5145050d07d9fec0fc8e40f096b3b96d74d47d8fae73ae4e0cb18e8f065d2ac27101bb588f2fac9f2a11177fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cef07b49ca67b5dfd9bd42f469c9d882ef43a04c0ee2b35e23dca93d8ba69b72da83cbfc2d94d8f2394bb1d143d83af54533a16e1e4aa263551bfac76ba7c39c8ba98a439b142b41ec38353c3b518577deabfa5a1211a8bad00d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67a3858dd07e80e7b02b0661085443f9e36dd9757a4956024d5e38f8026d087631856d099494bbb19e30a049213f7ae5940c0c239f23d3ce6eef07d5dfedd405c03664fdb149edd42dc641074e099bdc97def6af53acd372fac100;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192823b5353c00fb59d378d9b685951c2712db9c868e2138d680d6f56cddac7a99a878a8cbbeb48ee4524a04289ef716387ced10be06f412147d314236f43267c435799321f9b46717d93ce2292be6f2c6c62ab9efb15b53361f03c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1029c15de9bcff6e538dab80af6abe2e4fbe39b120f34ecc72d890be97fc7a394b3697fbc4b3a9c589dc6f45098fb5b338711bc365f37d1d8499aed018e8830d6875283a308df0eadd2c7621174c03ed038ef939b24d055c34f2f37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1114ebe3c3a61d54bbb0930e4ee7c518f4def1936a9c055745ed4e4ba0ce69f839f2c6d11c107324640f361a77f5e4967670b9ba2a924588e53d39733258010dbea6c1d43c04643ceff33db9437f24ed19e20ad5343c92b1fe5a642;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c425d748f95fcc6a35db6ca7f4071e9028ad302d4dc1fbcbc06f3cfb4af4334746a34d1dd44add799745cd77cca227420b87450cd10902a6bab4b0218e74aa54c16837107a754a6eceea022ce1d9d273badfa1d8492f9fb84f2be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha80ee1512d93c307e446b3662742d8eeb37cf9e12a548d73be7af2cc4c07617b100223ab1ad0978c6489eaef76f1d79bc52338258e4cf817beada74627a7a6831a8e7fb63585e8e5167671e44997203fe673fb10d8b428bd423265;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3aa0dd01d72637212aed248bc440fad0281a185b94747e23c15e2fbc61b5f7e711bd6cf45f496585fd3e5ad26939083b0f477272ac75cdd2b829addff3b7a24f14b7cc8a5583b7a0938cfa605afa347dece49480ca70d25778e905;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1997dffa7a6488bc796bb50237f1775d1580af91008d5082c9d9ccf46d2a8dde741212c0f6c4e640c0cb7d4c750e9c45a82c743188d8188170e28122d0bf434f7cf73974527d0c3247c0d5afc7114e5455203d69bcd1034131e3d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9386bf0882b7ab021be181718b998dba74a2aba5c78d7988bbaa182c52b4274288c0087c82d49fb2eff035336fd928f9c7d93cf459ef73db251f42d777f0b059263eba4bf57abf07ba91730c5219a888852a12933c9cb5d6541e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4cac319f752714c2628f7de2427ecae1b5fa9fd36c1f0708172dbd8a9156b4bef3d67f7b7d2d1d5e7db9018ee7d45eafab51a487368968d79b98b4f1981f1c6502ea70cfabe14210d8a2355a1944a2c06afabfd439534aa8658524;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc580f1fbd828cc79d24bfdfcf147d8c501c8af0359d4cecb10f081775db6c18ef39ddc08c9692589aa3d506468b0ea95c0468fcb45e398e557a05b72c786de7051690290d35076cf2301d1fea1df3aecf932b5252a3e3ff826f49a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8cfba7da2ce93628aaa498e4b9f9282212fd0475c0671faac4ac2af5421c538938515d0703126038fe73323fefb17f38e7bcaf9934983df407fd37843d6a9fb19461effc96034a9e09be8e7765ec711703337a080319c1563579dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha19345e29b4a91219b935fccd15b5083504c6339e8c0dd167b35ccca0b52a4293938cbe438cb10201efeeb0f3dd017986a76fb6dddea14a03da202847456111215f675104353392e89e8d83035847661a90983b3f2afb0c42625cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f712c22ebfe5324f65dae95ed2edee04b8c2e08b974ef0bc3eabafe796b27fd11056217a5654a815cc768e8cc0bcfe8d9f81c8cf00bac0ab7b536cb28abb9ebfbd38993ed9797d20b915d50c9c78d1dc02533b162487dc7b8194fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbfad91b69ecf87b2272c8820cf3648f25a1e6ad142a32b0b31156a0cf9058759b0a5488c21e7e825c21562ef03d47fbd624d9304bca415a403e1a447a7d60343187803e179b9b04f1202424ba5482d087efd101467e2b7b12e6434;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19246f169c57543469ddd522fe99816333c3c1f82653376a0bb37db7e8df139e61fb61de753c0487f86094558227777ebe614a56085f89f9ae6e1d6277d694db2e9d41dbc6ec9f28bfae25bbabaf9ca69c3f66253458ae9af8ffcaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10df4e8b0beef37dbceecc30f2112d267d8d28dbae14a95571f74d9d2e1bfeeed4c05e332318828e13fef6dd476d468f90909e5041b794bac2761bd91ea6753c3882e55c8482b64eff82a8d664e5d5115dc6c9faaec442529a43b7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a38fe957674aa1f92ce4afd11b133011bf7e18b583e4bcd83982dfc449b87deae29598b7adc85645ae38652082b4bd6959d6ef06cf2b53312d1c74e1a9c76ed79e235d4a55241dffa6fd9f59814be6079d8b2c2e832268240a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa830bbf8fd508cf0f66ff50101f7324b728c8e5b15b02ec983cddb0008cf36f2659723406b106b2631a1ffeac16448141dcc37ebc730cf9d754b4847e6c4f6d23829b3c2174a4f419c91012b91b2aa771993cb297fc611f8d8288;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169a6b844005d7f5e188b7bf62db8df8df60ab641f372dbce43fe2b49931faf00d0520ff2ff4f3a9a5cab3ea790df571d9b07780c4f9c90d9d64025c4a145b2202feab598bb4da07bb1d794a652e2a73468d19caf24da39de9e09d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb9ec161c78e97a903a209510999b8f65b3bc79b5b7396cb669e3437d1c0e4e301a4bbd97d4d802b3a5182823aeb7efe815f87bc2132cd8c35fb09c4c8932c54dfa33c1a176e124c949130ee4bba8fd2ee7986c44d57a11c8f7bb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8229794fb3eadcadc2f4ea885d7831809ca9e1245cdda1fac03fd6333e5dc35f30b32cf9ec1eddc95f093fea2a31d4c42f9baa6f4907263a2e4639b9b701fe39bf99f3a2494ceeca02d15d99d55ec0dc93dc67f47d79f1e37ab5c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17062138e0dec8f87ca90872f6e2205bf514942d68935a21acb1da66e8c5bba8a7fd8750beac504c3dd4b9f088e4d8d431d35f195d97e1fa3f017e308f9ba65b36b958ac6a56bfe1223d30f9e2fb34039a05801199e899dc9dac7c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12782dadd98c71e381a44fcca3079838ad5564faf913e28349d96ce72b626e02be5dcbb3ec7112b1bc30f197bde0e7efd24cd99567779db171a543e7112ac5a690850382dee12016b4142c386a1790c40b07118caa039e80450fefb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1650786e6dd041973b78df60244a3df467507bbe0704615b5dbd5c854d4c1938901492487e36c1487e7c3f9b50bd12591fffe5bc8ddc2b48f38c0b92be0da3ede04d8349b44c47c4ded3a5c252329e400eb31e6c2075187b106372f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6d62e3dd55ac7433b4399b75487925569fc574d2a9a8bf67aa9f156e03ab3ea8258b4a8fd1a0944230771feed521b901ad56ac70604cc4d9a4e0e9369d8b968e797f46ac8cf447930b4718ddbb55b157bca55c715d1b9cd551ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fd5f3041cef73af5c1406c84b73b78a7c071318b5d46606274f99d386f02b385ce087168b4188b578f6776fe627096b3de1c39c793ea68bc8715a185aea3f86c4fa41b24cfd0ad13d117530f1f79d631c58da71beefaa038a92f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51d5fcab70fba700c57ceef909687b4f86989c3d5a5c773d02b316ab868c3b796271bacc91a39c1a01a3fecfbe9c8da93a82542eecb48f921cfd4c8492b2e50f56182347fcef9ba52237a2d9cbd92b7ca730ae17ad1bc38930f715;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc46240d6e026c5ef411cb758c1e421c399e92c33db8357427e26853c00a58e472f21a42ecbc1440dffb8b4517d5265740d7e44eba1dd5b67cb80ed53c44efae54a10342b455726e222ff1892f5f51e0d891b918e306e316cd2544f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169da3417d16b9c4e6adcfb880f21163d9b444973a946752289a44e6cf5d5d2015297f8a0e682b55971e136b061f98f4fa96f63d3d4cd2a57390036bc0168d13140fc7ffc06c7dd36f8cb6ee798edddc6c6862e373f44d3df4f42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f231666e1e1a1e4298660df00adee569087e55c9848ef53a1b98be2614b862afe649b1c1e5d2a223ff8c4f27267e9f153e5f52d89844f85630ff4155ca147b75bc1833df8d3b266c5fc8ff3b1b258e0e2e8ffccc1b456c1e33d5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d0fc0e3570466224552258a3823176b1eaaec625ef1dc9aa45f07df3ee64d9f46c1e497ab47e8758ef4dde2aace9f3632266e6bb1a5d0acdb1f1740e43750938bd48971c930e6b140c0b76d0d46585d34e83689c17b4a4521c5ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17233161548b9f3085c65f2028c64513cef3b5f9d31e82733381a23476ea46a708e9d3baddef80ef454d2eac007a199ebd52c92b5f544b7015721153c342f2585d95e47e716897ed7d504804e0e732ceef2ab87e894df935e2ad3f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157d96ff179ee7bae2532e45fa27b0b6bbfcd2803125ec76d22c5889d43b99b5371d1c44f76dc036b103d9e1ecbc95dbb79ef47f259c1374482e263f7aaa831d443d5ce767414132cd5fbfdf9f7483252dcf8f1a2625c8cfbc4979b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1090d6d352743e7d03e8a4430ec336ba739a167d02efd189d72c8014c26eda07b3be86e352f5c8692520c9b744b80fcfc35115324ed6534b0e48b384fbc4eca9a50105d67736656abb56af880e5b35fc6dd6df505b29eaa7528d79f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64f3cb239050172998760f87da424b20dedc064f225136ea1246ef2ccb74b2b7a38a24fa6c705efd312cd5b22bfe0fbd68548fd0c334f7186cf1184bdc870efa71f218c3e81d70f7000522c0bd6ef31516f7fd9a811f84aa211a1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf013dc578b5d11a4f151cbc0cd2b60a7e05f8b7ef2511fbca41b37686ca91b215fbdd96cbef85a456c729ab0ecc52d2b40281ba0f23f0fd2f5517eedf1658718a2a7e4a20fc706c754a798db3093cd2ee2c470134c9725886d91b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf344ae1a133b9f225ab2d9e45d710ae795433000e83d758379f73bdc2c521d8b0827bbd8c5c9585a8d352368aba777da4c4ad9f05f9b10f3df512168579dd637658c4e905250646ddbc0d3710bb2689261160602b771c4781ba055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9090e2ae94b9fa03fd91e5420b72a5ae9a673cb4b01e00d2fbdeb9a91af5cb57301a3f9e1c2b09b3cff14db42b6d6cc5a59cdad2cc4b5b277a12f1a945730ed2da0d97e0e9ab8db4f94dbb5d446e94e55c88439a45c5f2b2d82af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15392bf31bd9bf59312b773b5c87fc3ebaa4ec15189a282aeee5ff506df2bac1fcd2d2cd29c6c1d8da549c3eaf7bb18bee653c658c9c469aa1c33b790c0aabc9a3de546d288cf47077be7cbf6c079fc05b852859b482c06ecf63e43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195b4f08e66693179cc837c555b91c409ccd4c0d10e6efd12ae51b3a87af766f7ce47b9a4443022d30f4e1ad0d0dce4801036e820a97693674938ee125d6851d26be121b335b391906a5c2f489103f9fda3b7988a35b835c20722f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16443fee3aa1b8e1117780d2f5612e779715044b94517e5d77ff79c31b778c130b0ff39c293b7c76ad531757cb2b89b24c13a8b63b9f59414ed2016a321d7b70ece2e73e8fae91d72b4158a1c81f5f6fdd7a8d5ddf697e691f64569;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d702cf62869056320e840494a4d30b753d06161f9f2539852c934520abf4482dd8fd5575b60e9fba1c82412dfc75c8ad64789e83c18885aa31a475fb774e5458855edcb79f88cf8295bca0674018ca745e27a1cfd431949d935709;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff763d97a74b04842adaa840cc00f7cfd44e66011f5b50493a1cee9886913cd362e8adb009e828f161bd807fd8873bf18f920225b347c57e3c4062775c8332bee7db1e887795e6514f4b967faf7d4883710b45129a7e7e4956a8d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h824d8623635f6d9b80c7f6f852b626523fe8f174e966cf9aa9b045107140f4db7fb7ded1d89cdef5fd6ef746dc2b921e630f27fd78af7fa161f5b32806093d217da4bb2f8b93a9905d0569e67a4642f3b4aecf1dab5dfe1b7ad231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1168d64bc5c0949461ec41bff77af8a3c879556ce8bab87d73784bb1dc01ea68b5d40161ff5d16de6d31d8fcdb57d01dff0ce42724f063ce02d91b6ae8b6e44ed1b7d7f3b4ddcd6dd60c812db732c387af9d1613fae769a3b9b3f91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ded0c97503a7b2fe126e599028c96cb02b2acff97d62d4e82e38c3ff9d4ff7233cb1742d33f789baaeeb8ae42eec39bc143c58738839b93b6810e2bc5ef2649a3be5065f44d19b76804ec8fd34898130515a961fb07c269bffdd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16afdf95ea88415827cfcdb25f14a5fad00a655f3e569f776b23a8c64f5537306252591bf566825fc8cef1f42474d52b406c17d47c0b971dc2f869fdca98ebe063986a2b822e17f731e4f52ec5059aec547d8687cead8e7893f12a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133c61dae2f8ae37a37f276257e543b644cd9302918da9857c64a903c9561a8282ca50358131acca71eb5e9231f57d7ddf6a89c36d3f4bda7535b94f9b32af33daf3e3b83b5bf4976e83e429f731a11fc32aa52dfc23fbeddc475f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0e83ff07b1460299d6b8b5c40f4a70ffdf12fce15c92b2e7788b86288d2eba36f29be23b6a1879c050a7265199ac3531099d63d748534b0d1bec8bfc5f59d88bc1e9f10b8bbfc3c36463bcbe3ba81610aa54e3a1d345afe090b31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c7293d5d607ac069a298c57bbf9250f1175f8a980dbe0a14bd5556262e84681f7e1e06a65b02ee7a32b301e4e7cc2360e9075f1eed476000be62afb93853e892c0142fab05f417417b9e9efa0e02555d4ff8311e3ab3192eb757c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142205895e43388ea0981e3b9a9e65c50c202a3f6dd182b6bb0ac4624fd6cd88a5c222b500283e3f5f96bd91e93ad981540bfd0535d6971dacc224142e0e9028ef1cdaad3bb8026c0c2238414403e64c8f2de6f4a36b95affaa562;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3dabd4ead262f840106d2d15e463a28d3ea9e37dc71c69d3fa32ad37d18987935125d8805ad4fa5cf4664219997e19c1c0541a7979d67b7f90d9dc6e46203779f5fef9e83d31ea7c197cb69f4d78a120b642072ff9d0f3c0311b55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a5645df0aad62973ec714a02b2bfd1c9569d7d2a5ec6f0379c151933a134104220e9537feb271c706555667458414391b250aece0892c6ca216e2a4ad2716c7f6df829a1bfd8941d1118cb22526a2acac6bbf59810a2d4d8f8b94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a1747d4810ac9eeb92c051d979af4ba9bdb46a4d8e39ba360ae7280fb847cc7942e17e1efe6e7f0024c096ed22fa4cd8823f16084ff2b7fe3d804b743aa9abcb6a1f172258939f2632c22fdad4ed5dc9c00ed2f80fb789ffed582;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168feb6b216f041572e20db86e4529dfbcb3c1f5ed0c850d0c22ebaa9d61d1e1570d8d826e85e439cb46773ded2900c32a58b19cbee0ce6e614e4e2ee14e836017093cf8035b7d89a8e10bfd9ff6dc503b830f68b7f905905ae02bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14079dc97d08d72d901ed234b46ab65dc333a466cdc526c376106ac36fd70c4695857741873812ea3d62f4f0d43a76c53a32a30661cbc76fe04cfb7eb5d4bb02f34dc1a8dafda9bac23d7cc7d1a5a50d4a85c6e766a6e25a31e1b53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84114707eadd5861a56ea024dd55bbea2d8f7bcd573a0978aa9bee95e9a11d85094d68709e808eeb4fe22caede5e771d4c1b2276a32f0ddb788dc1e173416438fc42891e8db3f84f3bcc7f881dc5148abd51a9a2acb9528774e7bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d01bc00f962c8cb1a1e394fa7b1db91cffbdedb7b99667719ef59fa46513b10a6d76eb643ef4da6bd37aa07d588433d469a7513139727df5445354d507ed90e846f23e2576af9a766028fd97efebdf31aaa9e8d09fa715a82d4fb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143000a9029f667af8e7105bc9fbb3b816218cef98f85fc5e0f7de711a2277522b7c0fa312851f1257e6b40b67bde6b37ab690d0f5aadd396387056be55a961476f2f471e4dafe0144eeec0e41c8726c3d05982a5e5f95d9fea4d05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc55045318a9ba6d62762cfc8552d8ae719922d0bb973783aec09595a61bcc1112d7255fd344bc69e86d2e05027c7c8541ccd6563be01ed887c45d33a28b270403f76185a3436225eec840cf2cfdfc7c547ec26292bfce323c1122;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d285d34055800be0f99fa06175f1f3ea064c7c4319da33b960aa300e62d2574efc505568635a7d9205a60c830dec9a96d2c3bd728e31a8b379ef6fa9d39b6b6bcdaefbe913bdd0faa964ab1280a508a553d9cc1d4e0fb28a691094;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d25d2732249dcb65b84c244b459f98a3685caa8ac3011dccf39642228b642e270beae7fc2f3a4d65984a417a16da92e3eb502df99e12ae76be5a37a2461f89a2f8a64918a09002c7ca82058c4232c139ed2cb90bb4daa4ffaa504d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad23ec1698b7ac3e2ff9012432ba4ca9253e8505158a00047597140625f7846385aeaa562c155cf65f44c183a61a2d99f03c00e2cb72f1f71ff81eaf3c9e87c81142601f35f3d2f366598e30e1d6051df08712216843488266e213;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17efd5fb8db32ed2dc9f918859913dec3ddc52bbfdb8360fa5cff241eaa998b709e975906e7d3948a397fc77ee4bce794f55f1b55562191a8d2eeb7ee3c31a451e8d4703347f9256e7c85093eb436f47a1c8bd0f58a549a8737378c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1014d066f9ff40c8435991dfecf27096ebc02f7d75e9d9e5a3a871ef6a75a009dca08d8d591d89180a5aba932f68ecefb08a5572410ff5f1733b0404897ee64500aca5aeb60fe52f226e116fa8ba620f3b8239a33bdfcfb696512c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he546a03f5ff5d29d6d79035de55d50e231b2192afe99323eb3769a79d5efbd188ce0455f2576488881e3791212cffe3127301d4ca7c567e4f99540b3ebc887f88cc322bb772f984abc6dbcc9439dbe87a5a20fdc81479fab42ad90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f69947282744d9aca0756eb9c8feaf0ad64450841d15f19f0350500f7872279b601b97ad703861f00141d0f3c216b6e29e6a2402fb597485f95f660dad13849e6435dda18e0cbf5174065d0013ed83255403ba74af9133c0ac646;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h773110e1b22cbfc734a4feb2e8146164c4e3a689ba60cc52f1ea8cbe8f44d493d5ca559989485d5223748def31ebecfe5ba42e7d460a1abbd2988d137a1f988353a8c05a92512a86efa88f82a3275ad3f2e6a88a897d57a173a882;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151459e1f0bd070ba08854ceb63ddc03c318c678ba2d110d3106706d439ccae26c6c67d2c85a8ce96094036708d5b4386bd8f162f6f096738750423ba9f174d0c57c4e21da91034c78840ed335d047d4777ebe1dd7e66d802a738a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf520afd89617983042cea766c5db65c3462443d956173c15454c1cb38123f33a26fa96a6c90f23aa6066dad7acfa1730f220fb0112fa237dc79b704dc1e94120fe59ec8f90fba55637f018e8f2d405ed0385810e6c70074b56f00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10514cf6e560add83302a7c61b817434f50af11eb5105f120d6da940b11d887f1b2c45fb52125859d74fa0ceaca21ae9cbf923d5f0dbcd59eef74320f54bb3af66002d0d7f6f0b822a4963870768ddb072638815ca25ed26ae0d338;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4ce733e7299ab6622ede8008d0b953afb129126abfc84085d49bd08d30e40c45103d56df904f58dcbb1e0520f69fa55b7b8590aa94fce266e4125d7b639bff6674b20f496654ecfe0cfb64ef81eb3a1f891e9c843c796d40e4633;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169796be810239d31191270765ebae17b11853ed35ed348651e8517e4dc6424f06519414cc79df4835edc1f9c51929a8af091898ed9abb4e7c5b37a5a1bc2b374880c588cec53d3bd8909f046c1f6268068ce5cb74503675e8ba009;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aeaf6de1bab0ec374cb2bcb1e2ff00fd09c61c21639bb129f85f1fcc7568c85cf4744439752d5c57fe0b25357a1c0f29ff0d1575517fb10348f7e4254157a032887dfbb5e08a716867a66aa4fc2443d433ebf497a4e3ccdbf6db14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133c26ca192a42e46a941063542f912f1ed86baeb499ce36e72a8a65c07e4fd742a02cac43abc425ef7037f207c0679e161072b1c51b14505885aa4ac17f503200635c4c095d410dd28943ea0c2e0f6a96187214a54e27f3117973a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b5c57169ef50ba644df944f57c7e428ee4385e7dd66088063b7f10ee325b4469d176004fea99299076d53691a82648c784b6a5d378e7e3cdf157ff9128a9519708e4973817ad499ee3c66cdfca433f066b7d2add7ca6850e66640;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eaf61eb55602e54711b3b39af38bdf8613029baa9342f7b0bb83e93700f6747a765a04ba847a6bfadb0b1b2d7975e76ef9fbc1ea33b181ffef92f01c22370c48cb23b6e8f4fdc62e89e2fbb989b73e593397c6fd5ca0bbd4872af1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70154242a7fa1860b836abbadc4e9aaece7c23fb315ec9846e7f834f65c2120f8d1fe2d908c4c4b663805405fe18ba98f1b6d9fb10af0014f8793cd9c71b7c57da1fac3af13b7f46d81027673b72153971f81d340d8633b64a566;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h916eb3fbb9ba676930739ea7b9399d9a76cf2bb427dbeab12ea2e380cfade29decdde4ca426cb1abbebace123779ca770ade77086133dd9f899d5fafd39ba8e0dfadbf73b6f647d8c1b2a8d1aca4c75fbc133195ac91ba26214b3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1385dad32c5e501fadb3444bc53668a193c1dd16ecde909611cfabd21ddd78cced6998b748cf018aeedec4c7dde5de9d99b555f89369750a056a5c0dbb9e14bdd31f8a89331cf2ce20a92543ae3f63ce10c8b2b6c6116f77749a460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86bd785159104cebfd6ab47ff3bfd8f414704f43737a9f04f5455ed43da9df4effc7c928d863559bddc4901789b50422869f099bb5e942e986416afcb1823c2ca6a568500d8551ea7abd00e04ec0b0bb968d2d9fbbc6d82731e3b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf32080f7d2b382b49beaa567810715a60e6a72c9a8ecc1ba52bd5088c9ced7d0f652de6be3fd4df6a112a9db85149e1e63ecb90ecb3b7a3392459cc2c4d6490141ffaad53e48428071a36dc371cb20b17c229c7784a55c4a890d6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e79295a2b7ee73d922cc483b48a65e938e9ccece6ea3e9e39f2b176a8f16edd3aceb05f7fde6a607215a62ae6560298a11e2bb22f35aba0215dcbebc0a94aaf3e8f9e72aaea915c3bc2a497809a9b2091296e8e4a16d8abc6f3a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116a2077b2f5ab1c00c22a48d8914de55e268233a875c15b6b3f24672647bf15964841af909470411b8aaa8844910eca094dfbb655f2fe969856ab80ea4650cefb320634e8e9ef6027974b53e7f6d545d9718d6e5937b0692318c5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb17277602d6b30fc25ad1c78cf42312daab6ffe0b7bb19294fc13fdf52be88d03191509fcb24209a1120d81a7496291e765d30b210355a6f9d7ad8bfce5fa229e9be8c9e084b74085b483db41c2c4874f2428523985e9a3733d69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b487083c722ca95fdb56c3e99ac89023a643a3fe13d658848be22045be80df96868e17f59027c4b029b09a451b4dd7aaf437962897a94aae8dd4d9c06c266adc88b2727329faf1d6dbb8b2a399de0947032018fd0054980453792;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158a132c5d152bbc9579ce4166b5aa5703b36c19c6fe3b3c55731803a7c923e6ee5efedbb4ac7d95e2d058dfb30829ba092cd4b2d982e1e11303926222521cb8accb03b94d06bc646de3bdaceb65b5111d7ba7b59ec65e8b2051cdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd42a78ef5d0af23dc9b38a409cb87a4e3501d7702904b994d88e762e82e7685f7084769cb7705234be2da749d2051001a602ab9cc4b29442e689eeb74c59366997c7c6a83ae4af3b0e9bf98ab11e6047fdfdc49d0f6b823dc06949;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1e4a2b6a02c3e4a820b05e1679817cf5c598c93daad6cb5bc523b3e079fa02b254abd8c4a21516edf708fec5d690eb0f7b4706fdba2bd64c9644d2e314009333056b1221be2237ac8d64baf75cdffba14cd09792705d20249079c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3bfa14552a274508975658f394157e8093885246b5cf271aeb9741e1e27ca3e4d6967fb4b70e0b74f6381d10906587ee4fbdb39b5ee83e551bca9014149d480a0eb91cdc58c47df55445597fdabbea479a1376df3311d4092f265;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7b456fa155d8482c031da5073fa57874745a08ce3eafa647d338f4d2735861daf204628be96558e34beb38f0fdd6ceff1d880dfdee7e5c801c0198800f4a42992e2a2d41170f085a0cb606d8858f71e3dc5ac3ae10f31bc0ffdd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25e4d979b3b1b34903fb43455948fb7315d8a98c215fb87b7158d74e4a1058fc84c4ca3a736d3a343187f8af7b84e606aeb789bf691f788217b225c0e30a089fd9f08314754ef075c11dc85d22407efdea038611f1896dd35b6fbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185688d352cf139f7c5dc1fd5498eed05aa0001e0622546b7bcc2e50412bcb1af503ea47cae6b06c39d26fabdfcb6a25c7ce5c4f81866e772318377a75e500ba32ed27ed30c8dc3c98c8892ab01604a0762d0791c53cb15c074baef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1d7babba2108ffb73b4d233395b80f825086efb2c9bfa6c461e0cb7cf3196203114a63a91f517f698d5d32c8809bde1c6cd4b2b5a6c157f1b133ccdfb369a84f655bfde63f153fdddf10af3663f0e9f6346ad53df1a7d66d5cb63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b79127490d831b0ea821b44db47c75e5d64324c576ccf57989173c29cddeddfd52206fea405552978e247b29d1f342a26b1960208f7af7a6e817d4c4730a4df2bdb7172da8f2b5bc770bb3a806146c8baafea48f12148ea695d8c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd489ab90e22c04528483035f4b14109a5598a93bfdab7d16724ea70bc138d9ea919a8b3757ffbd7235b9ea4e77739f3760d52ff52ed96837e884438edb281e3d2551e2121afe61ed4c6b0b7c041614966a94bfcddb74352083909;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c8b84da74f6aa813772edf71ae74d822cd0660304aa46e5201a8088509155fd307eb99f93dfb376b0384597fddb056469571d71adf1bb702dc2763ffa57cd1472d7e561e03551d167acfbc688eea6e165c4dc82660bf1c50ba7a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6611edc49388616a3f4c758c55909c03232bf6b6865089c7db07cc2b7d5c0006a1a2f5e920c4fd3019f8cc0db5a1661d5daa5d00edf522ffd6a732f6aa4d354a81d11fc630ee6fc9dcb1b01ccd5a771ce45491c202d1804d8c9962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f63f7ed091739c1144073d452b7b5d86bf4aa812705b8fe28bfafc72ea25bbbbe5554410e50e4c82825613550ab6ed0850da154bf63ef28651a1071784c4d0f66cf7afc569da4d47ec76770f3740c937cca011bbf7b904129fc35b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1997d3b8e2476fe9a0cf8facdc681c2c7d3e3d3690c13b6b65625f867127b7397ace9ea52ba47d3610ed120a4a18edfc964443109a62e25e99d4f54b6cb15273fab3ae79727af046da19101421b266cb1e72c5c529ca74f25466edd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha063d188cb6c7d45c91c79cb6fe916b65454a4967ec5fcf0a9707b081ac37fdbd2803dc624f0c13d3933732c9e279a57e74a975903e088cd1f1d3c0e7533b6680a2f97e02533d7b0d69fe3ae6eb5b9af5c5cceec89cfbe0dde0823;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h952da56db8840c82615cfd7753853eda9ce79c1594616b016455226c0ea05eeb214fe3856e43ee30fa06ae0c9252a3f805c2bf9c4937e2aca7bb5b8ffadcb428ec81d0441c2617137be1085fa8341234a779d8883ef3b2bd31bcfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7f12b3eb30ce5b6c9a4ccc5851547e2d83e5c5f59eba9122120fcffe313be732cb79983fa83aede0c651e4e7f5703143f43f8267ffed54aa2439e492e4c712c99a60175ec5a30096dd1868344357a34203d88faa8e5cc113a6b48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbe989d565179cf3975ac94a87dd84d154819f58eb42ead92dc4c217d441639929bb8d2ec7ff5f8a4b9c1e23ee5ca432f625d748b0db94baf5becab09040249e39d844b34e3fb51cb273bb469bde605f9ac09c61ce90f35a30bd657;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16318de0565c5d866d4d910ab90794ac57a2df91b299fd5b1ab2ce71f0110ff0961312dadc50f22b511f91d4f711f51ed98f7e17602affbf7b63c206373471025d853c49084adfe23398ec6879351b6613af89eb74f25bb29f15399;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf60eda384b456b04a0c31203ee378a8690fc6e9e6da306ea99517eedbbfed784d1dcf36becdf34341c60cc80aff1ccdf1e713343b093edc50ce6d5baa308750c5490a6d00901a54710f0f5c7b3a647ae0429497b5ce722e0b1492a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99ecd36632f29ab6c347176d80a99c9a36af436c25090dfe6af5af366d079451c9741f7a2c07fccdd7b4f39821ec35515306b784fcbc9dd028c290e6c2be2825f8a10dfb8eef0dc5723712caab045ade382ee144439e4ff7339f97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19916881de45f5b37917af352be58da59557d6ade14c8175c1fd64fac7b81fc3e77586d36cd9ff0769282867a3c966ebac4eb72a1a2444f19af58ca7cdb900f726850c37ce4ea203aec8070d1ff3c54151e28cb97d94d1d2b35c0e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb78dfacd36db7109405c512689025dd240f225102917b26e983edbf70db15cf486b5d8d0d068d10e64205f25d7c6b04798b43f82ccc23d78efea5525896710789b9c4cd0d8e99faea91ab6cffa58b3a1e6c9cdfacec82f59aa998;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a45e60777c9855d40b8d52d3e91aac5b83bf3dfbc2bd6826faa73f0c4d34ee99e1ed174d3e486568050866e66f097ce221302b6a6af5617adf007eac4f200fdcfb1890dc7f93c97739f87211724481823bc06787f2c4953e6aff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a7a8d7287ac056af6226e88f88f47af66f32f4b6d99f27ad0915ccf66e69582c4670576f3639ef6ac67490e4b1d0e8d463fc840152d5911d761fa5b17ebf4ddf39d6cc7b30d5a27a5f6e39524d451f721ed1dddbf59c43d589c5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f9fec061d823cc3d39f21645b4081815052c09b75451307cf8a3f4713565e0403665dc7f73112850f6666a06a8834931082b1d1d19cb10fae08c39dc1dfbbc1e4fd1984aa634e9a014a240314cc2158c864b8be62d03b9500231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55d3aa98312cf987232550c097c820989d68951a2dc3d06960b770606094e0789378715964165fd583da81ade4015ac5ca524cf8cc50a7cf5004bcf1c49f58592ff27165b89412ffad6d5805f9236f365d1a9afac86ebe840bc2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd2a4ab49559d2e274c87b4beb2e8a4a057e1ff14be5c2ecc7c0064f9063ff77403a4632120b912fcefdeb37c8b26f5aed44ac3af4987f671a70e5af64ef4c19a415fecd13e9f21ec657b3c879e5ec093b11bb6aade704b135d6fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baa8e7deb6e5665a2aac86efc9253013e7365066c4e9020d791c0a2d75e8195aa2a340210d1def3ab40f3b414c0d4bd26dad65e4ccae9a27b499961a3ce733dffc6dbb9918b5f2b76ebe386308a780efde119e50e23d203a1e4340;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8b79cc2cf55907b65ba00f718527fdd02f81e7735976f52625ccd8b4483d2f3615c78ac6c332214a8ea3d1cb0f9a8455f66e2e225f46b79f60757cd8b1ea823ebc8b791340de820f44612c79e9ce93b13b8e890b33cfdf43f7390;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7323a13027a6d4cd6e9d81605f4c0c6d5379ae65032323fd052570edd5d7f724115b267ec5df97a13eded0f1b18ebf9cc008e117712db48acbf19dca4412bf6b1b5fac4696cf72d8a05a2fcdf0e2e0d224f9fdcc3c7721a8937dc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189962d218a2f200454ff050a15e28f37ac5bed6558633d99c9bae1364faf7f5142748beb3482927f6a82f314227a376690e9c2aa5c028e0b47bb389b1191cf5e372eb407084fd12d3eb80a5938b92db450d4efb6899619a4bb5ca8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37ecf5fd3f2eb773d156a0517c1c10a879e74c027231c8ad870866246dc550903bd77ec3a2542749de51dbae33bf8a34961a7648c3831c425c89f2d52b191c4a6bd81302e158c1f3170fd370aa8be0a388784a16eeabeab0d1120d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32118d9f179ee13d9d490f7969fd971670d01b121d98e6138fbca21f14317a17095d3849e1d35455e953117c7b606d5c967d45a6ecb839d3150d6497094cbbf019a7413e446f273cbf5523f87552e52d4a1b29810ba858f1ef7437;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c589381a937b18249b79240812f1216ba277150b76d33d39506933e57b810b2f5e43d20ab687ecd30529454d205e62d34fe89989b9be4b9bba2aca73a0351034e1b6f456dd76fde858bbe16b3845de7438f94f0b98912defde7e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h445cb0e4b9e720a42dce6e5bfc5dbd5a5e628c3dd1924533fafe58cbe9461e943ee91f970e0d89ca3ddb0280b0e0fd4d709690063a63b3c2b1680dc42258736e4c6a768b9ff29c90567256838ed2f59df716113128bee337f50de1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had076b3eefd41874f117cc312189e186cd84a9059d650f97e720191b1f43101e1a7361c831d932b8d89f8a69766498733fe8e228d18ce49ccffcf0efb47f872e3be04a17949cbed1bc4c1d5fca46f84e351ff10f89a58618032b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h539bbce11900287124d9063e85e6314dafe73c44c95a8a53b6fdb5ad26c77b7460974528a48a22760cf9f2fa9e67d892f60cadafbe7ca1b6443d708b0a6a4daf4cddd70f2b9d5e2a6e9d5d3d194a1d3fab04a5a8a8dbdb5b6cbbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbb11a98bae7f1216a7c8b2dc7a7d08fc2dd48dc4621dcf3c82e63f2cbacc8f67428d6dcc445b90710fbd2dc4b84676111f7da86a10581d998b2fbb6d6334d3ed3646a1efa1c31a600ff136e0fde6fcf261a0cde32b606aadbf3e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b731d764160c9a46b2ea260ab6dd002a29bb4a43e07ee8a211f81df55f04d1e1d30f3c211d8ace5dac159861c9676dd41434bf00d67cd390f829968365f1ab41eb2f25ac9d96ab81293c50ede100ce3cdcd5af5cd2c17313bbe86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fbfcdfe9a54e060c6a12c4effc7b343bcb893251ffca82246bdab3935f0d1700edbbf667f0bb807188520381fcab6e7884009cbf291bae3d151a3857d30630ff6ff37e2922871d979a5879ba3c281031808d107bba2b1fb4440d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1106ee05d69411cc2aaa88eb30a41d5c45c4a5d5411589b0d3e7f85ed17389a39e617b057c33b89016c4e0d3018733870e29456ab28633a88cd6939a8ba0506ed2fee23e513817ffd857c5efc24ecd6bd69f9de49563574a1c559d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff2e0a2d43ef72819e2f757da77970306c52102662b1b6928024bcbd183d91d64159c4c63c7e26418387772cad0594a5ddd88f24ad6ebf0630aa176e2e7fcb041e01a869fd57eca0cead91f2542588ea483d458f85df2689ec2a96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16266d583b1f2de24005842069830f63ec333d402e507fb1747cfcae8eb98874485d03f895fdfa5ef0789455986522028c35f8c740810347776b57b3deb43858421d6358756da5464c668eed94ade247d0502c8bf806dffd2690c17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc07ac69f6323c9e37de3842c119dffded9967527249ce01f679bae1178f88e113db9af9470e52e2f76aaafed2dfee6f19257307a5a7f0d9d2df34662facdddf85d0049ca5e883ae2bf7dfe531d84e0d3864b9ce06e9ed203d535c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7661368bffbcebfb4b7a60427dabd15aca28b67d7032a11aa89eba8f965e3d5a6911a8f1539936ad07bd8d3c994162f3bb6dd9cf7402493ae7f833254bd3345ce69d0c41f514507a007baca86182b620f6b1b52acbfb13126c15b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had5ad3c677255b911a9c84953eb35dd83b0a003956c2497b55c50ddb6c390528eb86b323fda9c16d4e3b5d6bb66a8cc919f999da4584a04dde93e23d530acd38deadbd4f06494d52be0a00f015c5f8f6230d655df6e7d27cd34fae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1328783f486b2887bbc5bb5cd90cae1b171a98e33df6d12bd829538139125ded6fe0209728b39e58f9b0a7e6de263f531469afda0e5fca5ad98c80abaf0e15cbc7372219af1db392fcd42aff02d5523e5813db61076ea6ff6b877e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdeb330564afb8b75ae779fb78aa2d1e93e6cc6ae353504757f3d067a0387cebdceb994b1d2da8667e765ef3d1a60398a5829859eea50f80301f116f7df5318963dd37600ab3434e67c6a0b915044f7e6051f6ec81396f684fd8992;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1229965979bef6804cd42cbe501055f41153732538fa1ba4176ac6c6d9ac011d4be0dfc951eaf7e2b1acfa3b2672938a978fb86505d802f0f1a8e8e32efb4769fd6d88e0e40272f7c2ed0f29f8120eeca022b768dae203b4d4e764;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c03c18a293ebd63e98b1ba3e957d113c625ca5725cea6a2599db73d5fba5298dcce65f2422b66a0bb02f50a0edf4924cac1c5d3e2c7495211a257669334c5d93bd1f4746dd9c4b9017dc4d40662033b421a09f5c46f8743935e52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdab9a6505a198e1dd81c0e4c3fc06542938562bde3de1288d1c93d9d5c4af712409920839246b250aa6a970013ae70a72bc0664176d27b61516ba1c2f7dd2676efca93141eb21502bb4220ebc41bf7c85ccbb2915b6f51eb1858;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h936985cfa43bf970cf14d501dec96b040e75ef832623118f18775bf4aed298022abda44180c7370693032a4b64409184e29a6ffd74b0699b4702cef6e6c7a75d04d7e80df919aed3f064a28ebd998750f48925333a33f55f62379c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e536728850458866e81eb168baf81b62a849239a70e4ce2e71eee9a28086c67dad70e14b5f5e7b0d162e4f13e12c46feac4e6967cf5bb920e6d408820a6c79586af64aa3d43c1fa94a1261bbb002d8a2b8dd3089443a7471fdb95e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f8f8bf58bfb186cb24d0a3109eca46c5a7e7c2c5a3fabd87522743860eabc52e816c77e5e58057c2ca3d6ea387fbc09cb972d073ee7752858cca03d1c10dc8fa4a3f763cc2969dff7b36492f7f9b48b8154bd567189bace8fcc13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd25a01aa8800114cf11e27b3780a2101a1e8a866cb8cbbdbca357263a0da76890d9db4f36605a43bc76b9ee86869206797e39b624d0155c5862e3b97c2179dd056cca2ed9d574d24bf62df74efa597aa3f8ac13ab0be5236f43363;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20d86edea35603e91b325f8d2cd83aac155d864efcf48fe27ba7e7d9f106741c1e8774ed2eb1f61b7fd10e32fe7261274257f212d7a06b81ee1f82b42ff8eb53f651eec9c3c144c61c6d485970cae11ec920f3dab5347ffc919cef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1903bbf6fb6e6eb19ccc5106fed87f006dc0ec0e70746db78ed8d03b95b6862d59efbb14fa9197fbe66e95a8b0227ee6851a2bfcbe7056fa512963786d74fd859a6eb82213d41edef160f25a0841e5db08c27c49d3769c6cee3a9df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d75cbf40b3313494a1c9f09eed6be493b56d83b75987fa956e50357975a580e6dba61759aa7e7c2d28df68c6406a53ac84434083e391b1707c4c0ac1c794d1f52e006183c09387b59137f4a7efc2034a24e10905f0a17cb1f03dd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd84213edd0a38b74ac46b3781ff8452d4a8ec4237cf2dd0175fd2f66e0eb4eee42ad7d2defc2c335a461f36f95b36a6ba72297e05d25b48fd3d64f5f2c5f880949431a28c5d26412105d5be074378149c2c59c50b10891e5cb19ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b787c5f0ac46d90c6914fa651c85eb66306a11cbea7027a453aa0b3ac35344c8115bcb4bd1d63d0ccff33cfb3a93ed2a2e8478a841c6ea55630ae1e847a25e7e4a86d056ca99d28bac7e390d760bb08519a337cace8086a779e19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c5293306ddc6a372e2a91cfcf676550186e018a994686f009cb364ac9a1488fa44946da1be700397380fc22c0fbd03a71ae12bf4c88614e90eee3a5e24b59a8e5f004be53cb3e28dac5856f3e4820d34a4d12c742087be354967;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb141faf50f2edfbe0e2f873d90a934e443a7029fa41a27a1017a8d94ba7eec042bb9ab819f24624566d9d130675864de9033178ede6a0900bfd49758f436764da7cbee6dcb9ae16100a7e59cbb0fa113c4278ba2f2efe6c7b9539f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d4166ce481dc132379e073a413c30ede6533a1711aa3a3709ad6c4df59965dd71517c10a16480ea4d7bb2724bbfb156e6b96ef114f112c4eacc0e1059d38ac9e5aa1f3ebc573eb276f910edf9347701d535c7370b32a5842a968b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e7bf22c96b0bbaca170a7e02dec0f368cae7a21acf15195b44e789d758681700b72ac73cd04c02e7555e452fbb6b1b25eca449350add431e3690b58cd4e8fca5ae61f07474c5d6ee3ea0b95b81147f5b4970a9d552aabd023a29a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d97399b9c3a529c1d70ad89ea18b2bc595680f70b9972304541ae408f94ab09c2be39bd0afed6cb7bedfdbc4a44197d4fb6789947a4d6a8400c312e3c91fd6cff448a14d5541fe27b4ed3797e4e3a2ea40ae2405ed3eccc9feb6b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h429e0358f76ca2045387952ce1de50be0eee11bb8e1f51dfb7159eba3ecfb6a6a2fba07aff43f9304527630bc2cccdc59736accdde312202435ef49f54b2e4ef296c13d6dd45083f39aa3673127adc72e949177ed5cd92faf35341;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11fdcb6ce55e01eeaded0da2e8b36e840e5795048096dd46a42d4de90ecfcf61a7213e30aa8f09d57b20190dc9495c28ff70d5e8a6c8c52b29f19128f239b1502cd69f397125d3dc682772e5add50bd65605120a4db657cbf4968e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106b3b40aea8a841381e316c3e4bd752237d56f287e42233b48d601cb0662bde49123b73af1e7d0814433d1f3fd40a1d8231b25c2dae1ed081afddb618ed54fef682e88221c50b278cdde6ce1cf6dc82167cf113907dda731c4dc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164e7229af311199db57f3ab770a31b0f23edd94ba4267803ce3b3531fcec51a088021d3517f0afa0c41b33bc9eb3c953709a06f86390df4d1799eac0ebc036d9fb9d819992a9435e30b43e42169c899b254bf2234fff0a0ee66e2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c38646bf0feb8f63be4a925300cba85c1274d3006c71ac14e494d942d5f56e6285de07c7cda8e5691ee0c361009e3b14e56f88934cf2c97be26bdadb5b0e386bc2c5000932629950ccf5747b0173986fcbbf639d95af11fd4dacbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142d39491d2abdfe9f0dfc2ac55d2ac147af58d648a8ba83221a3ff6accf3a38f390f6be9e09932523efae24a750d10d610367390caf244120eb749ef1df22e3a3b7ead8b895bd7e9de7e9a0eb4165c5d9993ceba4c3331c132a1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha82a7f7471dfa42feede6f74e892c82318db2fbb3bd0a7e2543adf56588aa2e105a1a11793c6906a763f01540b0c96dd7dd7c3532e4c060f509d9490f1499db1da147140674e7cfbb5b7c6664bb0a33630963c27377cf89383af99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h810fd020bd1616b3c77e0396267c68e82fae9b42b7a572754c0b09d4b65dd60d838fd4c481b658506c48e53e9e6b9320bba7d2d8f110ca3a69c48141039ab20d6a62bc030865ec859973563f19a81206e8985d18c6d621f8f89025;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95108974b4d8742f2d247f697c3e49efeace9f2cef1640fd553d78309597a82e50b96a24af47cede9f4bb6650aafa696b5effa0529c5cc5dd468299c05123dfa32d949680b8a359fda78c1850786835713dfab8010f6832205a53f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182799b71ca79f69a76c8e222e0f6ba7a777f62ecef8a0418ea070e8a260ca9db87d7506d02bb172bf46d5f6dbe848408c1bedc40c59a099923c120106556f7dd8c8aefe6d1578ca171cba6fc9691f65cdbfc17753daba325d819b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cc6f2e00152b5299c6701d442f8a269f394a6c65cd1b26dc2f6a40584515feb34f9378df085f64caeeeed3062b012e65efd021c7c3c5f1d8e8f924775db5e448df44819dce176992555ca5e0dfe4b13bb71605f56a815eb2d002d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105ea0ffdd36cf6bc9778a99bec52f5d1ae620e11b7cdbc3d26d6fc7f984540308ef3c5a831a19e2f57de0d074a03c7848d52ad7ebc0cdbca6adfef0673e49a4c92741bc2649a295315256e29611111fd004fc1d3b79c6754f16f37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d88a14aa8f2f44974f1b12f7d6981a3e0951cd37f872e815a9fb411ac804ec9afcd1763725e89820dfdd37774d64f6dfcf527baa2b8bd5ae983417b9aa4f866de650f07b8f86c1a785329fab1ac564d7b81758df356fb2233ed3d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5eda1cbf24617094250142812e31db4d764a349a5223c40e4c8040d2c92cfa51a10203741ce0fe70fda7a93bf5f665042937cc3710a8c607dba9adeec447a919c9c7157134943ad06b6ae3e271443d0cf56120be1b54ed22c6d074;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h398e00afe71edf907daeea7f099ab80b17e13a412bf68fc3ec88bec9471131d3cf3673125332f13eeacea79a5841f2e172bda5010945950cc58434dad22451a994081ae046bb8d62adb4f58393fdecc5d3c3b26ebc9a22ccfa84b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6328fd975d135ebce013699d3da06d548a6e23b30b8f10a29e7fb631b5702e62b32057c35acb12ab80139306ee68abd9e228a03bf62d2e73e587d7e8cf40ce45703735855eddccf7c13856c59b10bb18a9755f6cac7c617da8e917;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4eb973508ba664f225db724aaae6c94a9aa9eb4ca3a5b3f7dea08e383cf93f8de2bfd6f2c9dad36e07bd50611bdc874de98c32a1170b7f49c03947871255569cf46f6e330bff2927595f45e5f0e1f013430c9d53623a030ca82f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h734a81fdd9a7ed6c7b711fbdd3d3866662f23c1b200c25fcec4a6ce86f1a7518195edaab90642f04b455127a997d56127d9c181375f1e0d9d50caaec3b19c089a8f2c5604bb5a901427d220c80867bc923c0c9c73806dd550bda18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bb01e4a25fba66f981151561f13b829d174c0201dd9fbaf63cf18f7d5e4a315cf2490b7a79b7b3a224f462bb665a1e0cdea9c3a0cd566cd13249bcdee685a41a455fed353fcb14e50224b1e76f9ecb08ec17d64689af55cba6dbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109252f9f3cb7a6c98cef0aa115558d1a5a53bb7be885d503383bf62d2e209491531d77a325262568a4aa97667eead64f1038ec270988d53d67c931535863d11d11c74bd5cbcdde050b0c5df0ac5994b9d58cd7fff5eb3127ff10fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ebf7b8cd252257090be7c1412ff9fb4f0c33aadc2648029642a35772c962e9e37b38e5fd68080b2eec83404a5a9bb72bcd5f66a86af3dcfecfd53252ca7a3931a80bf1dd4aab19e3ad5b622db39e0d8701f57908b513e4d5dcabc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d989506e80b5cff6560a878f6d99b0c234042ddcf339c3879aab4119aa9417353d871665e2199f2de5d2b917e6beb37e8b6c30133544706f038207883a15f63971d580ad386f6f3fd1fb62249c8f0e92173a11ab56f8a8ac768a59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1289e6218b10b7bb88d9bf4afd6c1323ddffb8a63844bde147409c47f932c837960ffe471d3ca1638a944757e98c94885ca225a5c991eece14b5b85d2d92eb9826e137a1251a44c54d4c7e163ee9d3644fcc9aab4e38cce81144120;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4a6e6eaed488126a2b57cbde385db34a2f74416f2b8fcf455830700b379de2caf06d19a1242c9bed0b2f7b6752ea7d8005ae6ef1f11b03ac5d3377eeb3a67fc5b5c77a95ab4e11e1d8d21ddf995574e752c860f8f41c77d703afa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f6a4848b615c610f97bd117d7d189c1496adf98be06b2364b9b00953eefdeb426709003ea04d8cbecb3daf956a98d80e03a50d1fb7d39502aae30f3cd6ccc71d1387b6869afd13f6f6def6a5963d88f5e7dff3deb155adb989e05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h817224f15c91ab9f2fbef9c10aeee4a3c32ac24413756add16637ec1e752bb4e55ade8d9f47b1990009c40cedda5784cb28a835ed357f7d28d95eede143f4516e88d29d2da45d06e60e1f1cce940bd3f47ceadc701c4186a8e7f4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7e8900d938326ccd1ea5c8b73ee52c15e84cad0526d4bdeb01680ef98150c79df1014d016afb23b7bfea474ed661b9b07d8947d93a3c9be525ada1b3648c6ad31ee659ce9eeb806600913222c378d77775c30807f9b451f7c3600;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19091d7cf4bd328916aea9303c5218efafbede75cc1abe2371f17b242dbdff188c20837694edab9f40cf08c1a3711438a09289574e95112235a7e10dac10c28c438f08fd237aa7be0e4f393cf493ed266c0f56bc520d0839db4beda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32409dcca400f4f6224bc1405c5f62d01a47029be628538331deb7b51547f3f0be2ca0f4b30328201d75df301234d0d9b8134954d0b7d667963ca2ce67a6115fe1657b2121d5e0357c9517e4e491c25fa930d937b326357716a494;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdec30d28e286808d856f6b409287d2c0f62e175611a7e55e97502db500dca340c43084e3d359bb02e07b13d5f486c1749f210941e22feac2a70e5092e47dffd41b6867323e2d35bbd9e23c78f34199ab11b76615c885af39a3e91f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ad8b32cff75f6bd49177f13c26ee253ea4165ab71805703b9af0a4ed0135897d0be1a2b86e40d4e5378cc988363f87b760d9d07c9fac291dd8d8a0d5a84004f70cb9e4e4d5c0dfa15d6fd3a354f26974e0e644f203d8f05eec9db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187a2d23698fbddaf997bcad8d6d70d10a8cb0352b89138095057b462734eed3ed2847dfb47074ce2eddbd2de48ae2f7d930c7ce008bdd6f360266fc5ec55335aecc82fa9f9bc14b53f9a445e6e78b27405b2e782f1bf979efdbcb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a875bf245be6742dab682166b835f40872208686ff565d525d2890c26bc94316a63d55edc892e85a7bec074540daacb622334d8aee7fad5d9867a3d29436898833f6421050e4e389e6ee87a5da2589894350e79d7dc780f3e3f975;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a456b62b0693db1f94d174fd929273b07a516633342d13495f5e455d6ff5e31fdea203e96f1dac1a3f532ea3a5c68432d7fa3934b8fbb2b5a15509366c1b60d5164f2be8c2218ecd01a5513d3cc18d6a58eaf782619d2beaa53980;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91c7072591fc0933513e0fbc1c8d94c4749823cd17a8d2ff6b26856a01b3a52748d7ea6e235f4076e2e8d9c2afb992858dd6d820c0aea4e1581de64e9aa95f6bcbccdb32037f72a87e9bc9d817f5ea60b2a6f80b597ba2cf061c9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cf4541888ae347bd61bf80c1c036786c24d91ea6a4b341e936d6ee7edb9146b2b9b748720c64554b410b3f19ecdd6a9e5c413ccbd0bf89c99b463d75dba016b6bd37a15ad7c14eda39275b6275b78cd51907df48f749f37f2f3b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c38d801c9fbfaee1092fb23c437980d56845963d722a7e8d338c8bec93b86cd983ef853a376ad613047ab436a2594216a43215a1bee6e42cd34d8211a5ff73a5145b8885cd898c169a0e3736481d56039cc6bd7ced8fa65544cd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h415c497da080ac5a32b9a3a9b4ca029fcae537eb6db456b55ad3b69095e372b31e2a30e157d68f1edc7677bb0afa4f25dc906da140820e001bef353a3173df418cc2d0471679f6a3e24f40906f94a4e9e36ff5e02c88d749fc3092;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he07653a5dc6145442d2f9ea8d826f2b8aea022e24b76e5c46d3b87c414ef4241ef01d85d721c60997b4f6bac60bfa6c3ded2b24edfec426f39f27257c4a9ce8de1d39c57d910191478d331d41eac4b17e24e56f566bef8638f8d14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd87d82773c8f9c3cd458e7fd9c4f6e0785a16f165c0636285ef369f6826c69f4e0bbc4f8855a91561c2f1db7b77841091210a79bdaf089598489e7a6d2f1eda77f27bcea40b7c5e27e609e48d5cdc92065e866c0e78e3e3a482596;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb56fa07fe3713f202bb8c0c3ccfc1e4e296e0560202268ab5d03238f9d336cf3deb86ce9e34fea35b82b31845b7de5430df4d15c064d0291bdda14fd66b4dedd5b36ae6f11661d90505bb3db411be5f7239a09599b7bfd7be3237;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd85abba67929e87785d58f1a943ef3cb982a8acfcf75d4ef31da262ea53f7d0da8808a97ee601fe7b619c991450bfbc26cddf50f7d6a44b192fd55da212a197112fc8fcc3766c8f663d0e32cabe2af13a7a9c458124fb37c06b951;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1700be971ffc931380b2f84415f25f262c8b37a44b97219f1fa33e4c4a9f5da5d91c554373ec5b7e1cc51c1748d84b35760f0410d7bb5126b3e0598e5ee5feee0a4d5ae070e078455317045ba871b1b51d10f9a3ed331256edae2d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1258a07e0ec650e0bf92e6f6db2b58490a87a953efd111bbb00ea57288e454d5b492db004823f628f07bf58b27f933c5518480ffe522b82b9ef6c355aaa5dfbf3eec0a2e2fb3790331616abb49f5da4457a4f833b2325d55535111a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95491cd7a696b93721b056ebed8276c7f30d5d10856a8524b0981b51c5fa8913ebe6f7f12cc6904e2eceab1e3230e81764e8d752cbed4a5b7d3fd225cc0c96c971d956e2ee4f28439a90a405bc29ef82a234e4442bf352e6a55940;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14de863625aa8f480708998e49ddcb8a3e2213adcfad44aade37a38f5c44804c5b9a5b42995c3d0bf6a9e3a994f6e9395d0c92069548e773e734cf89d47db0b22439438e1aa64530a750a5d680fca0e18ce254d378924523204845c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2c287c35a8df48cc8470ec2815090ed935198202668cb867838b66fbde687f86c81308b090e9f9488da9d2e00e36b7d137382ccf51b0f0aa5d6a4a4867cbd68defd1a2d98c1e87eea62f9156ed5763ac02dbaf95e648cd8144d34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9831ade2e64ffa3e35ae21d4b99e6d33fad66207c98a42138484aeb2b92ad4100ea91b103cd6aebb0f83b1b3f85e04189d2f1ceeec8a405d581aaf2279b09497e087fe3e608ee562d6958e7a22a2ee0e1d49ce644654c9f70f7bed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41c5c12f44cb0ffeaf3c507664e89aefff63ac67abac8a46580eee66c2df12d1846c1f65bd29e1139629dec1982cd55d99996e963b11d338250a43d31911627e5fc8f5f6e62acd18ef170ddad1cc92d880a83b09cd4ea42c4993;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aea754dc69facd46cb7623c66f6cbfba02b13196c9d44b62906ee1b8cb89d289afcdb7dd7b7ddc0e9231181a591cfbd29d8461acbb7ea593f05f33e9a61e526858e3cfd93a954f430c0033e46005d78e2436498de476eb2f86810d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c47fe4f5dad6ce13aed333027ee588412ca2581dc0f6691ba9aeb572f9da75e481f563c3512ac7e33b9fc0392372d92fed6a1dde36f034ffc66717eaffe476b28e90d077c823d76671966930e4c6e23b75078482d4548a2d4d4616;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ee423ede6a0747a9941b499441bd8a583c1add79e3c18937355eea154165b2370248104c96bb1c983e0456bb8e7abada0cc84af1362488a1de4908a98d47ee3da3d68b3465304c918d5cd2441c1cc7010026f85fe2e184fca6c8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91f3e6732f8ba9ae9fefa6824f848bdee1ae71877b90108de85c3a8c95e13ddd1c9872a6ee25e264524d23b1b274b8c3e6602a27f18554123d4c45f6d2f8d1dad3c3f94c549ffb7bfdf879768258e442749205f55b34b0ea7ea21f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeb494051a511e405341d11d725f3529cc1e70cbacf4112a8729e6b6b3445d2ecc6ef85eb35664ebf90cce49dce77c0050f1bfb9b60a877fd314c3bcf26e50b28413c352a3817959577ff0a719e40509fa836cde984602a086b72b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4e43b321ef7c022699a84d4b191eb1156e12ff785df6f92d3914caa00e6b8b98fed334b98f9af97392bb9d6c9d8052fdf420fd35153cf966a32f927d8381442b1fe8ba33d25e01fa6812c8f7439fc2020540acc90201ca2108ef8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf07a35a533f4edeadbe879748987371a7f90296eba3a76f0f2742b4fb82cb71595f52c38487392e94bca8afde61c646e904396cd418b7060ae806e04f6434b015ce9c64871b29df8e4f7a876fc4d2bb3e0f3753d9b62618f1162b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc77bdca75027554120545e94f26a577ddc12e887e3ba1cd44ef39461424910d1530889d35bc9f2f1be08dd8a493c73282908d9f498aac14a384409b1f509c7a60eb0c98079edc932e26c378a642c4c1d6eaa046dd5aefe703f3a83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bdcc61a71205910cdcd9b340338148be2659ae32a48983356d386abd7544f345f125f48909b3da251c86a063f64c9fd781a0510a9c44de2d55ddf7a4dc9fef8cdd4e90cb01aecaf4c14ad98c98d9b930cbd0a356c865e12626f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1220e551ac03333df5966cc29a1eed865eb8bc37076de4727f079fad01aeae3b0da146b38c70f33b1b5853764897944518e5811f25a37b12661390d3fd3457d1aa4b8534e3a43a7b3e95e872bca55a4f8f3ec45f4762ccd8890cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ce6657c29cc640b0f8f8a7e5c2f4f1c282ca7f6a37d5df6d72db4577f1a6a7dba5759bd80256edab7adb1feef7a2222d2de55a473bc13aeab7b0d8a2d7802f63e1d1b74015a64f294dff6da4b8d7f991b71215ed9e9ea63e664af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56d0e80d96d99ac28be1f85bc4e7b77ae6a493fdd846c7aa6f75bfe563750646282f17430fcfc59d3646f0c0e61ab290f93c50b9908f54f92882722f269dece396413bb7110d00f8f44665b65234cbd321f6eb48e6eeda1f36155c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff3775afe70963adf4c77737b768c8adead5e9025b5ab516ae9a86f8838f5ba8d14209fbd6bac0c38b56a5362764e17f61c27330eeb67282838b44583dbe9c9bbde1a912dc6670fb25005551af680d311b69a54a08a25d60828066;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1676e3f684eec67fe13356e688b84c7df94a0088608618038142ea3b27050878716dba2f91254f40f4bdd60e50fbbf950e935a3d87e26a4813b7a1c92508838d4925271724d34da681e6c8fdee24cb613eccf675c2ea8ef4713029f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1585244cdff3fef93587be2ca18aa41a4fdc2dedec797dbfc20fbbc2f1b145a0091aea7cd3f44c9c01d0d1c6dd3bb5056b2b30950f55293a6153a77ca5129575dd1d813398a1b18e4bbe1613224799294a4a34824616f1260779da0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41750c4ba445a4309a42b1155b4bf4504011c4ba765437fa944d0d392ee4e9dbbbae4847c72fea23e3780c358dd9fb3c84bc005fa69dc0c6d43392ac43d7f7ffbd7fee8d7b90c1e99b03ea540022977b494260b42ec56121fa5e28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdc7e3655ee4adf40b38ea46c9c229274682c36ba6ff6cd006720e38ac348da34787402703384736b20b5fba74c2031cc2a0542fe48be8a2efaf5ab15e75e1468708a6cd4364a56fa98b0abef2074fde0130d0e7f7948946ccdefe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43adebaa77b7531bc7078cfbbf0e0e8fa0ba3cae65c47f683abe31abe25a3032e44b606d62229470e889c16863db627b6ee08e1e8bc2e2efc732ad830fabe43ec9cdcac6e31848717ed5bf7953513bfd7fae1feed0e87c213d8ace;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f5246f8780aed97304d287917f5cbfa6da48b65b92ccfb0748d453f349d71f386b24ca264bf4ed9e9c6cc4366a5c8dd49ba12436fd2261839e4e4bedf2d53ecddb5de04ce44c309a25c6dfa48d96e055a8678f68a77778a581087;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ce842ed7ce5fde8b25fb903b66d8ef43c04f2257cab3db3b6de350f5d47ce6d0f991c8652a5e185a1b9613f176377a32800ba4c0ee849762c40b74965ed2fdc9c4abc32cc138c46c4959705c2be3ccea0fb8ebf96673e07bbe914;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11765892cb1aa19b4b6cb20d28ddaaad2b5275ec5b043219b3528f966fb038475fd99016c686d9923bf5507acc2f1c98ebc957c060bc9441be1dd3948ff97adb22b28e57aff7c68e2d03d22e6c4c9aef79f8987ce727fb3b3d6f43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9275df028464164b1373e15ef06b2d0e0aad1a417704976359d0c3024a806bb40c3335259a1903dd41a8227a6351d7e845a1584a6d7c1a3524bbf302fc4f44ec975a18f8437ca103d255e025dcb1e5821db7641c42c373008ef928;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19dd8b704a27a294403a6be60e071dbded80f8614dcd30d0012a2205fd755424352cf285a2ff1d6dd6ae6f45deb89bdc87f313f69143557af330e11520648da316adf3c2f4dfac90c0ae0ecac3530276cf3090b9bda92d384a72e52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2503cf8e13dde6d8512f31a11f7f696a1ef481ad4b133b0237763ee660820d21c0bfa344de4f486f4091bb60ad1ef57821d4918bc799ca8db248cdf6fef94ec6dde9ad010a8c209de8ed5b00463f84ba0ebe702b4aa02f6a47864;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8c64125e93a0ea9bd4d9e987831464d0e2bf1f9916a01a8b21f4cce98a900a8423f64abcda73238d08f1fd7804d6b03e8de4bc40587ed3c98eba96febe982dcddb7d4a6199723550652140c96d99ee69ec081f4de5fda03dc6093;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb61fe8b95464d3cdf0c2b742fe9024e3b93dc773aa6058f77f4ef6cb9c105ab36d1bdf3547ff368d8b883f7f3824c17b2a78b2616061f51175702751cb8f0fb591bea63cf617a908abcd3f5f7c1b5db3590d819c7cf99dce4ddfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bd55d64766af50203e171f8eb78adced6d2df5b2ae0c3a904ac25a4c397eeaa7940c43ac43ebd8b3989338257f4b7ca267f95ea440535197c5a1c10581180df128d738a91a5b64a07dc34982f1912776357c7053d463feeb7b13a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2bf0e979773aa4cc1cbedcfadc2248c41699c608977934575a4def65782e2f16758bd677b37cb6c91445609bf6e0e40d6ba87510382be51d54692f21fb0b45804aba071af872e0a46add5108c9af62383a4ccc714618bf04c2434e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha21413e764c9eeb4b11f0b9d38d3ca2f5ff44b945ecf789ee6ab89da726028d38067a0624fa1b2d23a92a02b33b8646a1cd5095a9820bb4baad9241f904d82216ada8ebd5e5481c4533adf40107a9e4bf20804c8c7665734eb6111;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ed3019e713d35629979cb18d63a8cbeb4fbc5aba017a9e5345bb77fc90c119d698f658cc9fedfe839d64c52d24f81362daa951023b8bc73920dca7101371a0fef5971f6443b92da6b397daf3145f7a6c276d95e3fa5759140e406;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha90d4537b84436e62beaa2babd712fab6a4ce0fd83fa1c48d8076241ba7a485f0d5153b912dd23dd83c824355a96428b1b9f1fc8dc0a023fd43e138b42f0e9d53d87377062b52ab1c0ffd9ca3069e9c78a8159b65caba72dc98176;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef4126107dd72805af42f4be248f3d1f14b2888bc790fae4f856680cd3480487834ff05370fd26f93f72c4ae8bf9a5009f5fbdfa0624464c9f73a32e79f701f54c3c8bdf367a743cc775d8b73ced90fcff7bfeb2c7e37775888b84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf96560c9434e1025341aba5d5f5b49d135297000c6133a8cf7d8ab65c6d75f9af3091d716a1e6f3420e5eb6c6aeb765bd258f99b3de6637b0e99384b14585876ba366e19b46183d1340b656c726f354bcaea30df29b3fc16a23a60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc6b6a6dd237860c476476b697626db5a1b983cc5bf7f139819bab8c4baa43988d9ff20417b10302b40bf345d144c2c7983dd3af60460c4a4195944ab5e77626340a83a51d5aefb9a1b243b8dee6af9ee5d283e96d73ec3c3df365;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2f9e8bbc7528c9b32fa1cd212348d9e588f8e74f12b090f0d3fd075e005edf3e7499e48acf48f6d88533e07d51bc55ba1a0dbbdd0195a33aa047c3bcca4f26db6d6fc07a45307d6537ba449f9315c3f640d55a2b4cdc466ecf663;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93ef5cf4177423fa0e4f98532d79ad6f39761b3acfce79b6fb9b6d5e99aac1aa932afcf80f832146156c3a36b2ea11cb6cb5f17c865fe5890fb6b4192f060fa9bbfb8b2e05f53d4a01b388ed378c80f8522153025ca558e8227786;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba7ed66fcbb0c423321aa93e3198a0a9e4c305aaa3c26c52eced81af54b37ee0849e54413db5bed29d7a5fd26deeba25ba579d97226fe82d234907b789b05f1736327b03e21e1230a60b37bae1c57100a9b23157d5b64c62bc0ada;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18295a705bfe852a819068e919d8c5d2bb0409e26de0d73204b47ffaf46dd2271f70ee9cd6aeb36233c77e159cfa78d563f3791e11d81d7c955a1d73633fa4a7a20a3f963b95b7a07dbe37f6d66cc571a738d0d9b8b065c06484876;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61d9bad530309d1fce8d2bcd68fcff693c692cc13ac224acb03672c8cda2faa301cd0faf7a93810c635dbb86926f6d7b8fe42e664545b34c4580a924747c5103144c20c9a8d62e86b0ff49f0ff59e39164f64cd8cf1d043261d963;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2634bc7c69de95ccb4ec2d9dea316cbd1da7183a1d1071233a8556166f65aa900a4cd85e396c5b944db32f4f8465104e982d68d894c65e01db24db25da609200bb9abda051e347545d811304b4d3d8af793677a1046b2cf102267;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a206079c2bcf0de4c016e0925ba30a88f730b075e5b222b4672e7751d1bdc59a3783dd691497a48c14bf7351c832b146bced6dcf5332467254c7b501534a5a70e4a1f36d5a91069ad23cd87d2848c317fbf1c83f8a525f5ed04f62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1938d797a6019b9d67c73d2e944bb1a190b68007c581ca2a2a4e592ce4d31d8e743d56266ac65ac98a9cc6354099bec150ac6c38e6a18b1d8686e54f508322cc0f1de4b71432f803d9e1ae6f675c3ec1b75890e18b5f15b6adf2a5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42f6539c54c27424505dedf7f52973cf47dc974b2527b90a128ab3457a180b9bfd2322660243aafb1e9cfdcb29c24a1513cd39c0d45a180fca6e5ebb6026aef9251588bc82ab3999745af884a166bed12ac95514148c7de1b7835d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10404b690dc1660bb2d8a4170ed82ba9f0ee73efae23ed2acfed2ec05bbf7c4284c6f9568f13b6f86e32ee95c0d5a8d2c4e3db1b4863a5d285ae46f73dbded822441a997373bd5935cbb77ed1fe8abbf85d4008b7db6fe58973b717;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef98a78d947019bd449bc9203d28033060fd1c4f1b3e05ab531c551018213567a7acda28a0c4ca07472fbdc70a342c7b56708cb8c40f82dcbc68dc469ec85d0821777b0ea2ba2bf068f421aabce2a11ce10c109f4cc5960b9ca633;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1220bb0abf966f53f94395a28f65b97f025198646a6101a2e4ea72c766543a8f9835f52330101574f3fa23ea2e2d9c05a4aec87354598effebd8a329db1b92c9c607775b4aa25638dad5f493f51c02c4f9c673054186f0a3967753c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb2fc663d452a31cb05d578fcf79ea98dee8a8eab215e8f7f35dee89aec4295fc2d0f2f7acb9f6e8f421ff274e89a00f7a9797e04dc34118fc11c667601e05c80ff593f3e051345c610bdfc8e5b4a6c0e3185868cccc4117b7cd59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h540842f86201e0d3b6fe421bad9751631f1532ed65e5ef503bbebcce388e361593ae3ab3ef9b1dcc7d2bc2c21dd8814c93275544d97d6b85b85cef0a307fdabf06f645323739e6e4c0d8558c1c891c55ccc2c40281926d07e74dac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbafae1ca91cb742cb3deebdd1cb77413ccd697d6665616e16f2ea9a10718502039b67ec397fde9863a2557bdc8d66bc3a02ceecffcdb0749e77b00ea23197ef53c2a8c928c4be6c6b23fc58e7a7e0d0dc9470fa2debface927b64b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111c6d124eb9bc2b946d7d5199b199d4e321507725ef24b02686e502aacf6357ab34a74eaa463dff6cc79f2d52e5ca5a4a46c06d036389da9073012b0aa20f6d04d05301026e597c589a8e1d861ef4404ec7fcf116a2a530192d7f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92600a29b123bbda416942f9a6f049f49306a354507e31a182e23fc90719fffb6056077a046f71eb308ab41221c338a526006bcb4cdf977181924afef033e6617330505999ad76b9e6e8d7ef13e8f083ed13bc5469b9615446adca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1debef32107d6c89484c51b6f2daa74ce2c6014f212b70ddd3de10448aa6c7f2c21953dd267b01f3818acccae171b68c5dd3aa65644eef33f46a5198730281bf0222d456056a71d357f7cd0887b9402d98ab78c51b285efaa410e10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125024ba261defef96241830f252d048cdf75dcb3abbd26363bc808585770c2304c2bf6588a84039d2ca72674feb826ee4be1be4c2133db98ae66e1c24718dafd653a633aaf3190a0d41d5f8190a66760585718452e59f4dbaaaf25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b7632d5f3eeda61ae3c2ff6d9c154ccb60d8e652839f5bf3301f31824cb8b68eef435e8e253c7ea2bbbc29797e6acc20e689b8b68d4bf7484be4cfd0c6ee0220466c1586a61e6c72e9ef84b4e99e4f0d10e04f42f5cf81cdb1774;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1925563b589888995d45c75718ba8ac996a0ec711704c7be1b93a9b70f4521f10a7d8ee729b272a615d1d19281c771a321cbb8d6a9337ff699862f4c72149ea2dd400c1b85c9ac12f97dade6fc636a7e5d74c0f888a06c758a8ea99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbcb70e39d286b3f9dfb4a559a5d3b254fce1912d5d460873ab1a7163db016b209ced5ab574ed4782135e74216c52621e8fef3fc24890cc9c7f252a68a357065e16eb4bd643376d17bc04cb70d9bd221a14a56235bc1c67323f0310;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2f6325d60b6be0b89548af88959474d8530eb233fe6f8ad56eae51f8e23a74a2ebcca97d5115d2112027a3810c6c7de637bcf03603bde89a1fa6a7d3bdb84a02b8fceb202b49bd90ca9301e5c89a0d489dbceca9e0270685c5e64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199bd576a30ea791045f898bfdbbc229555d3a23900f8f64c634d4c278353bd414e115e4aa33e925bd387e0dc6e3c788a55380f2b21e52f6c57d0b3004a5a3b6b56abd53b687b9f2d5ef98b8257fb4ec1d9a1656ced247958302fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141797b39d754eaf12b8a7c02ae584865b2a677787be5a407ab651d500b5845dc54725b593ab5369cd05edb00f88286ee9f4c49191a40219e38e94a6c0ecf2eba433c595a8583c1e5af361b7d5b97ec67cc99f2604dccf4f391c36d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha88943adb237fb82b3e78b19e4ab0211a34e91c3ac3e6b4db557d0240cc0bbf10a2f0120a03afe6aec8c3280e0889f108267acc1ae581ca2adeae302c44169cce4ee2f38b9529a7c5d32c94304442677072cf6109e8bff8cbe75c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde819bbbc901ba8a3d6d38ec71ffd3b04a4312e66468c327586fe13764402cd40b29335f4013848d3b93f7f50e3d45ced80ebeab1e5c78bd07aa105238ac5f38dc4ad5c5fdc720acc6f6a60c70f92b28d5db63972e950e84b8ae1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd6cd46758bc250626f0f3b80d75edddf33e504b47dc842d62cdeaaf737f5894194a9ecd894dfcb9c1071cddba60445bda9105150b2a34616e1efa89010fe6bf68c9cf272fb3a0a16e8120351f64618c8b1044c74f8815f9ead50a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50396a3493c0be49e27390ab79015b6f257d8f769168dc34536f6cdc1bd99f3396ce47071b9414ef5e01ae826b33568c129fe34e1a8573a7f5264d34e2a865c23ecf1ea14f81ba053126e05fdb2e41ad4e873d1b62d6023da782d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84e5171b451c16c9dd089e34090f1b2d09e87be1474a6b644d921033d940a5416807e72b1910842f18c1b977945ff083a5d1fd0565b1e5ab3ded92693ff0c5a05bb25866f62f580919af9b78e64dbb11b915832927cbd7b9674065;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h284acec5c1b4e738bacd3d98a40cc0e0fcc0d8cd598121f2c245409421c601a707c8c1acca4c4c07902900a209ad8ce24fe009d15bdbf2956a2d734f4022c7d3a17fc5568a2282482e2bfdc723a3288f4fe5252f2abe80aa8a4408;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h926acdbf00cc6a66b8f066dbc8b71bcc5b8a3cc2614db1ad9a6b0c55e25b18b41a81403e5fa227a863fbc60550ef721d2cf2a2c9fdea9402b812e4e60761fa00ca9719c1065f7c5cdb0902ba848aa97b11401d1a3da238691e730c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1cdb0f14ee65c11e75458cc2d88a7ecf0bc2d731a07edd447868f343abffa9d8b988be6b185c1a16370db1a84d64ac5e9638f769f9fb5f787947e25258272ae92729b6e402367065a5138440181aad96585b5534ce2f953c0f2e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51cb3d5338bbee57ed36f75835a9f091af14191f1d2552a5f71c79a6c575131004584ec22caa0c0d951fff681467759054213d301aa0d5bef3b8203acbf908cd743a12fdd0a62e6b9923d98e0f1214f8948dae051b4ebaf6548a24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5042c60bd20fc60b672f7b59aa2b3e31e56aefa760393681c97c9aa1da2130f72ec4c552fb433a2c3284f344b58c73a13f5cef9714242550d676c3c43fbf9332511772f0ac1b793142b28acd0b83983abb4b2afe2c0e850d7f20d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d96c4dbf5e8d8594a5c62b8e292044ac761f92a60ccfc160fbb942cb75ec10bc9fcba2df0f06b6755b8b86984fe4fc3fafe69c9936670a45f68cd2322e333023dfada9da9221510d2da0ca82ec644c2e31658275536a967a585b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db49a2501be8b96891168d895dd83aece69913419168eca170bdf8e7328cd1ae69a9fa4e99465d990597b173266c0ef0c30838edc00a21cccbf1e0a920a9c887cbfef1ffb02ff92e032d7962d153fc5474d1bb9c0ff20b40757f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5164d75e14e71ab0e1dee7e04a42b59f15f16161a2f61eddada371e261b66c9367fb1fd16a9ffe419a38c5d016d1ea684881c9df234cd5b4d651f5c9b060a6046f0498d6700f9fe2866a168fd5b6586f96e0d5373315a77d7d9323;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12751f6afe155f16fba8a31228b235ac3d34b9352da6f9287c38fa1bf340f411910a78d2cedcc03ddf9b8f0133cdb5dcfb341393b3081166c1776d62a2a8a90e8d9101009645fdbfde946f7d74ee132facdbcfa793594b8f9734102;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa249ca6720011a788719c3da7e4cc322f2e164b354f62a048dcd73753f803a052f0b89c08a62cedb59b5536aa3cc74b2e642d33c7a0e92aed6809885b9aecfc12593e6a91a213428e5c7abcd0f27c57fd762ed5947f031e135a36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a455fce27e2f4d09e7df2793cc32791202f04bf4a2af80d3d9251f68d17f2b6b6aa21e7b3eca776b1470729cd092b124ecd07e9656e50b1788836f4bdb0e063e8227d390165783af0f9a035adfcc30a00344bd1dff7fd2be0f359d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144a8564b5600e64ab081e8b9972c99ed25c89aa3e982479c54c14a54c1fef2d538106c3c9d426ccb5b5bcb5d96f59430b59491520bcae5df472a7163193a17975830947823e74ebe7819d979ab2cebb44e7f9d71c274e00d153b60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f31ec6446d959195df67d42a530ab065a965b55b6776bdb58152bd9aca1a0359fae24a32ff896716a11417d62f9339a4176cc19855272324e724d636860ca58b75c15f9fe7fe3168ad15902fc2eed1c2b0ac50100068ee17398db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18aafcd1c01be182ed1b363a734570b60b3650f3809c34f194619727cb8691c8525113192c7953158c99d5db2b7d69a9e0a5bcfe4d8e27ff49975a99ffae73d4756cf94a63218e0d624473cb279e3e23ff10ac1e01c459958f17ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd98327e6cd07360ec2f84c229c86a6bce8862a75045231b30e653de5fcb93eef08f456b759150fd1156190079cab5e2f49d52c9d15d53bd2344d70cf9ff6482c6003066b0c277c091a621c566ac1488417fbd7990942473604d7ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efc721fe4969ae38ed1be114f25405c645e7e3de69829423e0bbdeef977a73e136a0fed4415d6432afbcf20fa566f353247da3929eff19a779028952e51423203013ca0915d45293f4e13900b6be6f6486b6e347a5396895a485b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffbe5ce08f4ee8364ce581a484a0cc55891bdf4ee501e9e5060071d60c97b8e58d1abb058dc04631d69818bede82dab62c1251143eb76f2e23d060fa78507a9c341541a60af0b2faf872b629b068dd5e2392a538a57683e8228f62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c74750fbee255f77a24ad6fd15a244d01661fc90fa9099289e9aa549753ee6054d4e27693dbab541d29a3b5a26fe51c79718a52a9f7af726b923131f8c042f4d652631b7d077133b0aa829aac26aad6459475fe2742233453da3be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55076da3728124eacb74caf18f81581add1193e78e3d5e590acf44b92d5a08da7c0b24bc470c70cf459e06f3feab4dd13052f17d41131ba8b642db30e4d92341af23c5aa23d00416dee3de062687f6cd26443a5f41b87c7515e3f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16da32d897290de7f22838654f1a415cf8a8394e6fb1fbff48d39d9f24832522041f52d7ad8d9a81734e07682d9da886e5d9bb01f5b42945d52f437ef732a71a36f94100ad6e84f30f3c9135633d75ac62a2fc8a131f70b1b41d94b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2a4399db126945fcbf85824aebaf9fcb7d55e88fa86d7d22a374e352e3c4f1d2a1ec5e6fafa2dafc10b15db9d6bddaada0684054b1856ee2b1fcf67637109425acaff6ebe05649e4687fdf97983442a998b78bcde3375882638ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf147ad19dddfa3cb2bf2bb5b3afec8beb2af15a28874d62eae0715cd31ae5b9691f6a1f7e60a6a4a64a06d17cfb119ec6486b1d13bb20b67c805b873a109efd70287ba9874fefe88dec0c5ad208f4267de7487a16c97c6fb48549;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h404e76086e1c2ca6ed4697c57c3e19f889608deb78f6e5a7f6dba9719e283b804124960d548bdf7744318033ba7886392f715d76f6296552dc79bd307eab934aca1f738adf9c753714dad3a8a3447a972a5a7b016dcd936631abd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1973f6cb852c64f62801154d3b79e49cdbaacb753ffbe88c8078f9e500079f151be63dc72d2cefb5e49cffbfdb231ba522d008adfbcdeb55ed11c959d7fdaeaff86ce2ca216e70ad3ba10905fa52934324d1c30e44d8a032579f2ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcbb9d2be6bc659ef36c299c1e35d5d478a3c8029800451e7b7f5d2c5a6d8ff49f8cd041ecff478001611d66aecedcd8c99c21974078e08d5d063daa8f72e5fa670d2854a8b043a39d60b1d6cd37177e318d98df6d4945d162a829;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a90ba05e1d52aafeb9efe5e83041f5d6dd44a18f419fb914dc2e3ef7004e8918c8d2f0cd58f10930fc978f123cbb76d95db8b40c5d75dc27950dda4ba6513c082eba7fcbe4aa48595c582f260e41e6f909b257fd1b663a136bc91b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfdb89a83b974dc2a4d5967abaaae9d17adb8ac73d6b488d55ae2468b6829af89bf9c738fc5295de0157992bd0524e4dd1d710f9577e52db13ea2d3159b99e5c14ad4330d256bb88a26765a878fdd0d1eaa059315adbc919878eb3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca91a324835488500e73832311a1e4b870a9dc3673799586d45adbc92464c159846d5edeaf8e0acf346ff6e75866d0b90b796e8dee372230e80407717d2687b0676e7c03ec6e587a1fbb65edacd1044c38a906b49f37a4c0b96c66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36ccfe8475da2a0c3f32751153da7ee5362ba58b44f4a41a4d780d45c2384eed8ded93f5e6069cfadd0a55aae51972512bf46cdf50db8060bf2eceac789c795499e4327ea3b1cac79f40e6f2581c30f90ab2d3b2a35b349663546b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116c28bd482b63f5daf3eda08e22e27881db8cc0b62fa78bcaf58593968214021282a13f55526fc8b45c9f5b0c317882d1b2fb8b59f3520404751490b68a1225055c0ecd7cdfae3b41a04c60958234dd560ea8bd1ceaae9b4a6d468;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf050e54420775e1486969a2cf7eb7df1d80b85882f6731a44feb7987945e66242adea9b46aaaffa2f8448d079e4f04c5f93e47053a4d8b1448e10101ac656f5178b2780051f390f05c8fa4b743343951f4c933f0d8c927259c55e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b72421554ab29b0bebe304a87e02e5b83f6c0b9dad36b4fa040722425b77db4f6f89aac41101274f25a5d5b5fc1c02d4bffa4005cf983cb757a26fb985d7945a34e84a20425f231cc7c863ab9bd55347ea6840e267ed69d13668e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed3569d6fe3170d141abaec91f4c9e1f3daa57294cdd38600a5609856cb166802b409e40c6506656d493de457017b42a4cfb39c06ba655071d0bdcc7dc621df154cb8f8c3318a6c076b05fe1016559eec4148795571d6477953904;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b1227988efae1ad1be29eae7291c7476f02cadefe7bd5975054bd588822c57862351337e2afffbef347757151256ee5b967e3e0fe7e89a8032e8f645afd313211455c1a3fa62c246c55df0466a59fcaf59b6fc853d47ca7bd12c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefef52ca6e211f64094c9eed63bfb3c0a6f6e0ae204dcece53400436d94093d6bcbf6b592cd4b4929ecbff22f9ebbf45c6b98744b9e7d58ad743bfdb60228dd0346bba9190b7c0de5c53bb8946ab4896f878daa80173277b2b17d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed7db6e11892d5591e9e8ac2db83aae1dd541a90120f5b01dfabe9dd81875f87311e3d788c4469d79b3137a5f109dacc8db6ff68de1c028626b27c8a7333a1761cb62e8771c9d11d5177645adfb153321112d21f949bcca5b3b312;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1adca3627f0dc8ef6f997a8ccf51f0df8530468a7ed0f6408b38df03172271bd841399176e248fe61b718359ee72b8cb369417679e3c79a3a0c639b52310ada1b683096f95f09ef53d411dc117e930b1b7ff0e879e1cc4e361e485b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15af1e9991b59e8d325a582806679f6fff1b894d3150aae3d5054b67e2c77e44d54f29b49747ea1c81190640b9addb559ad149e8edb9d2d29a9ff6f8d444e74f4362f053ab8a8c11bcbf96f4371286a4168c29548518877210bde4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1883eab20c896da1a1f20b236d684d44cc1fe999918a7a1dd7653e440a2e092153fd250c555c592386a59479b639d870ce3f6bbcdcb64f79c3b4abc54f7477abcc6c06b56e758cc832302b2d073e9bc0fa4f24f898bce6cbc1d978b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b71fbf11a546b5e52c6342cfe8b624c64941f15c1d3c9aa5f8161e08a62ba6936c78362775bb86d70d25a410dc4da43f9bb29d8df0235fdd590ebd9442842057f037a8825c8c4a5b673ef4785f184993af23795c669722203e392d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9b5210a959a2b90116b5cb9cc02f6ef5c904a215bfe9e2480e6dacaa1f276baefe05c133d2a0ead3f5bc2dbc52593f1669c995d61850e375f1334b39debf5fddffe5911fe71538f8a4aa61da17a5543a570e106a03a7c81b84b3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haae865b72d05175b17a4f9d6f6dcd6458da26a161eccb67947c05b2b6798ff2cdf99e008dca752d635a719ba75dab5742ca5621cf89cccdcd64047e632d162e701f40705537d2ce2dbcfa92cb9706e67bf3cebd629f375de3dca89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddd0fcd85e4e939db3cdd32d94c40b179655b79d2a0234b73491961f9b1294036dce8f13e1b6bd291f095cfaa12828b18414653203139985f44bab70b6e480a0311090c622658a7c25f6214d9c18b3d4b00639cf7bebab7f47a6aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebbef8da1f1bb53ff7fad22d0f1f812bd54c36511d194dbd349d436787fcbaaf7256d0672956ea15e3789db912a03b3b809541c2387d6055aaa61859b084782bcf5c6b24c5877d724de7232ab68d8cc2bdb7d5f2ee2d76b192c561;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43a38b8e923bf6d2d8eaefa3488a12797b1304ff0a3cd48eb5a442dc1903d7620391eca87d091338c2de2c7ffb20390082314bf3400ec484a5d5303dbfa8ec292007e2ac042b3907d63784999b0fb541068dec6bf0b8ad18c2d886;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13564eef2181cff79eeeb91d0c1f0d6611e67f034eb116f56d3c914f4dc533e4eca59e82cc8c05db14e963becfb483a271d06e34b9f4f96d76405cebab62de5b0deda814aaf78052473f527287975b4fd0f468f0fba1275b42c6052;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2f8260fb6ae84e1b13ca156b80e2c48743c6dcf7c07a123eaf6144504787102297d3bd693b86dba32a19cfe945c3af45af56f957fe8d42ff6103a9f515fd97612b591a774cf4af86cd1a0a07ac2cf4196cc11bb1a7574aa908c06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d67c985a484c4927b46e2c92e947bcc7a960607c07ca6496e078de4f9c70803fe289e454340291af68ebc251b60a25e553b3ff442082e84788f696ce042f17d6d7ead5affbb219f530294020849687811b04fb1cc31ebe2e33d24c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d253922fe553a53f5e18b1d3ce95af541bfa7a3d8abecfac565088f5432a19d05acc77dff89244c39a5450188cfe0f679df9221be3a39874b0ff224dee75e35578d6899c64359181b4142f8f85861a63b48e6d368fdd4180522508;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63e78d38f986a2b53427356c5d70040cd691a2ea137e4419cb0514ca21e355cabcbad6f3a09e5babdc4e617566163bb24f4039ef86ce6bced19fdf370ef53b506d23bedee1cc4cfeecea28b4ccea578792c9ed3f583e01bf2cd4a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c08d2e7726c7732fe7dd16921c38313a49ad0421c712a913d8de58b38abf9a88f14d7933b729ce9bffe6137dea520662300adba2714fbbbdc10d41d3f49ae7e243758c01a9771a73454e725211a83c635218ab88cfa6df861d02b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc2f68ec7ee1b6ad33ec8fddcc81ef71092ef3d85ff7481a4f55e50fd204ea734e9d7a7da11afcd91de9452dc518dcb1fa5c664cc5d7d8d4a3744a9254eed1e45cf5aaaa49b876713cd35401f5c7992ea66c15578a8194812424dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1168a9ff1fa1c11faeed94f21d3f3e74f9949c44b1839652385e153cf3a513f99ba52066e73594ccf9cc2d2cee3b8bf8c7f7a4ffaabde627ffc263969fabfe311294b443e4460f1feed2920f94772b644ac76307be81e067ad711da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc152e609d45f9187fe0e4da8553707824f721304e149079ae35176189a2af992f283b74e9ebfd6b0448cbddca28e74aa25929aeb8fdfc1673045519d3ac14020c7768d8a524b4341f2ad7154196222a0eac9c9c82bcfb27ba729a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50bce19bc8440b5e794bcd9b8e5c0f61a94322165d6002773b8e492544e00dde25cbdd437df8c69785ab4f711aa4e93daff9824290ecf045ac631091ae0c8a9f551cd832870254889434fc92baa681593eaaac6abc9984df13d6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1512218792ff50f301849d1c541f54e042d1e96eabea27766369a40d2103831e8ab5a7e6216a3bde9769fd00546f25723168b8602684f9c51ad8b077f88e1b9cb7c52f3e66e0cee90d1ecd8a1c394fcc81e9347068e3c8382974d6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c985ae01316b8a3375fe98d405e4edf7fac09825786a514670920a177c54b6610af2b3ca4093589611f4e5f272ea83946311895780275dabbb8f7b59b33b7415af6252657cab0faf3292b6f5988884646f1bd21b285c2a6b4fa93b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c5c2c4aabb11b5c971a8979c773836f71af0a377fdac6343557a3bee8c0acc1dd0cb39e2bc51dd0bc428e8a06bb067b138b269b207e84b46b162fc85b77f6265f682e7a42b90c1be45f717a0cde7f10bacb9d6cba830e5eed0bcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b698dd99b6812f480ff473fa7ffd310163a2cfe7ddb5529cfb5dc02fab345b37059b8a909a469f3181e0a951097a76dd4fbe114afb84de5498b6d47dbf8d93f7017ffbf3857b73efa473d8225aa1e16a2519cbac8fd7ab2f8901d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c628294ab21f774c839a48f9fa95eb392e38076b6f45a484a344f1c43f94c6f4d53e26131ac4264bdeac6c9a37561f91016c664aa15b8699d96631947734134e6f0781db58eb8db8b3e8ca0dedc53b467f333e9b9fc96557be0a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a35d3c29a4f0c176cab3f6d75cece9b04bab6d800eeed37825ab9e0959c3fc6a11835fbf8775e667bd8be483c96e2f3e7a97b5e0399c6869765139b2830ba3ff94bfe11b4fdd2e0a8596f5d714f7edefd9e2ae5e44a9701a29210;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15306913229e58332670e6e1b2a4891873424c5a92cc30f819cb0468b72edd234cd183fdf28b9d82938560cd82b683f207ef34395ed9a645b85f724ce9579e971a3c14fd11e5c8e2f73ebfae4604a455a59fa0b376f515146c29dff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he299221ea664c80133a576cb0d6b4c625c961d89f2208bd454ce5e79bf9f8247c40b706991d7be96a0662eaa6483db1fdc22cc867514f60efe508c9828a8f52f56b8f272ba6d2cc981bfa56fcd06388793d97c7fd042d90fdbfd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1051eb119e39db7c290c3f00764713ec281db9bd0e376451506e84fc02b7728b350ac261e51015b13d0e21a326d37232c2eaa42211d8ac5c272ca96c46c03e9c52268a299cd12d7cdb1644aced15432a99ff22aab9b741bedcb4046;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2ebc3f97959ba3a6ef67b7f5fdb6a58fe9430331e032461c031ba6a773113802a6e91df3aff67f70b371b01c8460c3342079f84da5bd6c05cb5ef92c0b6cc9a2b515241a71cbecfce3e29b8e69f11cdd0e54b18d67a85d7e662eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc5b59e97c69265579488c6489734cf3681339d3061e9877f2b4c69e3bff2ff54b31884f020e780085f4080c499818a45d3f9918b9bf983aed78bebb10f120edb55c843907e2aa6380266892c97e509a9d1a36f9e729ee90a2634f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h150a0b3ee4c5813240bb1fbfc540cdd869a3ebe7093dd7bdd2e3d8701411fe0338d7d8e1c513250bfe50fe31a446e0cc76c12874f552fcbe5612b357a928923215a13590bee70c65178d8fcca4afa21eeb59d319ccdaf5c2f22a82d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f7753a55353c0c0684ad05dc43848065df064a440018438617c5e88084fd8a334d2017b0876b983985e22d201286134eb314c8292626371bdab89fcd834058c5d7d766d9e8b5d8f0496a77a4770ad53994ea03b6e23b0a33f047f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c302359ab3e5ac2520c78fa1c6ef6d316b2cd0ed8ed1cdc05e6edb02fe2f9356979b364a8a89855fa9dcc7c56419cf8ab98d221ff44611c7d84230dcd6e860aae9698bb030f57f864c1ff03c62188fec0321bfb67dda5977bada92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h515dd6ffd0f722949a6053a3e7e08ec1e145da089371cba5122bcc0cba80d9bf77b15bc067844ac6ca4a5d0b32d734e471f75ca714668ffa1a45cb81dc7d059dbe5ba1a13a35bdaeaeb0439aff867353679728c1b7fc3b9b3d5eab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c349f91ee6707828279c69dc7a24f0c00c71cca5e3e08f8f863c8a4b233270072230410b3f3d150be3fcc1d04e25fb53ce1f6278f3ff43c144d47e9dd8c33f9beff53a5b1fb0bfd4a8283584650b33524e51d04a2023b80531cc80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf239ae6fd1fc868b5626f2e4844eb61ae2899c237687b73a46b4ee4e8612830ed4d7f17eb2f0c0d11b4b695924169af9e129d398310260f7e079ab9324b7d65c3d9e4e8246c2044e1e21da180aa7221303840581db5a708a77f3c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19526a177bfbbe1d5b02b08614212362dc90733837db36699b1ed199faa6a1c6916a72c03a3dc9b26440d022548781322d5496d8a14fc2471b37ffbb32a0e52e93cf3d45b8be083b19deccdd3669258e95aaa5e31ea98ba2d7c5728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1372aae1a62d2ff00dabdfe94f4fb7515577ac981be479ffea313bdfa793c95776288604402a60123133348cf2d33c7089cd695b36a97bf48d284f6a5468ba6be880f76bf67d2320d1ad0aa5ae96f7e715e1763a36f892705f9d1f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fab72d8f859f17594dd35526eb4b5701804f7ce262490d8e6c74b8d228153f4a8cd2c1110bba411bc553fa6b3b9b24f44b6268a1c1e85a3553105419adc52e7208f05a4d20ffd4bc0c003c02bbb6446d47f92f2cef195cf660b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85137e5fd01ae0788b10c561bf9af3b1213569daf83d0a1e727db8158ff59148afb84a71360cc3533335677a9084a12c355c0d72ee95d81cd98d1c93b868256463e7d7c6e54a4599fcd90c07571f1802d4e36d1b6a4f491b23cff2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79e69f50ab6fa4ebe140f4aad68108d734b20568f86753760e51749cbb184bab36039c094e336cd21a0fc723c396d57976da9e5d11cce6704e761219bababd84f0af228a79de417a575c07851e0c01a670cea3f4c08ef62693c9ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47514b69a5e49081f7e86a4a57695dd670048e4d8be2da1d68936900af8955af62d6bbd56f866c84925495bc448252d42927110abf6a3736c53f98c13b1c907d55346438f29e359b7e54a11454642390200bced0d790b060c6228f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1787086b15036301e143538f7e978ed8e3458ffa8e28ba1924b9513891fb67a710522c2564ed4e6be356a33ecfc82d222de20dd48ebd5e4c112fc55fe474450c7540977c6fcd77d80ced9c22edb0b581ab16a191c5f164eee80f84f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h222dad78e95b1bc3b32b878b3cf286882f1696c04472782b61c4c715d1634288a540b84da23b39601687581819b6a4e26b6198a78b84cdd8120847c3f6622f871e7e788330a2527659e53320d34cdd9e9a81f13ae6cdba270472b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19932071c76e582d615e4826f2ba34176209b1a76e68c2b74fd2d01edf8d347c8a9943da07b42635e2bc330d8b5ed1879106b49352f77b318efac268f6434db6eb04ee42142598c19403d58f0fb72497cdbefeb74fd8a0f9d6fbd34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137f943fdec740fd46c0ab2387730dc18f61803c4ddec8836086b39f0489ef6681d53c386361052baa33cc9b1faf5eeb3f4d77ab42a339bad4ea28f7057339c24cd8e86d22f286dfe0bc3fbbe38b12b041b4fea0542f43b2cc147d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162285d81ba742451c5c5ffff8d765c5dee5c34c174b05b789bcb85250dc3aedfc5101e2e968b3f63a087cae07b4e4be4db9ce817ea894dfc6026bbf4088e5a11ba95d192600e21103bf9f2706b8ba8ebeac3165c159c0c1200db5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14eebde3f7d5645df863d9b881d46264f33e9b9dfd4bb1881f67ece7654bcab8828bd39445b6913405f2b8dc5dfb9a2695178d60e3fadfd2e4ca7895ec9f0a9b46e413f28f7f36318a3617af278e7a1deb28d7b751b239d4691bbd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ee66b79aba26de38d8de7adebf05322a7bf164fdfca3b7e915878e6889b23bfbfe0e14e10ac7c37642597eb2adad5422db0f9a6ed48f8cb439ed3f89f921470e889eef1f9fef7bf5ab0d37a8f1c6106b47ace25a5b8b06b0349dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h774abad2eb157b8ac176682efb60f92b1b8c7fe44059d95f1e618fba17305fd73a9fcf797e1710490735150a2084c90a36793d4ed8d3e98f96cb1aa032519ad33a8ffef431fe595e77ee0e5b6a421feda67733c07ed07ffcf6f40b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caddd9f5f26d10f6b17c36798930ad16b6658ec3e4c60b9e98bf1735fdfbfd4eff97f6dcd308a0a1da3b1a0513cd87bd4b6a3ad28df365788cf9d2b8c37fe0b82ded15e8cd90b817c48f83d85aa4c6202f5df1bc60685af93b5382;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165038ef85c2804b550ea70b67aa2934a1e0426a21cd208c6fd541adc165d342b9fbf746bf8c1a070ea64d8d1129fb3cfae952e43ffd4b68e153a1fc371db9b2296f51fddd765198f480006dd87be6eaec5b9580dafdc2d293e5f27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176349ffb78be005681a26d7405378a1bbd5c809687f879960948f01e71871a1566e99719e7c8cc8e76f7c3b53220774e74fd87ecba15f1d9950232103ea873bf3ed5cf8e9cb60e237f8db5491eabed36072e3a7988c64a8e576201;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11560d8f0c160c182831e10298f7ef3801a1b9fc6c22db832b5e7ee9712a483df11ad868c5db9e84f97a0dccc0c012fb98c34b203b558088d3ca814f8420899cc5f1229ca0f47586620ac1f3ee33a130efd55d87f5e71f452a42f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15735877e7f4bf00bb896ef5f467135ef4f620c102a192960b1e071f650306103625a72b0bd02a93955354b7f17ca86e1c44ef9d4dbcc6b6c4b7c3686de0d85dabc9f5b978b793dc27436ad1ed0961c34a0a5d297d44252bceb51c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc13241aa153ad50edcaa1899a9c19e2c260d8a2022d47905c162813b670f9ec3d742615da057cd5d336c6f49105888d1e62804ed9b12497da6f58884f7c34700caefa547ae54a366d763d6bdd484e5a104b8f5bb0a228e22c876b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1e31ebafa5b0171b3efa443220c18e3dcf8ff90c41ee9a2b321a5b7902abc82c1eefc4c74feb5e76737d0ca5f5f25f6b0d61e401b5a10fd7248c36378ab2a9e1854dd90b85fcb8751b5cf8ef38b6d214fbc4497f86ce1d16a4720;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104aa81c15d5d2246020ecc8ec427722f46c4049d67d5c0eb8e1f9960127eb633cd9a0a87fff7a95cbf74f2074ce6be8c2705478464764380fedde7b31173f23cdd02974ba2bb2789905cd8ab407b6dcb8db1c3aa01054640fb31f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179d593756b2a02d3e0839c8ef0273b3e5633e4dcb8afdef4b60d2a679f2456e5eb3ed4891b7124a2fa218bfe21db4ab59f25c4cd7a0ad874055ccec28b9fc048750aaf020023f10bc9369b30057685328c02bca1d7f37f0c9f8f8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7750d601a204a5f080b7919458b2c85ca4132e0ebb8e21139099cb9329d6304e38cb0b354751595e2e148a90fdbf1baf67b8be55d1a308e5876a6e9d2f5a0144de2bef26a245cb753c621ea403addc1705fda70e37187c27938ffe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19540a23621cb759db09b85714f85354d9885f1aea2f85aea994eaa2408715b931ebd58a31751b2be693fbfbace39716cb1be3e99ec64ce1ffb5313a68573619ee1256121be084defa3f3911864e73065ca310e05626d2f9986a9bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab9f6e9cb05ed1965298efbc06541c4057e79714fdb05ec99b2839b783011ea299fb9c729fa930398734c37c83e7db5a1f2dac7265eeb75368015df2c16294e6da70c55ed938e4153a59d5c54905ca4afa16fcb200dc504374c911;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137488d8f7ef35d0bbddb86f81059998ed1b8935424ebd87d8d73e6b986e984a43bc9d5ae669fa51409e967fc0f0e5ee514ab25078c41be17de2846b8df97c73773eb3280588c203961561bc1d352650ba64587d26116718b809267;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h743343c4453720ac7883e14590de0d786265c14b745aaebbf0031000d69614de4cf13e40d8cb8ae56d66793934264c037de4eddb35b0d5fa024859ba657f121fb0278cd998cdc5d39301db5c18c4a4aa4c85e4276e6069d70389b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef3063775d294f171d86a2956a03a630bcf931a5031f03dd4d7a0cf90f93db334bbf38d5912b47e8ac238b5d5959133113297f05596434f6c1f71d24199f7bdc16f601e739b1ef09439ee7484712b912f993eff80bc3e91baea08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed18c1b9ba2b54dfae9542e35db5de0012152fc310252031ba179e60a8b7f7401d6d65a95fbebf6d1e7cd4e5bd58c0576025ae0d6d91d12d9eb8d65ba5b8964b16edd5e7df97aa4ea226a0dd28fdffdf3879841821fbce8de2d70f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdf548ff7f53e05b80759897f4c00466a41a71752c718c5204e17b4f83a41403a6ad05deb7bb117012749730126d05608667678012052a708b833889c5e8825ef1c9fc979ee8fdfb22f8d056e79172da3613a41d5626d9537ac4e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec64c23ade9726d173b3706f52b263830551519815c320382bb163cb6249fc436da8a4625eb853b616b9239ddc445c9565e38a45f497e7d4b050cc620fd946638381de0f9e4f15ac34e2f270f79fcb319a4c9960f42c74fbf2c926;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0805046f6f0b136fec2b159adb73313a5919ea3ac92412f0a9a88fa0a383148881bd048541fe2873954e853486fe2a0ec6c8b47b77137a058a57d059c82fd6491497e8549a8972ed8775d55c3f106cd05f345f8fa5122ca8f6aad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85407813ed45e2f5e3f811aac91fcad86dad37ff63b766e5e7a27a6cc145775fcac51b169ac6fb44e1dac68ddf60d9b637f30e910380aa35da68acc365a00f2a19e09366b4061f27336b167d7902074df858289b710b431180aec2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bd9a09ef99a0f002e38e7920da14a69fe3b19da3f8ec4dd084060255bdc8bb964d2a345adb815ea941cf75d1ec29dfe4df92164b77d63227adcba8be6d83a53a5d919890976bc5b0b77b39c9203b509b53e438a14030c2dd23f1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6553316afd1862e1ebbe6416a2892b04eb068340c4f925888b97c3bd9e616bedd9afbcd36591c800a556ea300721e9cdf25131ba516a1f94d8ec13034ba8f0fbacc70b5701862c8ada7f45c12b9cba24cc0ff3e367a0fec375c91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1081be91817aab073472be4642910ad67b30678e662558369a6f4cd4d24afff4a521b96b26aa73ee2b3d0afe533e881ecda423cb8bc653a31b907cc84e0e61e4bd3f4b5b03d64f7135f55f6b14381011db37e457090ac5b29b90264;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1515dbaff8b469eb0b38d8544d12332824fe2adc8c4f33be77510a6244486795819bff477cf1633303ff4de77a2c7441849ff1b82c6cc8142077152f244d33fa66ce958a2acc95ba3be74c3f614002b3e8dd0e052ccd75dfc402931;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd48e77e6e08469cfceb171790575a5d55f02a350e24e2631bd6f44e95c802cb887336e217faf72c2137dc3126768783b3cf7289c39f5ac7abba39018dc821a1a3dcae83b1b77ee25ca10a48d5e2c0ca44432deeb33baa667256e41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h824008d0f8c4890c6760a8498a3f4ffe54ff135613c18024bb9f61f2c966155823540d3d55a08df893d07614594677e0969b535078e01b48c337dd75633cb5f83c868e5c8a18349335b8bda603e31b6ceadfdd4ec04f6f1813ca26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a6fa9c0cc7d259d7516faa1f489e976a41b1e0024308992da7d39cebad3b3d31a2ddf299f0624fd677c8ddc3032a5af7ee4de73f4a7cf63d58d4a6b52d4f70fc0bfc24468ddeaef8cc81e6a4c09d180dab32f25d0f43c8edf01c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9cc64166b872038cd7fc8feff5c936a29bf3f0dc41cd991159ca67438a64f30d1777f90e781c2f630114d0f888b8029b49c039e977bedc0f49798af0c288c23d10046d1858909df9fbf09f2a2442626ecf0e038cf2c2818e2f858d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11dd44b3e7b251cfbe98070642098a1c908e6465a0639bd45c28d0c32f50373e01bb5be77f5ecf1c291cc7c4ee325cceb13f9cbefde949184bdf4c49102bad7efb738d1e9d38b66bfda73cac133d180ff2e61a3b6598de813a11658;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h720f07ddb2e1a268839a4e569d411cd27dfa6180152d82f7e8d0f094b2b8efb94d8d3a8fa3f5eb7686f027af06e2e45323c5f4a4d5b487ad4b3068f3991e7755d117c9dfd4a91ffbea83eb1b5cbcebabbc3b946a71d39d150aa1bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2443488be220c78aa91bb49fa16976eaaa928c127bad506008b41fbb185828f89bcbd292181b4a12e347368796df9ca96cc71f5ffdf3dea3ea23900f380a13980b86d9486fc8d2ec9f5b382d0d2214ea703e0ba08c1a3b29733f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0dd7d77d98268afa235cc433ca6f2bed7ec76e160faa105798c07e8b32d8558283011f7fd20c4941181bc73af7215cf7a173265e2dce5be72fd00a54830037a45d0b7f4dc88fcab823a7c31aa41b9cada30bd92e38f24112e4693;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebb58cc693f78cf7bdca4153709c96563fd5cedca4690802335292dc3b7a4ad9ec868f67030092bfc0b7d99a106d9d8158baeb1da46e9548a34270cd1d9c414efcccbfbcc8d6397a2f4db1ea0aac9754a21a453985e298555d4808;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c346f944856e3dff864b617336611e582d06d2258f7a32e482c7e72ae8e06827eb21018e4bd9ca92067a5421f400e0f2365f819c175b1655666474a3a105e7cec1a24a58ff2e09e2a7c746726c53974e1ea92d37d6eb946d1dadd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbfcc598e6336a681c16538da376fee627ddc1e98ca937f284911301d3e20c4c8d5196b90bc9cf647a54b780e3892aa4a9ff3d827d3ab9a19df7fa4a939e23906c746c8775f39ce2d691e37006e81a3e2ea304fe129b0f0930a49e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3bd97d13be35c1c10c0918d2b8a1e30dd44cb80d5ac0725f3d1e81f1bfc9d766f089bbad6896c0d1e844bea2aa141ee6acd98338e9d7367bf9983c04695bc474ed31ee9fff33524e4f1cc36fae79b3a5bb56a3730ab3d858bf09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5641cdd1a250ef259c55df0ecd82bedf62e60c36fb1d7f89f98847a86a01102162c643b0edc13a4584efebd29252069466faa43ab48b3ab999a8cb8b2c6f6f6593b05f614d5703b1f08af2c78cecb78d936525c2e690ec6458e48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78a1879d3326ed6319f8eb25d741f5342f1c4585c4cfe646a8c70fa622e8a16f30265b5fdc5d067d4a0f4d5a363e5d50f9f1a5c61d0726f90277161a3a1e6503b7f63e0cfec0899d08e5724498412e9ae1dc340e7add75a79c49e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63821bf729f21d11aeb09637b96824fedd1ef98343278b63d521275e14fec70d3ca4dfb9826901f057aac2cbb25adda3e53ff04c98b2a9c4b5fad0e106c331f630814f84e627b511f2fda78b6b0396b4fe44c511b9f48dd8e7a105;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114ee04a79fec97ea4f6e607c879ce45e655c811f6b281c3a23ffeae6b8ebb3f62cf91d693afc258118aec9573b85e2238f4adbf7fcf5d16d94ac5a63b9025dcf6f1f7af8a9a4b312c5402c0d22c860341c6cc7c4f35fb34155233f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h865491e3c1733f6872ab5ea6bb3303848ded55c1a68c1753c9c2abb9187428b9138e6def6f50c6ca7b7fa214fad177d295208ecc0d71eba224ffac5d433301d4ebd89d048a794ccfdd786134a6ffa1c5a2ac0ac1514b10cdd10d04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h456cb709a150b2d7bea97c5ff52dc3f8f0518b8b0ae797f92821289f4bafd2986daf91fab08ad1f2e4c8a70d17bf054a512d8cfbd651d63d928a7ac2a6fe6fc364c16bf3956ab94ef9f027f16d8734866e0586211562e824cfc195;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff1d3250a1ec5fac52d72a60f246c17a3c30b8c60b4269b52e8fa6ce1b00f20d5061e96b4dd60ae869e809fabd8514262bfe7dc45a3013209b56aa78b10f8c1b88668890e6532a2a8dc9d4b23462c1cb68d928aeedd9c77df3e116;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36a64938b9c9511f469b369216b605e6a7c07bdea2483d1b2fcaf5d1730b9a90cb342ac2f504bd80306cd0439fc0675fe9918611b707b29ee016de3fcaba477444531fd03cafece21362c09cbdca651da64e5afc92dfa925334888;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2ff9f6fcd510fa987fb4692001c94a3828a35efbeac8867587897ea52469872e0186b40136b9980b4d9468dd71524e78693c4123527a3ec6a45a543368d998d1f136ee62829d515043e3792166da382057a3dcc88faa5723a2a3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c085ad91d3255607a4240ad015b85ba051c1b00fe6d1a7bbe5dd49fa806c8974eb764c28829a202399669d28ccd6ec9c0208db563ac2e885bbcb71ffe6f00a84663c11a8fcc788c5e91bb6aa1ca61187dd8ed73f275d1b4b6fbdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc207d9b76eae4b87753177d755f187bdb17de35903d934dfe1387c22911868f12b95fd5cd46e271f64f9af3ebc6b76810cb170ed64af4ba915f422b53a50217b46befed25ea2d79888f1bfcb9a48c9296e6108b2aa2125c3db35a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a95f23c23b047ad0c51f8a0e8732ad02a4e999ed1333770ee6b13abd6ba9c17429373c6af504d15ac1ee368ea830e9f882db8b0b6f0182812b28777ae1b03b55c1092da7b7ca75be7b948d1f27bd0b1a5f8f422c5139a577ca303b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163cea7d265f62bdabebba3b47d97e81fd7059b2f39c42c013b52e14360746f83d123207a12d328bc4648e1ea5c377138ecd2120fc396d7ec783462fcda0f063812fe2d784303aac1189cc9168ea370a03aec3f0aaa63ead32feb97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc435754196e645fd8d5f2a5c17a1e86d56e848e787023ac90f0d19acecf51c4e85665b703b616d38b455e875225cbad407e0708e2dcfeaade7bf02bd3b2d2cae17d91b5986141a8a931614b7f8a01c0ecd4623c9930a6d72a1898;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d17dafad93f834217986b1ea1925fa913561f4dddf6f6afef5e348f946ac008d482d5827afcf0303f83d6d0372b7e6bd88c54248a9d1fb751bb293ad1c788b698a1eba2dfafa31af849892dedf93579ead7cce1f95560cdacfa86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1835fbf9ba1ecf567d4a26942a0018ed38329ab122f69b4f92c0699a7a4117a26a2b4b32b9a6759a814bffed2400785b2f6550666315ef5c659fb27a40d97df74016a48d883fb029e739ce5f4deb3f87fe91b088e8ec750e0f32cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129863102d60d5ddac7c8d7fb6f601b11fe48e94d0f2c275a33c85db5c9aabd010bed69710054f289608405dfe876c83f238652afe1b8f93d78f12d7fab672aef1ee5c20bba63569c0041db89d99f5070d5c483d2332c150cf84d07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1ef932a16e0d7b2db54ed6ba675ac6d1b0bf620dfda990f2c81abe2ccf19d248024332ac7367d0e684ce3b256b32babcb55f50c9e794f43f00b3ca5309217274017964fb8227465c7cc42563849921bf46569d7aabc5cbefd37d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155f881a839f1307878a96f2aca8687a1d8fefd7f169b67a16f69638c299200bf4e9aec36c5a7da68900f2e50efdd75fbcfcea86a1757dc7afccb3ca677b912826333d4d4a469e3f71f4704a11b0bcfddf8f653d90615d6d86b521e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf973f895677d3ef03d478e26a707d2e07400b23e8449d4b0626dfb686b9c19bf62c9f8c9d8d3d4e4d999fea55630f6f443d7158f7129101221ffec1eb53fa534a54343b09c495c36c462bb07267fbaa715d38c48143c970379481e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d137637a38adbb5f732077c1cac6c09a13237a9e1488263353a0c1a870d1c5771880d34609e04f6c321a6a915088f063b1e5e7ce251344e4183a9e0a9ac79df9790d1a9769a2b6419c41e49d10499e0c7a0bed3ee3d45eb0aa226;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ca350222ef4fabd4e24c795d1f4b6bb8bfc3df517372b4b9994889c1f71ee204026f4d285db2a1c90f4b8fb229b945d168e47f8d58f10dfc01f0147e2cb7d3b13698537b78d865d351a36ff083dd824b7cabb907c81467f20cb57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hced60f763fb91f5b6dd08bfe74ef3b5d4d092427a06d7bb554510269dd5ceaff15f678d542fbd4d03458f3d45ce2e9b31f12665376bb51d6552823f7ec8e18766678855fd6ec32845daea3c4986b544d2f0b32214e1296e47a0409;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d8707403fef2d6042603b92ce44deabbd08988092fc3748ae7ff2cb8a7ac296dabf83502cd459a6bed4d301f4c17a1c751f3713c8fbbd42d393b82c2926396f4e389c545279693d1e1e48d3a8f14eca02bf5a427f0fc55477e30d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114c9f47707f8110a3a77411e2ca3e23314bee9d2fb04d4679b6fdd9c9edd414392c7493349f8da5476c55244ac6f72639ebf00ea23deca397b1cbbbfc1fc65b0d92796078bc2d165e3383805a402d2d926927fc2dc9dea84663032;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea73a41abae7b9faadf9244315af6959bd55459fecc89b1a3f1b689f096880a4437f0157a5ac3e9d7357212385f5ac31626123f498019344f55dd245c1c5cf26a934a580b40d8acc90a51bab86b1327fecc100c537bcabee777e58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3dee472bdfe0a6dcff0134f08b9ecd23280613fb9ea09f18759ac1fa8f8270c58649d31cf532b8110b863640eeed21f937e98962ebca64fa8e37b5d6631cefc9e99297ffb2c5282347b498b72daf0e00edf9c422018bfa0900d26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b320e58d2e230cd883b42a6e8f4f659350d216385754feb388ded9f9402d81c818c3bf88a0f9aed80af25021c6510e8a25e4458fbb6b408fb7b5cbd9841d4afb3ac1e9e94afda862261c25afc15ab8008de7be5861019795f28a05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf98542d806e9e03bcab51c096b122e355b09515c3f3b8d91a1002402cf111208272962d29ee2ca0c1ed687c80d58edd971a266c84a9fbdaf62793b53571d60932e09894cde49284bca3a0045a314d4b769b9fa0e579080147de1e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129b00f83faa8dd5d9d18dd0cd7856c2efaabb8fe83bad913fe026b3a9207cd5e4e16d285e6eebff3d213e0d7f836b8a28ffb2eae3498d9a70827b98c4ff9ae784ad9f7d9f42c22afc28d236f4be28c435b91be238aaf8a0e6373b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb8f41aea2eacc8fd97cbeb491d4ec323b3ee5ee1f33d303d6a2e95e86b1c4e209912aaaac90d841586dfc85294ad294673e19c1fb9ba9f23b444e834c75ae6e39deee7fcd4aa5fbc26d212482d4456088a633e90157c1e26d0b58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b7873b335b3c1e4d796da1df59704c323efb1cf6cb9860c67c4c51673310104eaa8bf5cf2f9a2acb507be892cc64d7997a4c5e42ce0e8f6f2b797ab371475a0348baa28e57b38b46c25b63a02c080f1eef92386ec1b2f52b9a602;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa01a67e55065e66471a691790f7206ee2abcbd004c47a9a642a4f4155f452eecc960a7d5a99141f7ff49f44449e261585922c86ce4ec5bf5832c07ba8c6239401f8d0478314f79ac58f6c0ddb0be50b3739e1757b0699ae422d3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h679e96f90661af0d4d16678a1bcff4fa7cc621a0e3fbc0d44ade4d831bd0bcfbb1d47693b23c2e7c82f75646dd3b61b3b9a8a882de3b3171c9ee638ae1dfa927094db8ef384d2e6f98e9e5337b3a4a4ac9c857f658810b7fb9ab3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4542d03e35d5eb37d5524800fc3ae3594642a904fc0a769c84c25acba451f8071941a830be670fcd865e90c183d9db639823c1fd4439c8dad52e941205a47573a9bf1aadd9fa86210fb449e4748af25ac272af3ca13f7d90353e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d58b688e2a9d0ca5c94bd6c38fb7d60786b1a738f96e3c45dcaa0a545f02bc44ca909f877c99dd2e6d26d49be5320a6aab18570fd20fdd0ed123c4a5341786e446a99b8a2d1f708bed95a7f67f8e2a35e1798b39f0e7ebf8ff516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d77a95c619671efe89cc10233045bb2fc40a3ed1487ccdb0f61522a9f209ddb63dee8f59fdb6a939b83881315cc426810d18c7f972b02fab63fc984f2a108b3c3f022636e63e207e499e0d445c3b85bc4028ece50d6b5a628ff45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb82b8ed39adb1d91505a5cd6130d1896587239e2343be957b88bc8b8cc8ec76d3988997b18d3be4594bc7f48d141350514a664427d80c9ec4b9b8ca0a4ac75acd42cab56514d0d9f487ec660e68a5ff19a41a5c23f29f8348566a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9886d5c929fe87149d61db5909a98b99e84533915becc07c97a271fcbb96b24b0ddddd412d791a9d1a535d2a7b4a08bd41b9715114772de0a4dba62d752d89461ef883365834c65a38742bb38bf1b31e1dcb764cddb40f930c5f60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86e148a4314e522d316e51a49fa00712a41fa8ff01d34bfd0dcfb05afb3cd5582a040bec4de57ef3fe2f9a5b3cb12077c9a9f3766849fc431168a99ef5ecdfc5e4b5d1770f1f8f30f7c9e989ca5726b1221d6883a50d9a3f71def0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f9580585520c8b6d36ff8f8c131f656509da9eaad9443daea918a04050f3af5c00bf929b89b0f34881db975f54b52c58cfa5451b0cd7de34df2f5cac297686d18f1b524dcba0870a38bd1a9611fd5cf7681908f63069ca40a27b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcab30dd7ef975694e35ccf515b583a2be2a2721355a3145d83109163a013466043df3035ce7cb500eba583d05b42c1b2a3249fee39b9bdf4b2cbd0f61ea2c591c91d1f108d23ad0fde12c50ddcd9da41c34f065d498a0fadccdd09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7b05092a658a1ad2214454b97c836b8c78a5903bac074a84f247c35e3c2475601d3e57faf9222a3e9fdea4ee0a793826ae971343b4d142de90142dcf5a63a32206dd559b5b21e926a28e5b4c4a774c540d77eda96d2c5eb9cabcc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9b1cf3d5e0a260e27ec75cf5489349068c9eacd352484a78a51df940d23704a11ab7ecf7c2e8dfe8a47c34578d64e77f7042537a5765054c48f4c3f4ffc85c62ff035c41f83819982995ceeeef364a93ff355c4d150a688d49ec7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a60071b2007076401dc44ba10e38eca94e9615dd3055e3b59d6fc15234a697f74ea2bd7f76d6e847e2a10f21a9d53ee4e745f7b4308c72b93932461db0b014c1ae66f19246287222dab094692880acac73038a583a53d5dcbcbbf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbb9311a36feafee662aa0b01e252908dfce2490f6ab0d7edf8de9ff7400757d4c99a308c68870e04592f9549aa8eb0c803c2a7b611b3e2d4d12b5847b179308cb52d2babebbca42163aac774be983307a8d1e64a9dc427a4986cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ec838e40e05c7dc4aa918cd321a50fb6c815de2fad2cf5ed7437d59a59faa82125e6c38b0ad8354b1950dbf4eb7ba2785adc5aae85f5f0f9aa0582d620cf6e750c14e00dea92703913dd40c48eb5fa0910e4396e6d1f60fc2cb54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d79ecff2835fc94b46d182dac1c7e5220773717fd8f891036762b788d3cbd45523876fb53b8415f5fca0676ededa32c2ff505ea039000bf3a962b252fd4bccef7fd9ca3365ac8b85ff5d0642e31cd3c122dbdd8cbec1d24c8a4cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19777b5cb945ef7306551a7fc9d04ac15c45f58740e6b7533d1f0f3f361bb5da3c5c345f23781bf9ea7a14d53cd2f171efd09bd7cdbd643784c06b498b53c66fb9d3b28019b272eb93d0318549d74f54d334139c697d2de469f09aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9eddbdf2ac50110a21a0fa525a268c1406562b465b409b79f6052e99f57fbaa8f6ec183b279871677eff1b167e7e772c44eb201fd3fcc6805d1e10e7a0677499cb351e955d459dae0bb7301df3656ff4baf40e5608b1e49706ad85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bf24e3c38ff4966fa4b032939f63ee3bc741eb995ef74aa8a081e6358b6f8998b62ad047ef1b92b8d3d5691e04bba9ae9ed14aa6c0704d909b61a762bd16c302c457c1c137e99f046671e21402cafd80427334b1c3162bc4e49a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f6e7d9c736d4b24c487a9c01b36f8df75fd1ea43e50743d4f276c1e89063789df8dc8073a3bbe54cd6bdd452218eb77b7f5e5b0f0c82983ab3f0cfa618b069f8ac5e9266187e960f54257a1e991fc0932e978393c666f7627616d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae9f092537af06033ac772d3e4978a346a1672ef711959faf289d44fd82a603f3281ca28218aef94572a2e4b211f3ff4991e84599ab2d509a0aa66e96ee9dff6fa50e91592cd2e3cd1af87d2fb2ed6db9df352e26d43664c78d095;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28ebba0d43b5fefa907238977602c76c6b84aef3a19c62099d8c88cac14bdf020eb0418bbbd07f61a80e7b16a446f8dfed9a1858221d3a29edc32a1b01741353bd0bdc83ec7da41fe875a699951d53c2a2419c821922e175a60243;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5722894c21c05c91ed8eca38f6f1f613e0121b490026e564cfff01821f7aa2279cc85fd8da4f6acdaf60b6719cbc5c55d15c588f45721ff734cfd4640a10b79ecc3f30dee540c72207fa8cd50403fac128aaa16650522be7366d0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd10e0a199375b8641d6820666aa34672646d0ee23a98e7e06755353b5fce8b4b24d5e4c593ae53ca9a8e39871d2a72e3192263b3b57f9505cdca6b9a816df134210e83666658c31f3e2905af41cbc9944ec7b3008820ddb5a95c80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157d5861472eaf58adb918d44a413711a3a086e466f9568f1de3217cdfb7721440615d8738b23e1b212eabe171b796b319878e5d9272884fbf3925285f7c4e2284c2ae82bc848727d194be42d189e0f3097709e44869697f4f75fc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he67a6d00d5892efd9e5f4838ede6a92443e95e34bc5d73c6771b59051a242a8dd4d7ae52edfc0cf9fac024354a1f5a1d66443b4cc63cfe21aa71b4cb2425a9d83369507b313fa14ab500c9ffac843e2fc0cd46760185d2d6f07f00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6df655a90cda7fe35b100bdf69f4788dae75926980ba6c8327d9520788de99c0b5b8ac57fa87e79dec57784bfbc1bc1019f71cd8f23d9c7da8f84a3db0faeec606a3b39083ee86a005497bc0d71ab054c0c0e99f3816275a31ad52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed68db0b9450597ebb4ee2fa12bf152035d1d3f6cbc0c8eb8c88bb7a824f13e35d2349d585e2e89b2bfb6ec8c1bf3b229f74688eafcd93b6335e903694872db78c9f460281e399e689712473f45c4a7c39c536b35ff7711340efb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ad6cba764cf289c899d8b57975d64b82e33f824a21a86fb33c3543249d62f9b19893f103bbfaaf0273f91d28922792bf6157923c25170a6501531dac5970618a4ee89db2cfebe57429975d37dcf1cb659d5887d6b7d869fa35b5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he709724a8c1396b3af6a43a1404e900127cb628adf2ddf39beae930c5e5dd5e6c17ce52442b2a5c4159eb1ad360e11171245aada718d5c5c30d7d16b950882b6ce471f1eb49a8f3cd9e23e36eb302896edec65245b88073a5078ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8dc27366ef3d2118b75b354ae3357c4ccb636e530d55eda3a1e278684109e1a8074e626d2c02ac9d1a70dc01e1d14836f3f64ad82a962d4ac88feaa7bbb26c6a6f89bbf8fefb6159dabbbae3789b994bed5b382937880a0636c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e8ae348de9482d3373cc2dd555a4cd6ebfabe39981630c0be4f3f81bbf15079b0f9893707e342dee50d1ee02f6e591dd1af45e50358d4ac59bcd5c596d2cd34248cd9870ff4faebfac30d581a229b3cea64873d1820a404c5ff46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1769ea75e6a0a3d09f1c35eda6aa23484418f13a67fbf6d842d09a4ef20a608e427eda1a9e577669d47310fd7d8ecd3626e7fa9f685fe0c912b5e9f7917fc048aea4db99f86d62bc06801ef37085057c5a3083687261115888c29cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155dc4b26491c70560cc6726303b4fc8bd28e9144bb9d73d608810edc1191ae31f2e884489bc4a249482efa407b2e9c6e2e7d0d61d8be026b23401b2a6991dd9436499658b7967301df63237773f413c5eb2beb800765774aebd8db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87cc1c68ef907297fecd8d985681145cab9448dc8e6e1f86c729f677dfe18199d4f540a8789f08c499148a80469cac159a4b326333112430b771ae38aad1518e206aeb7a6bc6c0562546eabfd2d18ed62bd18d9882d4b86eb0a565;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0377c3b1f5d08bbaa18e55890f4729fb3ddb4f9ab7a7b310402401e3ea746ef245d2575467834120f6568f7bb395154c60df8d643037beb018f2fdea903c48c1b06411680a51842ff53e9d59e8a989739afa5992115764ecec35c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3865e5bf3dadb4088ed7fe04ed7a4c8b042cf3653dfcb10ad81ccb800ed4fa1c1a64337b7492ad85816db9573496d6f017d4f9740fc86b33fb07329e4a198d6d31a24fde3d1af14f40c9976563222c6c96817c17b57c7cd6b946a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c3e1658fccf9ca166367e3f8dd78159d8a7d6f2a9fd0dfcf8817f4fda399f50e1d6b47c664c12c1bb5e0726a52cd1628182bece1c78902741605a606d4bd2d93162d0ab6acf2f0510ff5910f9e48c08fe5afb237db75c47daf8ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff06b1c24ddae20a2256cee729defe2e244b6ab74ab2ca2b7d32c1995595949b797766b853916b0a46a45c956f35230e03599eba8a2d932084a65c79557318958dfeac57782adf6b6a25b1bb27e3724fc7be5a1271bdc7d9f339f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1047592b8458681511f30f5126158ee58438cf7a53fe9a3a0cff2ec88f50ceca9d72787fe24ea67ef67018d24ba7b6533ab35e788945419ffccb58f97bc92a49211fd4a58ac192ce75e651b9e58185c3ae1ad8de519e133f8f6a949;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98917808e4f1414a99d864563f0fc34b1b95801a33b91dc10ea998b4bf22438f7082238409e6ea024487390ddf7cc10ceab62659ae44e375ab3f4352540f42a742615400ba8d1a3645ff3598aed40aa8427ab59144c7091027b358;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb13fb733c1003097f5b858318364b58833b34f49ee50e289ccd6513b0775f91887f5298910b6745655bd8fed8b338c9b355bd97bf40ccb2cb1c7184a741fa93de0cea2120143ecb674b5ea996665b6b8070a76c53aa5dff55f0ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e69adb05a14c7703084e1a450496251bad1ff6508b80243d6154ccb11181f7b6d122fcf73b82682d618f8a30a46f426b4a05d97661b091d4915634ac0df5c5d8601deaefe9ad10d32601ab5a23e6c29715966ed6288b3e7a465914;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf4a7ca70bcdbaec5671ad4a148bdcdc29cb19dc9d5d5fa6998d1d301c0a19a5b5af0a39c3e49b7d9d15ca581eb414335be7e8f3fc5d800dc4273119280986ae635bc2a00af9b1ecb162712ed8c96d9d72eeb7d7cd21f6251c8f56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14433e5d4f94c2937dc4dc5639f0173ec33dca4048afb31276506491db60fd631e8b4d30185f675a7daba4aef4fa91a5b7f72f6ee7606ed30b138ee485e92ba38ce6cd679e3afee3648373a162cce19316064ddbe62c99dbdeb291d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h756da9ef0e49dba6ddeeb4b213f5985e03b2a82665993ab69237c3dd60f2ff5ecd38af570508c33405cd984776df900912e866b473c72e4f6a5e576a7d32bdb0b3a07c73c4555a571525f9e21c62dd65f46ac78f7e77c995bad2da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h543e0d5591a587d28bc91cdc26363e7bbebc2c02b077ea8e6d7b6a06d033abe0970311ffcc923991d9904f4dd6d3365e695639d3bd174445a27a22ef0d89bd0c5257d43da19a8c61fcf1a42a00dda6b368389545ad6ebda140237d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he590bf37f6075f5b3bfc678fa727ad8dff087d444f4d5e5f2fd7de31667d7d70453f2a7e69bd062c44f3f7ae4b880a5d0d700bc65d01074004517556a89f3055a7c6ba3d74453cb87f647c495f2dd62a91bb9939b411ae1c5967bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105bf165ecd1c14e6419a5965f8f133288f0c461fcf8b5f4d056d15c89e9e39544595ef1f2dc21dcec5e98022412790bffead5ee3c4f14bd52285672770f805d27fd5d37a024a8fb1fa4760059eb4c40d7a0f4ed5184187d041abd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6c5d6fb798c97af47943c2173eb6a8c11ea7061ff96647a862d64715a1b2d505dab40ee8ffc212a554e80a11288d26d8f48bb6fb66168d529487aba25de71f4df117073388aa87bc9add61f267e7d1fb530a35b787215c9e429c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151b95e429f2e9c5ead47d6bbb28d264e4b3ddca0be85c4d65789669415af552d41128b10eae8cbc6f1d65f93cebde4636917e50324dbb95c676d3a3b7e5b22731c8bcbf928c9cc79abe5818dca8fff6c40754b4fb30d307301403f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175a390e30ac5f792d4fccd1d1253f164d9b704f620618136c97b4b9c1af885aff0005fb552ecb6cdbbe342fb37dc5fc80836b2a14239a41d88de5883b69bf217fa4f10c6dc452349f932202918e274d4efa1b7b0cc1ad61e03f151;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a5298b569dabc3304f27ef17a093f4112d19532ffd0b01da90e0daebc230f8639b57a4b4972767e5583913a4d459d1939a5ef6064c054899b233e9008455296ff037fca056befd416e973fa648df496f16433272ef3717710b9b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1946eaea688e5c79609d674a3c46178bc3f9d6fd866d3584cd0b6ec8fdb180849b3f91eb1ec0c311f4d9ffc2850c5260d573a393a0eb9648e14d36fe4cd0e18fab3cadcfda767378bab23c1c96a53bf235ca952af3654210a76c957;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69ccf38fdd4d3af4b52057a88abb9ef5fb05f805edd7aba2b574318195c061694733fd4aa5de738af3690a18cd89d5f837a6330b627c404ca6d82e1ab642fe38843a98eea1755107f3f4c617ee4c53de593d8d0f838dfa0d6c98a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1647b17ff54d74bf7058826c46a65c35dab87d92b1b59c66fd5d1fd939b7c941454c763fed88cf70a7200bf148d2667c209f9d86852777c1bbc20b3595a8786e5eeaae1936aa43fe85d2e2564825d7f83070e38e83f5312b86538;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2996548ccbd424d40727632f04a4dc66da334264e75b3148aab690613f07f25f5f9507c7302dd8995c48495f3c885a6a9c84a158bbf8a25e7984274394132cccff019b3b0fc69bf3586c7ea5294baa69421569d446ebf8f3a40bde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e5bdb024b490b63239ed748c4eb28d201537625a21e8092e6cdb6a8e0d152d024d0883c9e73b18196189ed16cae118333ec54d8e41c69d4fc4a155decd62d602f5ea415bd85f65178a0331be4d61b58c793f6d2cd291ef26e9c14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdff6fb9e14af38bb08a231c1de9502dbe1866f55a0759299fe3d2c88ac94af4b07d016319800343a922077d2db932a74c74c13e10f1de63329dc387c3de5930a33f64a847e4a971943b0858c899c06dd1c5cf180b40b29f3ce6bf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b43b3f1882589f7174cc07a8d35c34f9cdca168845e23fd2ad99c4e6d159468bf8ddbc82ace86f68a74605e335c8f613182eb66f91005641c19229433093fb5c680ab3dd8928694c4d0cac89ad59ac72ae47310668262ec822a25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16931073456ec1cab2ecbdafe946ce3d6a89d9bb39405bb4cb1f7779c4e5769b2c7381c7c4a2cc621c6792b087885a7ebbceda7df113698a078ae667e1d02b766cbc8a49db1f9a5f9fea1c28880a40fdb20314c02db21dc42bf8ad7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he73b765784699d7406f08eae269d4b5e4500535152a9ea63719fcd94681d7b9957e80ee91a1a69461c75ec4102ab081dd83dd2fa85bb0c147a5e9019941eea9d84c3f1f189dff09137606a9b6533f86f5f58a2af57137d45fabadb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd703324ca3a37dd7c20ec433d487dd1817a824c2fc1244ae193fdb830a41c0e8e8e8286e9b5fb4d93c067eec9fc9e9783297258d9f83e02fe09b27d929126e948e145e3e0db1a030856e1f7e1f1c8a3ed3126f8e3ffde52bf3381;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5d6dcfafdab097620ed458ba7ca7491d3dc91d667c891fbabc1983bc62482933b7ba48d9061af92cc26da7167cc4b58b726086f57a0d531a2effa7e606841fad7cd234cb03e7180521e12420a2efb57643d990d5611b252ce6ee9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf61562cf6c316106f277421cc56744211daf2814ca35ad1011d39b289298cfc9313e509d2fb4c5615aac3d4b8582385ba44f1566cf1eba8746b4f0d55a63853ab29cafcae42b7a56d0a89e4c175d1b319a6eac01e36d157b35c6f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10755bb3f18ed5bcf2598d00dc39f8932b2192fabd14bc92a61982316637f50b8fc1cdf51f534d0e849811787e28b3a9e471fc0f8cd75e4f1042d5d739e1c7be5e69d92dd9b1135ce5c6d82f7b4c5b4efe2f118bd4461e6dfbf337b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bff23f21ac21eca0bd69bae3da985eaa969fc49ef21941b83d4762712e75e08ad6ff366d9beb79b10a70f0aca1389024277f64af1d9b842accdd797f7bdf69cdb31cbd57aadbc8a0089eacaa30c594da2573829d675bdc44e11d3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130a52141f96c07d5faccd971f13fde4a72bbb239556f7c3ef69aa0791d676b5533175c77171599632811eb2fe7d1a3a980e93bbcb8cae16243381be50a45dbc843354d6b65d3c16bfaf2b8090be775a2fc926e9d47929e9fef5c38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9c5a4453137d541a1fdfcd023ec1d651f3bd4bb27a0e5a8c1c4c9e21a36ce826394511fbdc8f1d57c8ddb86801268d4d1628c915d7f3073041c94c49dcd7a8340087121b6498008ab44dc6ba3799594fa87a313b104b5e1b3ab77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c122611326855a3b838bccefef9afc00b9b6080e1e6b8290764a13bdf1d7df4c58fd9f9020c50ea0941c3633bbba6e06191994b456e31120f8e67905189a939ba2a1d8419633b8ee875d95f08718c19696f2cc7075540274720cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42cdd4ac9629aa797e9f56dde530053232ff6ea5e35b4f189172630f51ceaafb9fa55d4efe7af09a9175f0582dee59206845671367e21e9889ad1a440013a18a93b1d18fd32ec5bf1463175538d31d7563a8360b3a73105dc5e0fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19598a57aa6d9005d9ea35c83bfd394e527c49a196203696ac505652e2d17c33f5d4b02359471e70fb5eb611bed3d14290928d86b73f5d04e8a322d7d5dcc365c0fe219bedb9ee863cea9d06791bbffd03f22dfc81489df7ec7ba0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3cd5535372424471e079f5290811346bd90fee218242b6df1c5cda2dce6ba36fe5c2f947d130bdd5ad80509203d17dffc61efb4424d5afdd98fbf3ec61809f09039d94ba6f06c18bf268827c6404d2ec056cf3547e0c1992055f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1858060b7dc6d313a35c2a5487e7bc87845024cbbcfdc7a35f8c5ff24658b2e9e56c1d69ed0b3c530d93cb1075751ec4e746b04e7760620cf78bc4feb71bc59fa127322d00f688240dd521a4e84842ddcb0135dbcedda2dac0583b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb472c20193276b8cbbf9beab5f2eb3337e720d4ef9a12550d604765cc46aae8a7f9e3c2dfcbcfd70256ac9427ba1bad049035402b395b20518bf747c840436ece11bcdd912b8696ba98736de09d8f35ce6ae6efef21c7cc723f0dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e7c090fdb72d582c5c663aba49336c1c39cf0f0f7ec8145ed4040b2e3a25482b6306fe557913e49ac8eeb7a6866e4fce574a6545faca3fd1b7b9cab703b800465f1cbd7cac90c25badf63d676bc57a56ee5340068fdf8b7c57eed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1480d15e9a569305249c3dff37316eef934d2d76182ad7fd8b28d87fcf11147891e04b8819de84ee9c5ba9483d692a2c43f7a6b9de157f86088c5eda474c1f231492c52cb538c7e63b25f08bece923903299306d1c944cd3fbe9961;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4ca9d2f3a8e53564df294986ce9a21e7e4d0e7006ea2b477daacc25a955530f0b63add20c84153d5509d1ea10764ae87d265d7bf2b8f543d6d65f55206ab592ac09a99667e8be69ebb3fcf47610695360c2707bd97c8df5b0b1b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd9aaaf7f4c19d8672db9badb59c9b499d0d786ab7d0cc0885a20de24a47ea210d54c04740a2db8814471bbe30c12fbb295b8e1dac064b9e312a4bedd6fe5654f3ef493a615ec09bf430a9ca8fb7c5be8a2e0c1b3332b76a473b8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5014b338158bb3f9a19acd977bafff51eee33170e98cc2d66b0cf4aa824b70e053abc23090e99700de6633a97092b1816a68519568d1551ff14c3b283ce544d6c7b452d08b1c968880eb9d891e479f1f23f0ae11aaa0803d1f7c63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1481ec98341a93ea46ca282513dc63d641d47eabbcfe8fe43b92c398b50ca336079a4725fe0bf6e67d8573ebfb31c092701e467cf004005a1d4a6e56e69f089e651e583f9e430b17c0847765698bb1ae8c72beefdff7a23c6543815;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1617b4bde657b425349496d24c2e4a7370f43dd6c53c4480b70a32dd94e0dfffb95805f839dc29ae6ad974a99cb38561f11589856b9479e2dc6e82d04c9271764252c1074159d25e9f89ba6b509b52a954be486da4faf6e1cd07f5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7176415a9a41791a0e68dffc98081042b4b467d3d224f68d5ff1030871ebc914b81bd0866c4671a498597dbf21641516a133b80e2a4fa057e2c636b4ef57fa25627b9e88628f31684536aa8396abbdca809e21f813857129d196d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184681538f25b4f15377c2e757d528d90dd7866abfc311152765df4feea5de32f71666525218115ca58534ca2eabedf6083519044916b7f3006b680ca0fd994b61fe8c8b95f57c038b950b9ddc136530463ca3a16657c90e558829f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h584094612417a202aa71c743ce1fc8dd89d64e0354ac5680fab64a67ddae3ebb142d19413b55b11c73887e9ed8e3188d5398c8b928c5a011e57a41bb8a802d9717ae0c7a1f51fb5a676f23cdd4634639351c687890ec4ed898a10c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he004589d1ada01d058ff201ad39c4024b756ad5904b4ebf3b6ac83f55749ec34c622bdde24923ae90efdd5491577ebd0ec1988e8e49a3371c972c2e5afa9d5b8a97cd4b2d7f1bc465298cc11940eaaa7eff515ac1c49831436c603;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19dba846413e2e20a7c227a47d1455c9e8fb40bcecc34ceb541380d7a04965fdea8b515698552e4667c23720cf33376248cdabdc4568a4eb72a77dab21bed96051b4eb1acbb64cdd8d224659c9f9f369654128717551bd744029b7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffc265ad5a3f01f13db45ecc12a5322c2ae55af194a41ebd73f501b1047001541a524f553cfa8ed7b76117f99c3173be27075a204dffc06b772ed0225f9ab382ffa73acf65cd50aa435e75f3241640ce5e2ab2456f2fc3837acbdc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1030705429fb62c2512c3fbe224096484fe1f3bf054bd9e7f21f0c67fc2b9e28dfba3af9a74d66b777b4018deeecf572e0fa0d86ab86190015c7be1d7607d8d1af15e518726b1f9ed8a9f3374706e39e7bf9d0a3acae1cc8e87f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1104f1d450f2befa3f8ac55da0d6d950c5ff991fe0785fc6f21d1de82578e7b476b5dc25fe462ca812f9c64d6ebfec8496761b8c15795dd3eef6df3e5956dc8575dfd57f201d743a90837ebd69abc4282e2a1d80dd279fbfce8823a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5946a1772a9a51b7def5451faaf5dab31e11dc84e994b8c8b1a66775538e801878a8cf23a0f46d154c5811201ebfcb3cac40f66c6fb13ab1260caec3003fef090b2df339e38bc463bde5feb3a71ec107466356c36e155038b1d4b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d0475765f00da363aeb6242fb6ec3ca49a2f0e05a66857ac76fc664bf8d1cfd6054145841b8a9e1442bfaaf429d130611ca6ca3b49e416f30c08635ad3cdce99d96ae396c8f71a055c8fe724e6cd2cfe4c3b960e00bdc6ad6aa01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ba3a97ae5839b176e6fe65d4f2dc743e8d6a83affec117db2677ad344acc74e3e686c7aac8155bc9f05012246d807845acaf72f43589b5ddfcede06fe7f83abb41aef808bc1fb87cdc4cab953a7806ba77eef5b4161e9556c6e66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b84234552111e65452533ccf5ee57105c59eae6b35f4745f7c95964e563e8a2677977d61cf7ff10db1527e930af4caac96b3bcc309a413ddccc0afaceb3b56c7940c13b8ee09e9f540e4f52a2d2350a9b87913d0a9594330ad04ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48d28cab0cced4db48ba75a6e808f588abadda77e3f4f5132c8637e51f8226044b3e35763477385c6f7529560b7ff9802f66d302be100e6d0a6e712369fbc19da9128db290fe7a3afc50bc53c4968b452bae632318c8b0120207de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1aa4ddac201bade3e3384361650e89e336341968c816d660a96fbefda9cf380830f87739bf2b92230d261e344b86f5e6ba0f8754d0ae66a1064ef2b071f514c35841321bb04f7c5a25bb538d27367d1f507cd341fd2867c2a0498;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1f9fcf684ed93bf139625ae8ff2e23e3aef8e9521a8fc95d20a2ce93401a598496a5ee0bccaaf0ff445d78086d43f1da35f63143563e7f422d5ed9f8f35a5d72c17a50f242d2dbb40608738aaf618fee414b6cfbb2b9d6d7aec24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5fa64be8ee51720c5244f192fa6b6ec2cb242d2d9f643672c1dcb8db4f01efaab78c6e727616f906a351663c38fd0042ba0719657fa332f937a8f5a20a3a68ceff1f36456f20a3a33dfbe2f51b04c99625c9f46e81d9e2ae25daea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125a0e74fb66d8f85f79bb563f8d8f773669b04fd2b278f1676729c8ea543491ee67631c551f8ca9aff66275ea9843fe623ed16bc28edf61b9c96021099b3486f438a15fc62cc1dcfff5688eaac66e877ca3935241ebfe158906986;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b4202ffa5e3115b6d443b0eedacc61b836c4ad73759f9eeacf3860aab9d56d13c5a0a8cc52016dd33d5e49a3381117c1dc88e22736c136e90b81f50ad8a7073dfda58fc4124792c167548e6014be23afd1fc6d552874c22a300ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h161109521639ec851085942a0270cfc6ff87d4300b667733b59f034cc6d69cfbd59589a927ea5f829c2f76c120eaee82ac6aaffbeadc5d088eae3321a35ea622cc20c29452eaeced9a421476f8549f41f592b485a26738552c629b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b3d9b973b47bae32a86b3db0c7a505274a91d5a9a7db4d6a7de7969faa771a9f179baddf91e6f6df202ea22c89990d0e7022970efe29575b2d7bac57807d92a6a28ba82e5449b6646d62c277e6438ea5aabbbf258d850ba15ab7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha072ff00ac6cecbacd5611fb7db1e55ad4419d49ec775fa7384074619433ea9edd1abf0a6e1e48b44e1c2980b346672c8eb68509116db053931e39ac238d0a09f30b82bf863787b17b6f3e216d16a9c67038047b32881eca945af2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11acad0c66826de3b99eecd27e658d5659fb78fd15f6e303cf777e15eb580cfeaba283c4b73e8c4fd30b2c68fcc9c7085afce724ab8662c4db08be91dab3a75168ea0cb72a077dd5fc263f90273fab5baca0b6900b8a4e6e28e9ea8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b337942718d855ed0b0d2de645fd221dde14da30a419cadce26025b3d2a3c1c539cf7aa2f5b9f2537a248dd07ebc02bb57da7abc86b4cd10892d65ed8b0573a4af9c0fc46a15891eb77d82bc5f0d97f171a2cb2d6dfad987822d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc6c4dec4cec47bdf80d6cb268a59174d4a4094334e127291d6d9a4facdf1de24221ef615019194193ed57ad4b74879d04af95ae11b8cf97b28156d3a23b78b1555ce6d9b966723af00799190a8617d9314106ca881c86c05005f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28637e87bb6e85cbc70edc65076d6554e690b64d57ca5a13026cbf50bd76992d5da758b5fe7b1909a6f1fcd8302ff262ed4de9bf47026bb03547e0e02e1ffa18f7e6fd975b32e4860ca50ed05df012d4dd64ec9d71ba15c9e33443;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa7d725b1fe172b157fffa9b5099517ba9a0cbb896e548b8b38b9d71bdaafc3c39ee963fc4b34ea9005cb80b6a5f5cbf2d905edaa7673e7c827872707fd9111ad6d70bcbc25196a28a6ccb09d1f9bf7b988e2cf5d400cd916589e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haea6dacc25814423d52cf97f3005958bca29939854a247df12b2fa78562a1e4c6139b4eed5ebc6172024c77163b14344796936b51ad3ae696cd9a6abdd624cf8d150462871dbc9b0bdaa1be23151e5d66d3c693faeaa83131198b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb13fe5945e81f9ded0805a213a1b5d1fd32b4c76cdcf5a66db43c008b56e2a76cbe6aa490007437df7de670fa602a82a31f761a7909fef89b313e07b43a68cd441b4f58a8825071e65cf5e968cfa02bb4b2ceeb053c687d4b57e52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e6557107c69c2102f880d441b8c4a6203a6f4db386ccdd003c1067212a2bf21467a377744e8320bd651d1f941123343b6ad647b0863d0f07062fb0962f903af791ccb36db9985fc549f8ea03dcc3e4aa560385fbdbe147f36598;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26b493e56d8b9fc1fd759bebdaec7158d0dd23db15ac45c4bc98af2cca466ebfd86e2fc9efcd616f98ccca6f46da32de1015fdfd7968a042e15d503ccd512a7dd48137ae23e1df761135132407f06dd0a28c1b62cc55582ceb2db3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2f8c2034de079e220e12226f86717a2b355d171acd952e8498e0bdbb2789654201cd81a72b658c811c824cf148247e9270d2c72f0b5a735a269c0f4d91f50c0cf9a68fb672e94fc230064774f6b1b57f1b5652418306c3b5bea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ccb7520bf4c74acd527476fbea8b2918ba1baa627feeb8b71f504d86825827b7c7007e27aebb2da4febc65e2011f4eb7aa70cdcabb7c176d2c54908c6ddcc431e22cc28ef042b9c5a33edcf6c2443f705f3a9d240b3a42c9ae8ef6;
        #1
        $finish();
    end
endmodule
