module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [25:0] src27;
    reg [24:0] src28;
    reg [23:0] src29;
    reg [22:0] src30;
    reg [21:0] src31;
    reg [20:0] src32;
    reg [19:0] src33;
    reg [18:0] src34;
    reg [17:0] src35;
    reg [16:0] src36;
    reg [15:0] src37;
    reg [14:0] src38;
    reg [13:0] src39;
    reg [12:0] src40;
    reg [11:0] src41;
    reg [10:0] src42;
    reg [9:0] src43;
    reg [8:0] src44;
    reg [7:0] src45;
    reg [6:0] src46;
    reg [5:0] src47;
    reg [4:0] src48;
    reg [3:0] src49;
    reg [2:0] src50;
    reg [1:0] src51;
    reg [0:0] src52;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [53:0] srcsum;
    wire [53:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3])<<49) + ((src50[0] + src50[1] + src50[2])<<50) + ((src51[0] + src51[1])<<51) + ((src52[0])<<52);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c8e4f0bb9425c6bb319c4b43241be68f6f94e9fcfd2e4e52f860459f160f906369c3919415dc0eac4fdcb4735e12cfeb37f105ee3ac60126d750571e0971660a5b357f656e589338137d8df8d610251566532a18dfaa47e63a7d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd8d7bda953d62fdacd4bf5ac99a8403c08fbff917e5926aab2a70c259f896747c55b74d7d63892afab32fb6bb5fc7cdf63fd616d53861e1cf50dc4d7d6978d9b5ec6eb7434926a5b0e03c7d50d4d33242dcfcd4db96a19dc7ae5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb68aa2756065d291c8954444a1b649e1577fce09a2560a2954fc484933271d4f3e821f43e50893733d0d61eeead6fca543fcf7b171e194ebb51249202d5ecefa5b3594b336eaaf16654c97439926739a53e1b226dcbcb5f8d3e80b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f49edbbd6f73ab79cbfe6f87d2fafe9e2729b5dcbe79989f49a1207c5d28f4e559ea8c4ce1390b8c3891b59e937ba4561332a4e96b288809618e8b84f01f24db636933c36bf02b46345f38ccf420cd5b22951aae222c33368962;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b046e26e921538da20be41f11067da3c2fed562ea655c9d21801ca0ca229576dcce44d07afccb6b3d7ef57d46d9afe83d85f6161dd11e587bc05b9ec2b2e5ceab6f8c1fbd18740df5231d79c8a97d10f4ad2c3b318d223eff99191;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163f31c120d39fe3c0f9f0fb8d3bfc68c7945d4ec286a54d7f1c01fd76f794fce587d1394ac4ae5bacc263559c61cbf6c65e0162467de421cce235b100e1fd4ea364f1408677169dcb00ccd139caccc98710abdad0deccfa35a7dad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111d871af30c375d2fa9aaadd404bda83dae6a1b1697fb4725543d6e8057002571c99451d0acca4c0cb6bd20d36f847a631a24e4952e189466e8b3e9fce67abd01a7413ca4b8c51c533752d52addd4b4c1c226b745e7fcaab7d2e33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h605ee7e1e7ed4e5ddb671a32222c5d406149995689d1911417b30bbd662de5c5069b82d7e539d2303ee02f28ab14e0733baf36c1e61ded2ba6eb760e12c9b96d197328376b7eea4161e860d4e362bb1a4b2ed48bc001108f68eeb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e657405935f158ba5f46d07ff61ee59177704ced7a0d13e48d967447f48cc00e1ffef346107b0777cf5219130e83df788c4e9e06006d32bfd39e14193280270594b28d6e4e63c4c1127331c544319ec406643920a063ce45c11c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e8acff5199afdda6b3adfe0f43662f108b52f4032b0d2d64b761834431168ba4711b794e657a1e9aca0b0d11ea832e59a0073f812894f4b684198af98c0754ec8565399ed0fee44b289958ddbbddeb1a4696ddee1ecdcc4c9c5b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ef7b5c9b48d66715c3742cd69f4346d27c5563875e6587577ca1f44db15b07ac9a6e420011fb7115216b9eb8d3b66fdf2f073ffcee4b2ebae6b5faede9d596b634872c09b476781976f89f6f7391e24e4acb9adcf3dc3b0f4eb05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144b675d1a2a5c8fbc6e228b22333137c0691936addaebafa900cd6bf8b2476311fb01592355f7ed070cdbdd1458b3e797eed459cebd0736913ac7f287c9a5f22726dfff866900f35c2796afe3199cd03a4bc2f293ed179cd21ea4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95fe66faccc923930380e8d4f327557095c7408d4bcaca5cd2d86727abe0f5a0e210fa2ef00bd163bcf7284a91d832d9deb55ccb8101b4251473289c60d25577aa4dcc84deb8e598c20e77b06a10552f7fbc197e582bad64e266d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9242d92c4ecb178588d4df5549b83b08160683118afb5a90dea58b42f09e1bbaa6d5e4bcd9fb90e14650d48a93a3fda4cc2166f17a84c096a8c0e69cc7ace168e706e2f5896a8948304d08988edaab9e5e87f7dd06b7c59b9e5981;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b03b3549786146db31f64b53d1a25b61360f0e7b747dab67e8d2b0d4d8b0fbc8c8f8d6e460bef54b79034a66cca0fef9f816391a8ee1d250837e4a5baead1de7601fb641924cf6e8f17a104284d057d23f676c51424ed0ea08ce14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fde60be130017f7e1693ae4a8783965171446368375d5128356441ece75fcbcd68eb6509b831f42eb02a2708525e462057192ebd5edd319140a564cfa624449a3ec1106774814508dd457cbb380eff998de342d1667bf73a55d3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec57c59b6b848825813313c2d11f299190e5c4f2a96dc7e51f8f1853c95a7fbe0860194a7c03bf009d70af394a8521944c58bc287785a2faa4fc712e0a681db7b8d063fde9f29a90c5122f00baa07aba2ade516cc6bbc2951dee28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68bc13bea235c958464a0874cf966c58ffa35fa438044f6d44ed3f31b6f78bd46e1bf572e933146c5dd762e4226638e04b98522680a862c4384d4d949e14426e7abd79252aa2027cbd14a2b53eb86c6bd29ae0265b6215ac95c33c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26f75912b28102889cb1c1a2c0a3ff7e26329e8d0dab35dc25b588b2a28c5137794f1f147d75a9953dbce59031ba4dd1fe011db0128b9d52d9a6de5060b7e2a50fea0bc70a75e7028e704d94721cca2b11ac21f346c3cfca63b8aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6863cb8aca577e31a44e435e0821d63d1605d875a939a30e558b98ff41cdd801cfe80dfb4a9ffc3290f9c3ab5ee9102c93e386a0a5efe7f6e87589b40fadbaadac5a576479b1a524fcefb58d4a3a3cc49398e8931c32aff7cbacb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d5302b6a29287414277a4743ae9ce8bd5cd1e50108e5f11169f6a30991cd0a5bf5e7e90817644abd946c734e7648feb34993b3e9083c7f0343d2018a1eaeccff761cfff9f5d71a6636ff43c967a319928ec17cec0de070bdf8f17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa888b7d6eca87f9ead74a4ad4ba8eefa1a9ea066e56610b2ad13ad0a9c3bb3132bd5465ad4e50ef638a9de9d3105c101bd843c6493757bfa24f97ae036661dcf61d37c310a1cb261cff86fc4618f1269347845fb2cc1592533c63;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14784533cd4d94277469786a416ac9a66a4cc8db4c8587d9494754e3e19fa69bdd49a76d8b980e5b1ea1cd966954731191ae18fec921d90e37ad0fff00348a466a4494d9b6df7cc1d2ade5a2c44b77e11e7c17cb0e498ee31beffca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e219de0321649ed0fdc921727979b5378f1ea078ede021fe3413601bcbedd7cc56802320a9980eb71d6f269ce0c5db15122d5d29f69065ae47750ac9b0b05c16aaad0796ad9016422f7c3fd81772b7096607bd938db2758ca8e3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he556f8d9a0c59b270ae7eb734666ea4586c3c6ffccc3266277ad69fc112c0cfcd876c4eb3609a2cf6f017c90a30e2aba91762c8722e1cb0fb6195e893729a21562e43c4a98e287dbe207420457969024035d268ee6ea368cefa906;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9312ab120e8ff6a434c869d6d4ae54de60ccab1c71a107578de9546af0dbc4877a8fe0a9b158d86ea8910dc2e399c728f3aa79680182e06b3714586ca5ec49207a262223f1ca8eeca1f3853be2689538169c5252f5038b177d4b4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17849c48ccd2aa0b3395e51e04ee68f579cede55fd1b057a0248cd4a38479306a7e78679f489587a44f3aa1fdc722efddc043edf501e8a494469594c5af1e1b2fd5b6fbba6f10a04a13c21c597b885f029b22d380f1dedbfa2c06a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3f9b23a0dab967303a8026fa67ae5820329f7ff8952609130ff703aea71fd9fd7591c7e5ee4b2bd79bcb75fe3334be530d2aa335b58a046a3749a00c288af9324f0aec1d23b7e56f4e08faa1abe2ecbea178fd5a9f445cd8fa6b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e61a08a9265b175eaa6c39e0e4382217513a6ba6c1ba4fb95327cd71c215e43518bbb515defc0e10a982ed3bfa25194060a79e26c8308a25ea58cd2bef55f61601eec0b9844e78585c7298c076c29b0766105b7146436729b998a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d657a245a10a6918b8518ae7424cf1eed72e5616d84461d6c211a67bd96e1bf17faeb3462fbb7534e1c49d8d39de623fc31ad715899d43649ee5c6883867367c27096e5a143246f65a7118cc52306e8a8f798f93f059579fa5fc65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f56036a0f6ca0dac1886113c2c3aefebd56fbfe64298934d384d4e62705ecdfb50c4038defe90450642b26bb2d63b17c013d182dfe91151f0378ad8b980eb6c793a5aac2ddece2bdcca3da3b2178e95a6cf2ed682bb5f3e799be83;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45347520255a0387bda43cee57230925761ebfcefdb0a2b7442c6275c5d81222a564bb8c11881cb33a29637eb52d70fa0d7db4bdee6da7b782037923fe989340a469c77b139aa4913ca1a715b6796cd8b8b279ab9f72ef6132a080;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4f1a537d0b16efe0709b92c4bc7797498e5f1ae7c680eece67ac41c4422cb7b29a65778f08050f54d7026ebaa2f1c526663f98ec62f53b72145d7ca2845be6dfd90fc3fb08507df5c32d1437e4f0751db36e1f1c925959cb257c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a8f034851488994a2fd1f6646cae2a1c2e50f4ce3cff6945876185575b892f683822116974e064c529dc331ff8ee04ed5943671d1c39b15d1b515ca2ab92840309ca9a940a953c8bd1d632e9aa3918446a34ae637f393dd6c5744;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f14ea73523417e90717cc5515145e2274f383255a25555e2eac5a867a80e19e85ab3cf834ca8ac64b528a1f888e2f2aabbf52a5f4343639eee39c0514a00f005dcc1b24d567c9336b26d0a0e86a49cd8081ba4f1038b9e234a54d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d4794930532eb3cfada5387b6d56203673532d70d132e4749b94190850f6320fca1f36ae5c28f6dac49689f6bf2c95341bf54657172dffaf9d84cb8c2e04d0af8958f7f76d1c075768417301d9bd44b32056a35c035483a2f9175;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a2c0d53faf67ca91d5efeeae23cb74da839025902b056efb002c94af0d98833a4e6ad339a0b16c5726382d4081e1f8952f6b71dc389b7336cf04d44a4d24406bfdb5b1f8f676cb155295205de3735bd2a6db18177720a9605dda7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14704032006901e2fd5cf5c52e331b5bb9bfd365dadf6c6fc1578e6c5d40130e710aa7ec28d8ca5f3af579bdb798da56e4a8fab23f56e221f6e8f793884848c1d3003c7a53a6766ce79d7f2c438bb8889c4ba1b1648635eae8151b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6e44f4afb23dc4e94eb349646ce97f100e2fe674acb0311a5cc6f3d818f9ac434186e8650354af41a6fb8ff8e26814fd95476f9f7bc8bc2ad6433ee0136ce93071c96560cb11875280270106215c59f14e6e76edb054a72c97d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bf3712a3a4152304920eb4c929dd6607edb6d70e5ccc2566e389e246d8ed23df38e675c52c5a7d5ff17c4ab61399f52e84daced85652d324974fac099e3c46a6edbf3571f7ba9974f988862ba6efb67e05755ca3f084a7cd50fcb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6086d877b7f87c073174e13007dc94214ab27675874335c033e64e9f99d6f9de99e432029f6ca81bf82081abe795bdd9e17f02e64137100570301d3bf2ac692da0a4cf5b646fdb52174b29dce3f5c0d81214fcd7bd9933f70db366;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c814044d8585a2f51fa5f2faa8b54485a390b821f21495382b77b568ba9afbc1c453467845f64a0be7a5ff8d1a1f0281472cb7ac4b706f49fc3b9752ba3a3363740703a1cc914a3e12626afc588d20d429c6008d48321ec59780d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc144dcb0fad699b1b3201dd68d8e462ccbfb7ae100597b7edf1e760a1a1a73d49ba0c81dbee62e94984ccbaf428092aa6b7fabf6dcecbd19388277b924048bccea49cfa42fca02e0ff48fb8f55237beb31ce0cbecbcecd4f5200af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb39eeb91205734d0488a1b3a06a9b5620b2476e0249648ea4d228390bd797f96d30e24827390ffea839d749988089d81094c7b799c088911b5a3050caaabed22268fd8ca9035cc8d456a4e8637b049e8b2a82b4ca8ad68a096030a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30fd92fdafe3020ff2449ac9a233bf16056d0b9f50fbace55392e70e295fd688c2f63683ee84d95b6f2b2e296316fb29e8ad13a05eb857c54047de548f379c583556c4ef112c96464ddd4e58d2ca58e3e331d19ec6a9565947baa9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80c85fba720f8cc53839c78069f0e64ea85c302520c242c7a408e06acedeedb0696b94890c3ef0f9b1202047212bc270f2952321aa9ece8b5593aaa8ac7b56a357ae3487d8807c1ea3733d7744344fa9fd20958a81dc9b4fa25076;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1132dd652615704a18b9eab95af3507f88c1970977b248c46293169d58267bb98e4d5ff4603a51df4a92f66d767021d88ddfd41acf863dda6b2f152a18b63b97118c048200ab13733b99fa45c2aceb833bdf92b51370c9042432dfe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a79fb9b0207b5c1d419e42d7c917ed6d667aa0ba3551495531a0d61817be074b638f52da8991baf2782e1f6ab169f49ac4625e6962f0a2a2d7bef787ef7910abe88a23524798541bcc85c63d6ed06fa6616a82366c5a6eccd4f51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14184a9adc3dc3a8faa478b1a09b11a2d418ca5663681bd9db9013068b1faf5b58485ed55d1914103e42f5a56ee60e9082c71ac9442b3356499e78a7fceb20dd9f6819ca482bb95a80de0fed5d491aa71a6b4b75b6a19fee2952396;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e502bd81879e0f21d3e82a12857abcb80982f71b8413944397cd1f172e638b7ffdacd3b502ba3194bdff15b110e45d5586fa326860969e932910cdbbd7fa05e92874521075873d89117434afa23ce739bdf8d2b4e858205c2207f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf37f59925b9a88c68dec61f1f7f4d630d09c75999b143078f168cd46c44361d0de94adc1302dd334d3d408da3dea6f32ef688ddd650070af9701492d50c0c942790c1fc282e3b735b98b3129b88f06033d3f1f180eec223dc6280;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h898ec6f24f6a36cfaf0619c216ddac8e22c7ed22ff084cb24f5421099dd1059f2734f842741ea74220cf92b2afd92ef387f8543ca261412c233366d7210eed9b7a94617108e09b5d58984a17f29c208f5ff2c8f52af8887ef02b27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc887eebbd869c39e08827507b42e373656d51956fc9be32ff9f0b901da00354ba8628929a37cde80734b8f81b8bfe5e13c2e292cb381a1d9afd8ba729466b9680938fad0db159d5cedd52507b7d97a2c3623b612ebeb0d205fce78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b4843a8a26aac3da70976fa27780e74399ef0837d4fa3c4790f72d4b4d7e251270b61bab2e9962ba20063a7f0674bb2961ae05fbcfaff51bbd2a6cd671ce9a450409fb76a879d9dbde0f70595d203c53bf07db1bab480da83142e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6828806f4e393a9936545c003d7ffa7236d7e31a507082004addb07f06bcaaf5120dd85e36961794dd2775d8b8ea4385c9f11597b20f634522aece2c0773193f3fc43f7c93d828e020d9ddc1cd748c47786c04ad5a5101d7ab9af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1334d2759e068830798cb4e08322a6c27b6daf1a3721997d3aedf28ec9aa977e0b3e756a020d43d18768c7e71b1b157ea8207288c81cbc434bcd75bdb63a0eae9a8e338784f616d6ca20fd39ccc1c3d79c5185c2b7c19a545930333;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccf141c4465a913c90bcaf2058772e5ed3fdfa496309e712dd584b402935447b045570d39242b0760234fbb856129f5b28ebeff3b1c64f744a12723074a03bb2d057e0c97f58b20e35cd7f8044adf023aaa231cdfa494bcd303cef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb2e3b233742f07725c0a42b1cd8738ebf55dea47c6aa22a698858453698c20208c97617e1b5b5e447ac0395f0a04432297eecfce09dff65aa5e05dc7687b6f234387ad4804b39a3314f6fc0ee6fed57dfa0417bc7f2d112ddb61d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc2832e3bf250356620300ee543cc3331037355d0d10526ce1f6a51c2908569eb0e29f3cbcbca4f5c3c935337bcba65a74c55492bfcf8ba50cb8b10d8025436f572e5237e5472e918736c1372ffceeee708b31ce81fbaa66c21753;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af7b7a7f90a57b7a116c2baf8b72fb6d44c6880af0ab53ffc92b2027eb349b991d6e24e3b868b980d2a0ed0950e63660e18e41ee0a3e82794fdf5ca50e21ae36f389ac7c7b85f5d9095c2bbe7712842b1476c4676dbb1fe2d12c8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2234c6b229884261ea9f0f8469130f58057ff4eae61273f38e052d9a7add1c2f0a3fb680e553b2be1d2f5e45f0eaf587d0ff97be1f6b88be301f041eeb0a7e9c795fcff811841e0882908585082cca62beecd33e724d511255ec8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9aabe1965fad7d461e6e7dafd636eed166ca402476514f42e2edae536b292ab50942a55bb246eea49a256112300f4c9461f21c8c1739445e6d9d1d0445d721b343b7c3da48a4b3026f0821f6f215cecf691edface45c8386d9de76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c7c6e05e140a59790c67c2394b37e3c6ca0daea7a01cf797a1dcd51c3e1fd902a8910f04911848da8d8d45a4b6618ae19f3cd8f530b99959b56516c8cfc803ff0eed0c75617f9bdc4612f79981e580526ff0c02a9b170d4e7f1a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e93176b393905a9e4bc8218da7d7a1132f4aaae76c26335550f284d91a0af4c2e55f30f2858d216caadc7b9fbbefa0c376d8fb2103d49d6925ed3ae27a3345100132cc66f2736132dc0e6e1e7605568bc6e57da7203701122cd55;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca0db672bd214e5e7d211e098b6c73713aee3f710bb4967b9fe8df3fb6e426920d20a71b1b60c3ac1e88d2d118934891026d04406f874af50113e88206d1c2df65a918659c0f13d38205f607ded48e03e05191eb93b27460a451bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185c4ead7711fcf1b7a267e061d0b1c00a5fe0c276f6b50d8e4a09264dab212ffecb914130256f16d1a8be087ead473f31191d020bf76a46217ad5ef7ca93c905776b4095606f75f377af1f003476a6a40afa5dbd798c1e8f7c8430;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2390101f082cef6d7d1fafa7f7f4a2b8c20c1fd8df96950cc23407f3e70a5210b3679b8f4b83fdc627b5fa4231284b10b26838d4e7cf1b2b0ebfd420f74bd0bc06aa24d917df80ed67b809ce18f3b7ffc25b413e00a9add515008;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ff633ae634892ffdf86c8edacd9de7177acae62bade1f2446e0405177846a19632b4823806cd7ddf5a0711aed518b17309340533b1ae5631f554a98ed02df162063c09295e669f6fe2fb2f6a2cd6601cc1df2faef5f5b7b49102b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a594b17583cf634d520bf8c084dda818222860f7a7eb0226315dacc54aa34930032abc90160998cbf9275c7fd4bad20c11dfd3addb3f8c70ad449bc817415ec968804bab76043436d1a0660c6c23653559cd464d36313b98e296e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c179745f139975325caf81b7fc594b1f6daf9add67a65fb77648c88aa1ad2deeffd2b1b37b9bd4688cdbfde6899e59e8eb39f02ed22e04c1f538ac9813810b72048432f850be114cbccdae59163b6aac90af24c8945dcf8c6581ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146465aebe6de02d771b7469d4d5e3ebdaa4df5a35401801f4ab37ad37244ccf99e28724e35bacd37088a8cb5548eb3aa6f650d4c0441ee2c602aee216eda32fb48ba92af02133d1d16405acf810be907cec3bcebb0237464ad9d2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e5f2fe8f49799877528845b1c3f780e440371f3244923eea2301b927b942f11c9b971420ef413a7c25d6925df979aba51e1f8925d52ae8d9de73193250d9c42acc3662ca5d28d8cf95a14b47569be1f7ccc676aa0c86e0acc5e70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb87ffb79121a42eb4585f341c5241f9ea911ecc62571a03c08d98ae2f4c842b71dbcfb71a56a29ad931f1549e5c36ff1f0fefd374a92aef00e8ac1fb291cd00c7b8c3a65333efe557a989d12fe293abccb51afea108c0e62fcb0d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a64e61ef77f15528548386b0f23e3c9fd7f890163144cb774dfbb514f5b186dd537efe10d781a2e0ce5bb29f5cc17fdb72fc97fbaccb4681888e23b263f8f3f68448b39158d6cba29d83b9e0784fcc4086542f7c55e4321a299f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9bb7bf22688b8b8772c76505d18512b43e5363901f9356219221f1acd18fb1c456a98caabfd51104751a15f22134595c7aa46e6ae30981acdbfb2a237f0b70a3552dd2e3f5c083824e7ccafb9e6a9815c71a4b7e5d90545610030;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a6366619767c9030a548ae556a1989e8ed25a7f5f145351773421be329c180c4ec3e115d93d665454fdbb8a95c6da107c2c474e51139b446538be0ccfde7fa7654e58bbc844954f559f08384981efbd9cff0a7a3661edf49c1d03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78610433356dcd16232b59b6a5380ac9086900d794f54abb086f7cf778930d08de3eebb3a7746f2db080756c5bff440461de92e36f0c2f94193fb48a33824a65ab6a3068cb09be26c5ede23f138f47c891c729c06a73e86da7fa49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h644f2d68f5ef17846f47adbfa50e68fa5a00e847f3e1acbf325ef2e04db311ea0eb0b1724a249d9f3c02c319acdb7a90e0780231423a955f484f4c742f86afcf3c46ed34afa4c63af60cd35917bf0268a8ea9be173af62df118eae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad1b1a85e814893dbb88512aa009a1502393f844f93e55a22b857f02fc767adc6630d44f705d3c6d13cac47ba152f146dc0616cd30fc835a397febf25acb5b054ff144e7fcf757aa9b2c6937893e537724f48f74d1b107b0316bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecc8c2ba30cc5a50273240206d656a217dccca2553fa3fec296f2def7d43cc48f3fed80e6e89943d73a0aa063fd752f594b72042b0ce2d4f6eeb182a585be296014a9374750ac231b9975cd948f86d7af050c98c76ba0666c01cbc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdb9fa19767155ecd3d363b14170880c5aed62594b56596227ae57686f87fc9fa88764f786204a397707d5ceef75ed20cac64631884cce9a5ea5facb9bfb5d6dd1714fe072996dec51c374ad6b34e26475454ae9f5cf4bca9fd902;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab2d3a6107400c9207e70f0ca206f07bf301e6a0672e59935dea0ab7de2e15c80df46bcaf1e2af1b2bdf6b50adceba32bfeafd2799c2af41f80d05bd3db1315cdca8b03c2e6496bdec5c471b6fcd617d7aaf7f26269e79b09f1194;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1507040b3ad8cd4dda30c35fd9b07d32297d519b25b15139a75d54793bd57d138dbe7e3d1e42f560ffa9e88135f72d86da1a3203a0cfe09b015b532c66516f588f055132e81faf1a8c0c63dc03b5b34b26c2b139b8c20b0fc3f94be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a1e1ffb13a86f52622dc56ab0e71a992e2133d7a737636fb54cff6422fba3fa83c369f2083e19773b25327ced77cfb7ccead4d389a773854ccdd36e456316206308822481a168f83340e37b152dc6f2271d75d99f88535d8fa075;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a15c93bff16cc1066471b954dfeabf76791cd3fdc51367b45d6a3e571c029041784587686c9e265a046ff74ac8e4e70285d27fa721ef6eee7b4c97d85cfacbba2b83f4591fcdd6680cdf0f5b083c03ef39b742db8263a0ea1e58b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd2deee672673aa5a1b96bec7fb2437ad3c61cfe3eeb39d5dfed4c4b1656e36e988479d40ee490f7e007347eae23666e1ded967017f97f359df10c4373e913209deaf21795047707970089331ad563377f7eb5d385034767dea48;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da242a7f7ecb3d8acc39a1aabe3b936bec2368ef2171d7bf3b8aa222efe761829326f494fb0bc7e05edd789227586ae62d2b5ec80dcf63c064f613533e6d69963f40dcf75f8ba2879c88c3252d40bd5bf27d7a88208c0840df6079;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e3bbb06a36b3439ed4e550450f640ad71384bb354fb7587d7c0c670f4d0a22c4f12857de69fe59e4a9fd7a9f356225d631d91c2cf68e28a55fae2f9b6098db749247bd643a2cf9c2af22fc1ddd1213198a091b2e4973591b6ed8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194ca64668e025d3d2db28d0deefe9632a83f324a0a467cbb78acafcccdbd4ce2699ee1b8de751abfa5ed2edc90f6c774f356307d31c4418c66c3ce11dc3e9fb75529dd37ddf803baad97e747f08b5b011a65bde31cd4b6a2145abe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ce8edc9261c290155da0672159c0c82d5d23f07170242391f07347249824687bad7820f91d1373a1998151845b8fd269428e0b51da1a868fa8b4d4cbff120d2c1aa08851c39b118407f7f69984eb65f283805b4c308dc18b531ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d0b06ae45fca7dc6ca290037d6b97577b02f5305b7334c63e581f2bf1baf1ac0e21fffd8ec6b3d4e1095f027a705eba366f95485bf9f27a9b92d6660f92dbfa73ab73f85ce4d7f70bc8da23990e3da726d525d4ddade9472f5daa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6dfc73e8ba3324a848f9c2b4840dd958ee90c574026b8579aec741800a4a611565ced761e354aafbc547fa9b023c9e9698d06497fd0e23d3235f15016faad651587c80a3732989c4e2462ffa199b4b5ff304f8796ac49507019a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155bb4969367bf26a71aec21d034c1136ba66694be609bc38f0893cdae10b33edcddad9723bcb8cf46b85eccb067dcc6ef6053c547be5179ddbd2b60159aa1de95ee291266e7fe53b13a66f9aadea45cc41237592acea86a408f6dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5ad42f51f4437313f59f4926b20ae7a2e55c4fd9d7787b3bfc2d5df6a22f4febbe7bb6b159e4f4b3e0395811bb49db49019972353ec1ae0519b75da223a0e1d0122a14618957bd02768567186980677a6dcb1a726d47c1563768e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d051b064bcbbb25a1677e89e8b4bef72ee1d9c9e0f10d912b7801fdbef5411015d9ab07e4ed02de945cf4bccacbcbaebb425bd7824cd84c9a7fd071f9ae6b22d405b97afce23b384235b10cfcfbd6b1fb1f50bc9ab52ebc06bf8c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15203e843061e57f9500b3dec1c78c03aec16e68e57b9a52da7243df241e63e75e86c8cba2d3c19b2c8755d1e95f418c226ae677b0b6fda2dd270ffc11f770eb9ce093717c806f35eb4dabff1370129d3e71606008cd34403c72516;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f4ce406e3fb83a9331d6d78dbe2e02c09851a0ff4d0b76d2e1d56e170f6eb9e2f9c3b6f4d744272f3ced34dc0f5ca81bcdc8ce3db39d8cdcb3afe6cb7f7cb371ddfe8aa886eef5ffb703d210ab7baaa4e195860220f316167de07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4dc44cf83af58d4f30de20f7fb73f9d79f579a428f751a7f8093c86597795ee5193966f01f7ef0a790e67058d1a4cb648fe63c1d89f17cd3b7207efc8829954076d6d8c53abed2bbcb203393be535aa2d2fb0be63e25fa1217546;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e97c3e58dc1dc42f549deb1579ae49b2adc891dc3e956bf22008d42d1e3e309b7f7ef2d4eb7bc35de0928dbf1d8e185786beccba7f9bce582d2eff78fcb2d4297066e75a1f757b356362380c43ca70bc1403230a8c973612683880;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1868ed9155c900a64b6ea854d6c3fe41b8456d89d9a2d17593fe44f354b38288162956f6e4accdc593f417c997c42a1762b35b16092a11835271a255cace007bd00828e80b7da8f2f6a85ba6de30586147098f91029b9b922a14daa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a8a5a0178e215bc4626755d0d36c746edbd83487608184263f93545defde4c984811c178acf818ad11a5fcdc86ff088a458e6b3060eef32cd34be952e6bbe83a9068bdb25541a215360b613fa260692499960ed93148130de6c17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1050783799bc53f5357154150b255eea8608cc56ca7028bda89ec781bbd4c643d247308d6e3846bd926092a2b235dc8c528ccc48ca7717df5366167bd53835bff1e5dcbd3ceb68b8dc72aef6df83aa0790bbdf789db4f58ab09aa60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1888856e2466117f72b39ca19c2063d62a0558b2390c60be13df3d07f4313097284efdfdf6d6703ce7d5356b557a76be95c74c9fd1f732341e1dd13e60f9d2eb22c6cec471c13f944df6533de033fba2509e32b91983b2d063f8e98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1261a4140f5d37cbca978f09a0e46917655ee2659d761f58c185596ee4f76b1d82d7bee7bd05d30291515f344e0c859c9f66affddefe671172e3fd8d3d004b3e4e044e148daa7a2aece12676de5daae50ac4ce9ce776e05b3215f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12078029099b81eb9f4c7519271ec7a1b7f1976b8cd591e68470c2ad4c0c0803180e6dd31400b5cc3cb80b8d69ad0dfe9c416e4b895cbdc78fd65b9a80e3c9feb68a3306b7789d02a90581065a0a7db639328ea15497e4cd102df73;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf21981bd23400616cc769c62c51ffcbb099a20c08eba1f641a50e6d6e00131dfd68e61e547c6ccddac8a234141f137fb268d4cbdf2e638b944abf8a2da9cec53622609bcf0e60d2f4bb3e4806b21e01f205e6277c8df0426c48e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e6408d3042d1ebb750370f88be321de7110f28cd58c465576d3a46f2ad266853571c5628a9bc424ba4ffc69e027195614d9e55d83de31296c17452a4d59ce3fcf377671c0c2784cf02781f72eb0b6d8a293f847874536ca039be5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff2ffd2097c68644062f7c64be40262f5c06475045cb805a1ccf10658514bda9d20764ca81aebcae646e12deb193a9ec8e0010716f1394bdd0f0de6c55156d717347d475239e9507621ca5236b2480ef85a3f6a795c07d4df8e2bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a24dd774ad3322c93d8e61b03f804d80c593c9c1ba4b1a5f0504250eff81a4c55b4cfd3eb7d1ce8db7c7e4b3be42dcb8105633753726d65e2e99f9916ccffdf0fe4521ce65f43675e932746723ae36baeaa00c43884fc56d489cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfde7e48bd7a87b00a6368c08fabdc9bd78c430506bd9863e219e30b4c949af765c0185b82a05613cc1ae8a9b6e7062c3929c69eaa6efa29f535b8eabb92833b0089e84387237490108e186015fd59a445b170b2f648e8117885377;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6b9b07121d40bcd4bebc689ae6f9e1672b4f814abd3643bd55426fe176386571265feffc288d647996f0672f79499447ba05413c5823523a35252a490dedb9fe7033380d471cc0c79595c4240e3e9063b7693d73a86263408e783;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4291472c7f8c6ea084c46f37cf3d878b648aa51d83ef2c2c16d5da937a63892023a695f7b056fc15b80044cfe95409ce3fe90377fa4e7f90aa9cf468254ef0fa8459416cc1bf75650a569a4dcf850e58df57a9b5d157977cb51d20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1524ba876c546e9492ad75a18a4822f8096003b78be39de5ba607959c610364353ffeca1ffca8d486d91785337d0b4f3787c33333fd3bdf95ad8b9af06e550641cd322b358e9e70cecb3d9e4f7a63ac981f27b5ac11bf85fb362b74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fa9daa9e98417378d408e2f70605e7919ec7bb80a3a62eb59a4bcfe879f18bbfa880dddea9bff56538ef2a2fbf626cf84c6a0424bb821314807678337b4252c1e0361272ef8004250276e11a0756852f503e64b4356e7868d87b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93ed4a444cb0c02bd0867daeb6ec66ace8584c16a2a4e3236307abca2300465d191044a8e9888c69510f9bdf17888829092bab96648ca2f060b4c261678a734e8735a06fabc6710bfb9f74a4f2e1563786b8c264fb900476e9092b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha554f2572561b590b3bc6454a2cfa91e7fba9a3c4445a9c299596ce7e814f21f3aa4ed74998f6a614193d54f9109a5cfc7cfeb2817aff3cc3f779121b0b5b946a4f926f6f33ad2a23e12043b715573e33ccb7d709196b7842b4b9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76cc563cade807c0596c2ee1aa6c42e13b4f177f4a0fb85693e351ddb51d5803d8a47f1fbd49344eebec0d4220f0fee43ae4386309f3a7beddea8e1ffb787f70068518448c4fea95cc7d72bd2bd8a5df194e8eb79e1227734e32d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1edfe709931690dafaf3ba7d47bbd025d6da5cb48ebd4d3294acc2b8a946e9309ac143cbda49e2cd12d9ee13422a6d7e3d75b4b6ed4c737daf3599cb5b3a02885f83048c9ce23e017bfb23a0fd0a1c5ffdcfdce71050e22a5673e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ea88d74260207702e58c235170b9daeecb0fe3906eca4021991207375cd4606d15f6cc60157c4a2bf9f119753de57f41cdfa3293c2c02914d3dcba89c3da21db4c1236d63f2125ffb56e7227b08f2da4337d450f0e4ac4bb85ef0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a8341b34cea84492ccf5f14113c5b58dadcb4d05fbe1fd6b77592772550ede948cb779d94b0f9d6c3f6e7cb764e17cd1d9b63153ae5a8191ebef228e04621c7b5146eff03dbd27df3d24fcde942bba0e1cc657a81c909f244fd66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1192ba036fc1904bd2a26720ebe1905fc928a04fc555a94229fb9e0dd1f9e5f58af2555a53dacf836fb98b4694f884a5864537afa532e9a4120b9b764564847fc24c6babb6c44614e34a2d30cb907769b49d8b4dbb1b45b16ddfbbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6141bf235962d1a6c7091b598419b4e828c1543fd4c4f04d780e3556779d54fbd85d55896c717288f56f41d4397f245588a67fee359dec2987bab5498b78df22def2d964d63d45f3703f5ea6661fcdc7da99db14d42425002e6ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h778e4de91a9d02791f3d6b9c4f90c239551eb494917a03e28bb2037abbea111c2cb2aed1a9fe8a0c006fd0573bdc4fa16f566863e976518572d1ede0d3aea87d527e517f7d444593920245b2d839b5f2e846a7ae089bace4b28ba5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee44af54acff9b5774d746192b6c85f0072a1633cbf8c1027aa01dd19891ac3ba1cdd550047727f7cf55349be000640a5c190c1eb4efe69809957ad0cfddbeaf78fde7b065adc7cebb1a01b5e64210165ef4a070d55deb84d8609;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ab193a4d179a315a0da76f006fc3af1ba9ac999efec73454a2317137358c31de062ede9c966c65e379b7ac6229d32d53ed2d693a2b5691c505e7230dd4f66225a937a134918b62e9b17a4bb2e1c3886e268bb960ea6695cdc26d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a16b23e55f7b89631e9ef84cc14850a177bbd0e5b6fff2ba762f918fc52fedb7e5cfcb2c5d57f53e1a420b76dcae2b405c0a71607d0f5d2ea35abc61153447bb577976c81831cfe528e05fb843763820a7a10875b8ecd3014b4d19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38ccdd233fe51d10b9904d7139458c556f8256d6d9d61a76ecbe0f8c1d45d919f8720eff18145b7a1be8151ef9f8984c4c2a6fe99b2339059298350788ff199bac75e48410081412a6f414acd3c064d9b08b33f3bb377a9c5d3e2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h409687fe4d0fb5fb848d7f6f001079ddf34a697dabb57cd03ec202ebfcf2489537edce39bb91bdbf1a9ce3655e57f40dba6fcf0b13792ef918661e321fbf93b8b72f36f4580e9b05b65cab934978afe6e95c7f1e2a74596f4e4720;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1523ef0f8865919b4f33454cdd55252bfe2a68c316052da548b61f2a774c5e731c75d38aebb0fe95f1f2bcc14f75d8c1950691052cc6cbf0777ae55cafb33c97c590ab119f98a7aa87f5b9bfdc1d668b8ba2ef52c2ddf584c803d1c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h630e9966e4504dc85815d6d33784b267f78d0f58569f8f6df4375e06df7f360c444d9bad98a443b96688cb06a91e0df1a4325bc57f634b52bc18db2f11e32361c8413f3193b115569096e5f3cbb3dea27c51b8b5c0edd9e603f55a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6080494fe0cbf25d30ae813a492811f0fc6bfe904a8562ad236369e04c6140bcb631e06c1ae9aacebf95ba35857417c3f77842a26f393311a1ce51141a41f5e94846028160ab6526d027a4b33422408ed7eca8359c7aa50e3329f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f0e434801367b6cbb6cad016990e03b1009b5bc37a4d48420baddb7b342602a704d404b34e28776d14de153e38e2d7e75e808885175ff44d26b7d096e960ea9be68664406e1e652193d671cb9e4ba0611e2142c8e503a58884a60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eca1bd796417f99057b66c98f9721805b2ed0d73ac6e662a305e5fd57362b60e5d650470c723bad26d60c50194507c2c855b9d1e3e0e2088b352b936fba61f787b89434c424953555397779fd8476874776c40e567cc515bf0148;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hded86fbba3e6239c352d81561189fccd10a89ff4c5b5f234e7052b843bc69f1f7a8d0e7a68593f947d24f0e7c7b121f94fbaf32a4588acb924cf0729cea0ec782a9603217d038273e448b32e66ad45b39ea918451d588dda8644f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1292a555f973e23a73b759c7651d4e0b715276b54e0cf70c7ed7d42c561f03695a05ce4a951c62ba327a1a6c91240d041d96631735d14151a27f421ceaf7cc67b6f853b9bc54dfebe958de1861002774556cdd155074992c09a7225;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b22dfb70d088295c8facfa2979592952428cd24c2b69a96d5f531fc3f75dcf75f63b9635fbdaa9f6158988b56bfb619a429f82559f00c5483fb298f524435384ccd1f16046b3ba237ea7663d083924bfe15ff2845e6ef96308c105;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fa6d8091d2b2a8f92fa5b733fc23981b669cf835573b6d25aa4e9497b241430b4104e40382abebe01be7bcb19d62601eb9da8bbd17c7014c50720453a9e3dd6a3e71c9d7d58ea58b6844c7f745ef462507dce4c49297e2f950898;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cdfdaad221942ede63a5f40f56a57a10b18b018052bb1671339ec3f7cee7b13b07ff90997e23ea6d4ecb4c973cd1a2e06c1e6d45e7d04eb01c26d625637c2fdf09f8f1820af01494698bcdda59f882559e97cd41df7af773c9d7e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11275bd3c2371c44a695c488c8001defaed054f88a5510073862f07a43c1bad27c7b48ec81b4d942f2ca4d5c5edaa41f339543ee0b3a038e927f6c0f811f9c68df6fcb867da60fcc54bfff3768735650bec237568df18d10bc95915;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdfd5bb5d5da3010bda5d8ffcb5ad428b87cf94b31508c6384877af887157e4d186161767be4eebf19822423248dab692e80a18733468cd09ac7565359a3da5dd7e56bd6c10e42c724e973dc9be8543584f4482854d4f2afd9b35d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce99995365c4873e9227614558c6ade4b1a7382eb392bdc1655f43acdb391945bed547751622042ce9e381d5eff4fb473e2ff0d70ea5873c0ed1103e133ae0f26d9ef43b8e375e03dd597bc8226112c62d45dd70b177f8d329cd45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2343043da0676643aaa78423cf619a35d64197ab7a96fa0036186b2cae0f79da85aefb461c456ca790b28e7e7015aeb61a6e5619ec78ec6b31cbc64a85c10c41cdbaee3e1affcfe6b99af94c3371e81f85d0decbf3502ec5a8c0a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b8d5559bff062f19b95dd3aeef38464bbb1e9a073c0635b06b6c7ef7e265afbfabbd4cd58cd0d10de28bb2fe4d47d9e84c89e0f18013f326347ad49db2ea5d2515428f9e03f47fd8b6a174ca60321a1e1b6463078ef6da83f0b03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83d9c231f93e3204d22802c6bc1e1b422001528fba9fc54512af825b53f7257f3b1934ec3ab7a86b46f055239d438d5d635e3e4070a88e77c84740cd2b4424ecfd4d2e42e7ad2c2808a9985a0888ce80159a26b6c5cd66ce25f0c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87d474939ab711d1827b5a8cca5e1b8c9158d32765403433576c82c483f563b09fcbea995dd6a9d325fb101193091aa5b207eb4f3fc7f98f2c5a67b996b0d02f17cf21b7defb397011e351735644c02242f30422f5e94cd7b3600;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d257224cd0fbdc1904afb3bda1880df0fe04534e163fe8c950a9e50a31dd18702fb5215de210f7d666ee7d9be78aa6bec2117ada3634331275f80cfb9356bcf61f40d12e71b26c4d1a470ec0d6662d83de7207c59c58969c4487ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce65df9c86b821eec3135742cc9f0e45522a92a547be9428870f56d74e85157dd4f1ad8bc55eb1ead0f64b9e0b9ae96cd8ea0486a5f1e8f79774ca784982d5aee95f5771484cd7fff18a8245020e72c641dac09b356579673c6fc9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194b2cd21fa98abea6cd4c5f0fd368fb6d118fac2fa6e72bac008f6b32b7e71ba25eaeae5a10baf063157b7e45e16980b5a6f25c0f091ea90ae470ff1a4d1557b1bd6d520310acd912eb6aa47c304b10d067c1034780f3e5e2926ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c6d3109d704713d62b81c7ff423aa7071e3b377a0e2182ca97270f1ca450db8df0f76e5645fb523e382ca7cfc3fb9f646691af04ca9fd5b5589b23eb1277922c1a9db6b0601f0dab80141493c2d9209665424cd44aad95c07df22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63ffc21e25690d7815728fa557d06929428d6d23063e585ab8e784388ecf68fcae08969f72257380bec9395212e63f7a724d3b9038bbc6187fb91be4ab3a803381659d4c6074e2bd94b3663fc83391a13381218c0fc08b0fa81b3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha940a48889f4792cea66bf24e102f165b3324867eecb05c04861531bed565feae3837273dede5da789812d9e7cfe5fb617844ef78b1fd9892dd7c1b739c1e97894d5f8af5a604a567ee494efb2c43fd3008c2ff24db31f9a32dcdd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1152e645d6db29178970172277e7e2e58da66f62e10ea97ad55ca5336536a4f3467c62a91509d0b03b308c5e574d2b4f46fcaf709cc688157300e54075b708b5cd30dce1fb7c5e62a0626b9b9c5f7e8b649103c87879f123d8f73cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e6baa7984bc6d3e17ed83fb3f0ca5a2079cfc3e6c061ac56742f580fd4ef090a0b294ef519718efac2381aae6a5add5e064540fb42aad64d12fe915c1b5baf1b82a5a2447d2ce3fd0f17bf854c1c38ba433585e0cfe2b8ea7a75f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9c050ee526439658d78c7b9e0e223e6ea1e8f436333233dc622ce6fc62ebe84186035c00354a6079afd39f5a2c883e6189b5ae65800df40c65b593ac570e05d710929f7af725f65e1fea90022849b0908e8645e13cdbfe74f89d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182fee44f3586f2a8bd07cca9f815005c4ec4667bf1cc3e8f1ec07c36dbd83adf2b542be7e89a572c547b48b82fbf3ee4ac19f3a55f9246578d63d3f32881b4417d4c917895353ed255204bee7c116c482478154e8a012398990b6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b8e51b30f5e0b5b55bb7a92fb1253ee691054283e647bb59160c8e9ff69593b4f50bc90f2f608de625c5cef43b89e83b505b694c196280e3e92846199a6d102820abfa96931f9599ed4acaf41f2f63f2f6e18585c03458047786e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1991c050f7a7a953b9c7b07188e5e92885293316d64337b1bbf0ee9041b403c1a4239363a66bda467710eff6f67ec73b4309fa1005d535c93820e0eb359401d98bae0c3125f14f7426cfef9bf4603ee2154fdc8da12a997d10ce8e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4518e46070982f2b6d6ba4760863b8abb61100700d15b4d54f6146c1ea985bfd1b4c31a5d898724991a93487cabe90a1689be1ffba328bfa1f4c7f8a6f60cc703ece2ad0356b0a70bf93d971ae336434ee8c8437dcd6bd77ed176;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122cf566207a93cc21f94b8e4c76e3c496cc3178bbaf5c02b5068909ec4f8bcc2d25de4c58c40bdb0c8737238709b4bd0e085aab30fb90a7a7fe6f70610ab702a976f9f26d42ff7d1b806794d84f6aa551725029dda88b6a26f5295;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8bfc84135633faccae37ffc6430a78020d565dd9d3e3edfcbd39e1d4e7abb6719cb3f2b64975be3d299b58f7d109f7cadfc55903564e74c0b71d9db9d0d5ffe5ebf555c34d84bb4e31c6fe365622c7fe501f2d227d814d7a19d75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69470a5da5d1c3d6c77a9d8cd2e4334716d55f0680a44804c96e9e9d965c965d5527eede65dd7798f44a7a46679a973fe45f6d8837e662c3a18a8e7e08c01c043d8d967f1526de80e268124fef5abecd9f0057452c74643893b697;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e73f75fa7dea28f1a51c450ec4723e18a495102e5e49c4da4fcff5739e5f626826a2cc1eda20e63d6f80177ec701d0244cd381b5d17b6618c1308f604db15b62206e2d5ccb566681cb76692ae960434b3286f1d6a798ac9ad93943;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193c7c7f71c40862473766a4dd75e572f4a42f0c2766aaa867db584570b0aab354621b7e1526fd4eb1278d2d5bf8c0ff423153c3def239aff4f7c19c82ab37cdc574507c88db6ac631c2c71949f253a55b74dfec765b68cc783adfd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b804bf348bc534dba66d1abc237c1e9f65b3dfff80de0b0a62155aa1e4fd84067e41c72ae928d020826531ce60deb8b6a28dacef6e4d37ced715d5a96b78758bbf9668f586a16b95b2b29d4e700ab5a2d48034c5b0435edfd3155;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8f1a94aa08a58e310a9b36cb4a9f1457761a986a6ce1445af416a89667d94091017040037a037448425af93aa52c338630dd2fa6aaed33a5f0828f3186bf01ffc88b432ee2040a5a0d0393843a7854c9a478d3bb99e84c8b01972;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11777c46221665dfc45d650c9b27f86083612aa326b8b1ab3fb41323a6b2ba68e5c9167e4fb02069bc38cd4eaab4e533fa4184b9b289ffc468f0a4e1dc1883a6bcaf63038d40c27792e497fdd0c21f9a6a7e1002b93c0cc8e4c03f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c31d20af642b28ca6bd05d76f7336aff7f5c3f7d2cd73c7f1dcacb693925e6eb988787b3b98f934634ee6e455a4f6bab9903f8b2d148e2fba6058064cee5e43281548313c214490341fcb8c8b6a521b045105e7eaccff6180ffc9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba1e90aca625ae6484686ee91b0b95e04fde6f7b8c3a54aa1242af0d86a251a84e31690eba88abce255f5e6a69fc80aba4c2f4f0feb154964b54720ae1717d51ca7bc099d22fc26c22a2a7f4ef245a62533456d75547825cfa1521;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f803c819119e633e5325eef87fd510e4702998e9cb06adba0761edf5dee3035a957a9c97196b7502365e3426342975c979ee5571a25f7d343d5152b9ff1916af4379681838c203b915add74a385c782e6440029159524e99f8255d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf2bfbff793f30b854e29c0c1054cfe18655fab5ce678baa4bfae63f43e70273d88ceb21e267128d4240d4e817b5e17ab25aa2529348503e3587b9c0dee515e2744156b8cd0aa964dd32ab88145fe7aa02bafc6bcf1a4a59921330;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2765d77b98a29f94fe77a6c593729666a6218f3402a9e82725e09286b7e37842d2418c92d6f60f66597afa7071c12cde7aec307c29546999258906d1b0b236dfc13b4f4aa0c625db1ec377b835494d0beb2a8022d0ca9168a8686;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4852e39f76489697a909cdbcdd8c42c46b6072abd1ccd0c60f4a135223226708f6f614971433f8c64cd3ca1e1253b7870f4d176d7de1c42df396bb69d06a8cc3b405174092e18338302a73d919b0dd6fc61dd697b0d82738be327d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8ae190c0187688cd5d63afe0094352bb401839cc97185e8a6552a7991643a8f8a393fadcd7a7867ee2b198bfd91202d9db9e09f7fd2736cdd524f7d4dce00347245df8c4d18d1ab8503aed2c9e28f2ed21edd6a538d25df7045e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda0af5527e9807262a57f34da592b95a0eace142e34c7594abf57439fa5532584d74e648f65863fcde2a26dfcccba838ec41ddd94a4cce060f81d50c8cea00ac501863ac48085685f13d1508637a7e3e1779c6507051ee9fda607f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c662b9a5f09bb1f6e25afeaa51895e4092948d8a6ecc26ceddb3864d2767afc8c5520714d23c375961ab828c86a8712f5cccf81ad50ffd41cd0822b0a428642e0aa5859833bd2da5aa3f093da57a509916ca9aa30384f00b2ca5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1333fbb2bf6b19d3bf9a6105aca8cdb1ca623aa57e744911886d1fc13c48baa159dcf092628400e7f7de6c8a9d9d5781b9feef243ce3d89d8e87a27591c0cc115d2828aa3339d77141e5bfe206fe587fb8c06fcb520d3fa6daf78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fc206e3eb195696a6734245d398a4357f3389f52aaf47e257142c3c27b74edf2d8ef4117cf71ffe80510de7a1da0dac3fa774f8e63b59460b170f2f158a543767f6ab1ea80528f64899ec059f63ecedb115d24d60c499b2499352;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f55d85ce29c0b9e75c48a2a7a392c4551fc19a9701f843a325f1a3e5e58cdf773e0b6e44c1ccf5c511f2dd1129d60e3776f708b14c318ee4e50883498f49db46fcbaf162a082e68fa04f4f943bdcb7dcaf8c18d6dd41c947dbe72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0485a6dd31debbc92f3ae74cc901824631a94502a69b6d6aaa3dd5b1c1858185efd353fc2397c34ae4ad11481f9efaf9ce0ef5b9354534d97f7b1ab39dd9ede5bab4cf7e26e8949f59aff0d777b0a29bffcbdc53d99d572420c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177151ed400c4e35fe4411ea161fe1966c949efb1a7d7bc1c8ae0c1925ab42df8e0735601dfffff84d188ae63f90101535aa6db2c790e609ee0241ee9f03b923815f6d757886e67b962a61359eb4822868155a5f29848ab58bb7a42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18302a416f8dfe9e4e1c8b905442f19dc936d46738b5389ddbbf76d56158bdaecfeeb8674935ffdfb8722fa226814adfa4828d552fc79daaa06df88758389e10cd4c410eaafd37be150b7b776494a32062663696553fa6839b0bf2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73e8a182de28d71431945a157c79ad8676a52c3bb6dff8535ca4ebabd54806dfda68f756ba710adb2c1eb92856be8e889aac7e961dd1c8c0f136bcaa43117b071afc47f3f78a1c4953ca9181e333e50af2c827a113f32cf35b2319;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1476b6dbca9765228036ad83803a4ce3feda4bb2885fc9644ab4fd6337a8ea6d77850c4f4a2d24c56de616a95956b7541e629f6e151c735575ad0d77365fdb9eed2ffee0e2e2ee1ee3c970a79bba18fd0666e1792ed204185635803;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf68173ce1c7c80f69bb2ab86f6c9b902cd213e159cd02b061410c6a5461896759c22a1f988a3b993ba502106a83650220fd8b0d843f8f8a83e015471532229a2c4c5bd45cc8997ec5fb4e98b9059f524fb4b7ab10abf5cf9d147fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17235708ab7f6bdf3f33819bbd544a64c49364febbb4d19341e15bc50d7dbd088cc8795fc6fa05c7a68ea27db9667c6e3f39ddb53e2b3c87875729dd550ab977e6a96cdad8fa092c51d4d427f014f2e5cba86f30ec03cef5a3667ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98a8be015ddf6c1574fb733a2192b6f1ce8153274a760fa0152f962346443ea5cfdd22217755f7aff09a82144fbe566920f5e0b204dbe01eed2bfbf5c75f3de5bfb07e488b301808de69e4ed05ff30375bf68f2d53aac789e28293;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3676c7721a5abc2bd754505f924629d127cfbeba8d23c58037b6e531506ccb9fb4dae5e575854c7d603904ef92dc3a9fa5f7eeb4604fa50bdd2b9e50cbfb1685cd00a8268c8dd450a21f8deaacdad5c33ff7dfeb8784c7888390ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fd57a31bc69341411eca7c8c7e38029c9e326f51156340ef2c78a1baaddfae1e83fbf5e8e0f530e798b218912c5b7b409080f85db3504452a9b9e7b1f1f9731e1cbfaec036ad0dfeaa0a5edc47fdb4bdf9afa2edaae2eaf17b4fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1095a2ec8553d15c69dd08c4ecc7c4289bfbbd6beb929515807a90e17ea803bece39b217065aab6f27e465ee214159cb1bdf089665f8d218f68ddf350d9d7e008023b1b7c7b9776c901a04f61aac591d7994175a6b5cd8d2b8d0207;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10114c0de3878b5fa25083ecd9fa7fed594bed5ff31a8ac0d43144b3cc787551f642e319c895dc758443743bbe8fff4a7a8104693206bdbf1946783307bd3254164563ec26bd8e5ee332675a492524a20626f5ab32dff73fe04a9ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f4365a5c26dd836a15b50e282007c13c65f53267183d7556a7eeffd401340088385eed6222dab080fdbd856b4a34443d2a2f5b73d6582583f36125c36ab0f5986e0c38aa1fd3c69f4f8d8b42caa8a0d526f5fcfb2b90420fe3a2c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee5e85d76e31a2860974ba3a022cba261c7381dc93b5b5962d60615f1c14f096036bda8dadfc79a031a4cb9edd0139d6837101219267be4a2c8f0ecd858b8fc10ba4971b284e76bc3326e0491777d041d5e780aa99b89d6c9606be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31140ca25557567694d2f7deb6ae4a59c1aa16a7152150151efa3f5d05153bc0cc434854a16b5e45e475c3ca306c673c2207dc27be967d6b0801c2eeb72543cd558616748beba8e48268407601f527bd88a6cf33d47c7e7a45b860;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1fa6a69bd12b786652a9850304f06cbe0ed48fe2ffcb166afb1e9f62dcfa8f276829e97c012b19b60e7b2046c5a4b0dc1541e1cd1520f339401ce04bfb6aa9a0db61e51152d8b88e73fad80dadbfb5c7cc4247b04a7c486b4e696;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15faeceb8f93fe9ae39fb314d31147d6ed6df4a08a02c20927a86cbcaa5a71037365a76f71addb74f3cb9ba6d73823c3262b7fb79c4029f463c4caf453eb537c807876ec7fc08250f91de6b4f2285979fe7264ae2e1ef424aa0188b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3bef3a24b5e4ec14aa869fe8761e65a5ffe07031800a3446e6e17420c3540a7fe2759ea9aab1f8824e31711392684f08f60d0eed8110ffe2144ca5941b539a26f69d89be04d858ae3b1ea75722bb032cf68ba830b4274edd5d339;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc13f2f12e720922d7c4a40b133c10d50d29977d2fbf55817ed373f149d6db4b8e5deaf4428fd3d10a2ca2dc26d919cd04f64bfaf2559d9b755af82adecc4443711519b49308440c88800df6c9df7ebe69e56a208636ec61e6b079a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda33e94635bdadecfb6ff72eff999c99062f4c0503ff9587eff75f1ec26fee12ca5f901b7118e69b07b27b1e5b49f44878514eb1f0250089867a11bbe2c3377a6ef7957d224dd0f8f53e6184033823dcd2878f27f0fe151cb2047f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104af16a7d66fb5d79faeb488e44ccc60b897d075634aa052383ab9492ed310ea2783a766da5661f225ac902049ee46dabff5f43421395c48b29bec79d3036c6926ce3cfac9d2723399a5c5d230d815d585d4063e459d24dc07a6f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb2985ae31b2c8a0000a209a49dacec72bba529a890e1d6ac916c4ce08f9cb6b6cf44ee5fea20ebcb6bd0e9482ed56fc79a5e5bd7782899b854e933e91817f152ef7297438ff1de49412a1ff9f0565947e05f2b4f400099d5884bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a1470ddba86b5da0c2336a8d6125a65b3d1f7daa0697a534abed990b3cb626a9d37e25a721b5c5099e6169104cd3c5d9304c0180d5376b9ee74fc56189541f3b62bda58bd8a193cf912deaa0591d2d61de3880d47683a6377bd15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75bf5e748e616e079f7225c6f30113fb8d4e58aa27b21f35d03aa21b32fab99708c7a0f70d69fe4429248ccb4cbe0969d3975e8c8774c3f1d37383f1e2036f651ef648e46d8b0a9fc85081bb703e013635dac306bd29382e4354ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfab4a617b33c0906662b12d76d635f448f34b0aacf45883b40dddf36d3c405d93d57ca49e7b9b8efe0e15443c18b5a41b4c2cd05d34ace7d82a0515090f0c4f2292aaa84546e481ddd2456902a8a2433ddbb787969026cd896ed6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h800ccf64cdbbe0a128cec0c756ccdf6d050f2b77b5e9ab05c7031c7302289da40c32f7ce8a8e9518606f32a1b3d623fbdc3e6bd0f77147b422a675ae4bb0a1bfa6ee71d914f943b120f895f5bd24e43a3345bc82c798b99d597528;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea55f1550a11185ac6254474f6e84eb2dc126d723195d78be32b234e7bb8b1202d32972d6a66597677a586eeb217e4bccf00e3684301c1fbdd5e3b7ae05729655d8058e1a4b2298927fcdd506dbd1a716acd539dcb446d23563791;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1662c3c5670c6657f754503aa72671d95f904debcdf3a2a82f2fab495018d68e65da553ca436f8307191f2dc48be884fa1940e86878703ed0ea17a057a356960370c4c1e743e14f198bfdc200dad980169b648867a2170e8c9720ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10762bda2fc39dba35b79f75e8ce3313887186b64ee9728544cdbfd6fb6d38cd849383bd2fc7fff2edca5445079108d57ef311178c80e775b68285572b155072b94445f1c7b808082a526807b6f824f1715f7a42de555e451e76ffa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9aa62ddb4931730ff01e4df87617d4d115ca931a42ec0e70a0d96b75c59ea1db2be99000ff5f9371c006d8a70220142d55e4568e3768eaf9ae2a6efbe434e3e1c130e73742e540bbf07f5335977cf85921252b126b09548f223c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d51d4da89de868597c56b425e8288e109360ec023d16f47a2eb05d67b70b991ad6051104ae6a00830f7d4c6499840acbd67757335119ec17af321d167a8017c7683603cabecdcaa89274df8b93740a169ea21ab7e65a2b9ca3030;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f0d7abb51134b84e7d07f7ec382b874a9e8d6443ce374316f660460be26bde23e6f051ccc7cd4810e8c6701507d0802f920f593e8665563af83dac68f581d333e22af3f246fc55dde0b3e8ee8707b84fa4d0da5577fac075aa88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7b6c5cb6d0286ff781dd0c50a381cc8a53124d98a60f8999b008216aafb11390e5c544f08c579c277c1eef2be3e8c6f1ef665244e2b6d0df6e4186d0b34077477c4e2b2ec1a1aa687a5b6b6914a803a6a778951edefb80fbbed9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caadffbfa9b4c9a56c75bf8b064d1c8fc32146dc2357ad4bb130f411d4e7ba91de60593f6cccc1b47ddbbfc0ad2764ae59f99069e30ac8a1b9822be57bedbb96207814d0eff5ce3c1c9aa66b5e33564175fa37e246c556128d7119;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7745024c6dd365dad14836ee89ced4d9d49b0a291312bb47e1a7e3953000704eb023be6781b7441b2fc9131b17831db89e4b5c1c81b03fba74275a2d71e885eb7a189e6fea1a16844cf029328f812c1092399dd9cd88c2cb4b2a16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3ff64139e93932d33aff50ea873359f0aa5c0f18464bcd93f8abcdb092b29fef05f333b2a58b083991dcf8d0b65284418d33e4861ad93b357c1b9b2d7b0849f5efce245d1df05d898f27b2f19f2c92b598a316426c48c4bbadee1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1532125f5a1406521ea5c49b8e6d39f397631a0365779d761fb59b9917f95aff402e5ad5a7aca6ed86fbe109ae0c16681ea21e94f6c32c984f30f6d8d2aeb11ea9831d7d1a14dfd0944f03cc5a237c265762de990e470ec5b97c701;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1ae73cbb1d4e71e95e6c1f02972a296fcde220c5c0b529e0f494e5713b9cc34cf89c8a70defd8093e5d0c51f6b8184c8f2edbe0e6207f9f4bda46f7388bdf17633fa640fc76854ec22f10a3951adf50ac8044f803b076e4aee45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170bd4fea3d468436ee5e18922dbc98ca9448a373011c512792f70ea60d4baa567836ae9ba7585c15569f8496a6cc2ed8dcc31f9da5b21378e99018ad6d2a530ca0637f0603794cdfc5620344b77cb1249abb641cb7cc7c629101b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1e9f768b2b6fd8d8d133ce4ff3631a0d8e8acbcf07dc1b5c685679b0f414b8bd1cb4d0c061a053f08fbabeeb75e21fffa34e7da01135a27370ba8110630ba4f53c8483364b5f6cde88e9469810889d776e5d4c44058fc212670f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae9caf6e7bc509003c07e2e44d2a5e996345bb6698a22759d162a3c2df62b496da723488582a1f109700bbe46e4a50f4e7d1927069d5e185833ed50ed8ce7ede1d7fdeef2f90cd3ec0a4e660009bf04b5cb62f0ffb1e2421e5d5ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0ff6e027fe5ac5e34f578fc6b88e2e9d3ff0fa76187cc56d798e937c40157143d0d58e7c1b6d0eca4af974a32e1556cdcff390023fc135d282111278cfb3a1ee9598671d82b6b5b32e246f051eb61e8c722525b1a7fbbc5472700;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17702e27856aaac78d20f977736d6b2d02c8161d6987885f45ed5a3b81f33aece49d2e9f4a4f88687c52a96ab92e8e0224b8ec3d63e611e7eed516a1fab4699bb6f23b7734afff54b3947d3bf752b75552335efe974f6ad1119197c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h431d738e4bfcdc9251a339325a6e7af4280e0736fdde1fafd454835dc48d0bff69056065f28aeb745d3c442f2c6d37b21354cb4b707f73c3114adc680a924c173f12067794da36bf2dc42399579d058334ddffabe97d18b969b848;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d4c0ff3b2ffa81a1f85d1a93d7a1597fca80db785accf2aa3838f70b4723d7fd7c307cdf7d88c7d30d3fc74a28039daf5c3722583eacc341f9d1da5b43c4873970ffa35a02e5f4707f7ae0266b40dff2348b4ac52b7a8d1dbf70c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb15e19e0a615f97c9d398906b2fd5de0459ffce5deb008767496f6fa8d84aa761c35efc8ccc9b114d843b102ee45e58dad88bab016d113c3bf0007339a02ebf25650eb3a584e24964ed22029a8bdfe2b69d3f7f4f73bd0955e4ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbd7dda8c02f82455f446983c85df937a662010bc8ce4c3ec7b2610f8a3dd83d1b6f62653c18b8f3400937811e85ac830834b46182c6d2bb75fba136e0b82127d9ca73af033c0b150015751ebac040ae009f27c98b4e7ecab6ffe0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee0222522584c8c19bdd3462a340eff3fb58f0f338f3113a490874f4b96b78ac44ae792ea6d2c539be1d622e0ab82ad01c41138eb05cb1d053d656b4b94303e5ad8093541fc06fe5f46f86dc6f2aa9fcf40aa994f5e2d3a5163108;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h727f215ca21807c90e411c4c21a81ac6b863b223c0b6ab04604b6f93aba5dc2bcdd2545728ccaec303734d1a16e7fb1d3729d12b820b3b27c028c691bdd4b5ca5afa09d7997a20afce9676f9a13524244036f028e9787c61fa8c7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1993d23ab2f7238c9df25e1a0f8956f0c160d09d34d3d33a0ce72bd84ec03a434d468cda038cce13d01a54d468c6b14c4de4ee6cca3f47b75299c722eb3df82cdf1f42c37a55d7b8a9e083a1c7fec984f511608051a3f8419b9e4c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e12219cd48c637758fdbd894bf86eee30281ce6690d681f52f98b1be37e7741f45e1f50f58ef4cd7bf6e019287530100430ffe1123f13572bf37bd828ee2bd73467530e218ea0e24a20da4763fc56f94b15fb1a84a66fa3ca926d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3d4038cd8cbd777c717ace38860c10e827e9c81fb39779e56c88c2508dc2e1d71e187d251d28dd9a1048c62be8d73d4312e63adfa04f319cec2dc3a50566bf2a06df4e91bb72521090575f0568380fcd56a5717d1352b4241442f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd7d3d4187f7004d1190656bc17121509ac4de7c27a2091db28d58abbd1e81160bf2b849ecb2a72f4caac87dfecbc5324551970934b00ee18ae5015357473572fccbdebcad40648a362850532d3e2e17d15135687e73238971f398;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1691147a9559e1420d2d8fca5b3e0c6df8b868850caac892bd74e22c3e8c5094dfa5b94166dd31133677981ef431e3cee2d747b2dbcdf4bbff8e2a6b157e4915ad4cda666acff4012aa891d8ed242400427d025e211c7cd66014403;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd28871f0436edbac6fa8f7f554dac1aded70353ff7d5572c68dcc4699f33b824066e4cdad84513e4a8988039ef6b85b049bdb0e8205b3ef20d8de33ef794f89152539e5a8376abb9a98bb84a85c902ec42d13706699fc21fc805b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d71f73aa0a5bc1470fc23272fb591616ef6149e6f5203d23c0dcae5689438942dd20845b2e99d0e8911820b5dae5a5f119697716273e5d06824bca05750261c5f40477444c7fe84e28d2e6a48bf74ffb46a4e6a60577271e85266d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1612d421f3c3e33ead884110c0b93357d2772d371731c1466a669fbe1f077917dcf7058ca86d7949ef9055044fdcf28567303b8fdecfb06090b198a2e6cd61a59306c329bf1eb3b9132ab46a17377bcf56fbf78ba17da6cdf1d9e77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h278128bfd1aa21d219deb6e8fdfe457afae485eb2c6d06de9332be0c165a3d435db6b40475d93fc73fb041eec02b2e37d5fc96bd14db665e184a9b7a8b70947953d3bb412a8e786f1db5f8700fe2568b3307c86a14eb0dc949b902;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2986e8a9f97b14d7b22fcb63aeb1818e0d04211568520a8ee8705772875e25bb84a3c40f38fdc082a7a1ed6390273116cbe94f316c9731c7cf957feb3477593287d1a47f5550d7024339d3140043212e3f89377b4d93f1f1e5b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33485813fd58290963f49b3884704e54ca353e264e61c545cd6612e3136221bcd7b8088246dfdb375603a36d18acfa9cdfebbc4a0716e408401af8410c3b14012d78931d0cfabc897b4a4fd3b1ce4cbf90044a0771fd612cf7d8ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9228c9901d5cd920125b51ff110235bf093d0a5952204d7a94c35e5d48325ef8ff23b7632612595c31d38acdb66045c6233ed05b6fc2986b61c2427303ffc7eec3b339297313dcbb7482c1b621ef2ba34d399e0645e09ece1eb7fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b0fcb10856d2b57a6da975e93315b7f57d465630e75992066824c429894ab242cad04f5ca0db1019229c5f982549d4d68a8a9eace86e1f61a55a9e1aedfee043ed82fb6dc50cd1232787ab1cf830e195c55ca921725120a6550b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4195ce55622a35ca2c4347fcf8c3aeee069e7622000389ec7c45054a137ebba39510e8de584f22240ee603483dd5bba5c27723ef71a70b6daf1c50dbddc92281b3baeddbc748533e9e962bb979266edbf795d298540634b9ce5cba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17589ea809b20819148211a1255ace4f8b2239dd743ea64ec8f2f92ba85054260803e87177aa868285c699bcddc700f0dae8e529b5b0200a3193e9bada838c0928aac1a5bd6cc1a1c223e5e23288754c99a87acc3facf659aae23a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2fa3a2387e148abc4d0c304269b8eebfd0d8e79604f018c01b3c11300c55210f33684173df2a663120965de4c18f82f831658949b2e6b9824ffc3c64ba77e5ca3133d44702b8ebc8cbf7ec7cc9fbf02bf5a1ed53f540a5bd58aef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7bd33884c4ec3fa24f89c9dda436046bd1eb7c85204f91195cf613367d9c79d0ed942d3a86f81e9a69b4a970c4de17cada737005289d1baaad98adc591a618d9622d85e1b0404b90632005dcd5ef00e15323ef9b11b8d01f0a0d16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba1e9af2119fc034759b4db0c60b33e5eb64f521138af8b8701b30f178526c65b82982fc64aaf5172bb20da27a7381ad9a617edab1d9877ba6055d96c410576b7c585a9e6b6d5bed7f651c829135c1712a59a00240933d88963c7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3872e8f34b2eec66756a7bbdcffedbd8858eb59640fec2bb8bb7d281519154fb998a44fc647502ff8097b36499c0851b22394def76f5f812b6138f2ff7896ad3a3e464e00735e27d48f71c3faea66c4f87117c2210be02c89819b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefa3a1c12fe41f043908270a3a59caeee2c34c22f60fc843d409770f701bb49eff2a4edc8fdacf33886f676bf6b78fed8abd1ba548f43e12c0f2f75ec21890a4e7867c51a201ddd4e25637dfb077973a940fbdfd81ce44dd71195a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b0638ecadd34ca9e8d2eb5b9986081989be392d6c7456d67c0874529f2b91c00e5efc2249fb007c8d3db6c961c0a63360f6109253ee3600c803c5d344e0b19c94bac4784c1916e9c00c0aa17de97aee818aad971ebb11b2761040;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2dda7e76da5437f99adca8e401f314a315be48c0d23044b3fe4cabcb76473bd17537fb41c779b2b03dfb9b0155957bec4daa423de90d21047a041930551efa0e381a73fd8967589a0cef19092dad6c27fce66f5324ec316a8e28f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h809f4a1e27ce7be5f9317e8170ad427198a619f65b75f8833b5f41f079876e31d039074ea155ed22dde77cc38fcf05f2fac20c1a32aa3f4c407d991a646b932eb09bbf44a6769c67426bf14cddc929366171359151c0353322575a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bd617546ed3374dc85d55bd4f9845bb34bea15adf2b4a2a9ce9610d4cbdb28636138bece45b44873994fd17439b1fb8d9842a16fe70dea28a4fe6c5391f31308fa2fc76491333e6b22260e9e2c239c86f6da3efd2be22401f27b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112485b32c35f263fdf97d51ab6876df653610e7e4bf9d321582a5757440bff6e96b262de2d1ff6771a8f00c82568dbea5eb6aa074f5cf58c3f107abb88a29c04f9c4339fd12a62dcd05a30900acba2592ba6a7479803892e88a65f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e3f270fa85706be106cb0dc31cf845ea067107563362daa39a0a75a594ad4bf2fac5737e9af68f829949ac4a337ef55a1daa6ab71ab509ead21234879f31f79921eefb3798302ca819c29807ccd0bd9f9633243af62e8d98cc376;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cf0f15433e40d2311bc7c5a4c2075448f68d4fb3e13803dd442f263d1ef62565af65bbaa82a386865fd3edb6a766c312c7510b45de8adbab396218fd6bfddc63b8fc636c9f3ecba666b8d031c1681d25b095c3fa46d78af1dd2ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fccab059d1d7b44f5c174f477f40ca4dc1fba5907fc398d104febaa8d4f3eae22e4fe4983c89568b8214e92e6c1a0b6cf49c050ccf8c82cf3ae2f523f08672693870ca8d005645f68dc7bc054aadcf30ce99850f47458df088053;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cd0a5babfc6cfdf8da2c35dd919f4bd89cc354841e90016f09865861b782a4c324ca715700da5564c09cb5a9b10c4c907ab6515607fa9fba1674b8c1aa70120b994942e514cbf0b399f383f1abad33524fd3b29a0513d799cf7aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b957d1c4fd49619580bceda6b1f99bfd0145b6aadf361594c36127899436476bf89ac8e65333c10850c86a65aa4cfeb9168b24016bec3c46d9ef76eed812eb4e03a0b9ae23fb3afef986aad46c6a77b2a286cce4940dfc7cddbbe1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1347f53debc4fd6b9da5b296292e0b4fb921570f7a364ebcbf1f49ee1969ed64531136877ca62d3ab08174f99ff595193525c201e4bdafa8c04bb1df54b760b47e05e9b93fb2702ae24bd578de83322d3475ccc3c6601862e4e9ea3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he106ca848eae3c071aee88f96f6e494127bc27e1b8ac9ec1e5cb4aa822d6cbc53ea306f27742a20dcee434416b5cd56f399c15e9259c9d5e1feed7a62af960d22bf60fd5e690a6822c257ea4e0d294fabb4fee1cf91747901a16ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128995aa203ea8cc4f2034598fb9ebbf9b2c79228d667e8fa1006324faa238bf978e8fbf5397ce387eadc8c74054a68e3d1b4f839b89413392d35e8b292673bdff8076e7fd581d9372331c09e9fecd255482e943719ccb84fe671a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5aa5ac3cdb8fe2b31eb9f8e062d9ad2d61f684b6ca048b1d0e5e512916044ceb72ac826aeb52cbc7f7a629fb3e087c2bc14ac82e3a6d7c9ba7853a8c18446b29e22e39976d20ffee895fdbeaf07a3ade5e0b3352d26af71a105d32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18db40b231213eaf0f8e3218ef30f892e38dedebe45660fcce1b50d34002f8ae11ea88b72b852d32af97a15accdeb49e70af8d3431793731095100934227c21883746b2c52e88a71788fbfc534fa3bb73127a479df66466a8843a91;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16008b9d99879e58c2efdd599ab7433170456d198923e114805a44ff8cf03eec8eb89bd97c7e79593b0b65e45b81e885c412a412c38b7754819fe1276f8c6457e42e2a6a7c83fbd6ddb853dc0834969925cbd6c93aeae1531f3c3f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29fec463b35d317ff5dbfbc23a9af091975fea28abfbf724c4361868b3bd1f1578dd3a53295a715f8b353e9b6932541f5d66fc9f571954c75a5a6f2eb4fd2402b33fe100f542ce406c3367c76c7710954800e84f8ed693e3035130;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef02196bbfa01869391c81fd279842e49c1c4776a60819649066c6d39a9e073b4ecda4a3d59297fcfd2a2e9eeb61c36246913851423971a61dcf379c3529cfc0e0ee1d1215c4efb43de8802ff5414af821811da58e743a91fe902f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc7b02f7f956c5d248987b08816fbea3a0df58f51469f1df83e65b214b53ce4190735efa0e5d54507afc67df8bf93e02f42f96b92a7f0b056f46ed02d2f6984f94aa893a4df8823942db598ed3c739e34a2220f7548f6adc6d1d01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb86e299fa22800763bebd3b391a1dc8c4aa22b31140d174bdea58bbaaf50b7d89ae7f8f274ae0d5134b373b40f86f9b8d1e48ccf899856bbde1a78f27eeb1a585cbcc964f48c62c80bc0e7ac6cb4a9ebc575a58aff014f6417825f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h897ec97df9b7738dd4d8887d2962320d8b7f4f7d555e01a8d0f3ee9d8f01b3e116eb8833b987001bd06c130d741dcc0ff545cfbcb81991f5e5e76e7e11343ac32601bcd85a3899076a4bdf58d14783d501e979c2af6c1981c30e08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123f4d2620e110b1a2400a7443ee828f5ae2d27579d584f282ca94fbdc89e16999ccacdbdce2138b3cd0a56c8e7f19559b5f354d9fd15c6b832788bc3639a6afbb1174dc6a898f8fab7814a48866efa7ad0132f0af11f3ceea50f69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h940e8af982bf85b41a5bab7880d2447a4ff5a40d7ca8e0abd5b0d0ec97bfedc6160250c2cee764ae9ab82386ac7c0031ab99a1b1e90081da2162d1c5381c0e501605b5c407323f1a6b7fb68c601db158e1ac4c2c90424138321680;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4599e0f8da7723d53c78ffc7e35e102a4d77484b1980cffa4972cd0cfcfbb30dc8503919b200a9c3c923ec513e57bac8866b24854bd3e8c69abe96ed6e73e428b73f342ee68cc3cdbb9603c959a56595180dea480b46bf8bb9f212;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fef03f1d3480677109c5320b13575e4dbbc4ff55555a5fcddffd27992108ca8f6c9891e7b3d28493b9031814a9ddb701f7b4047f7f12f76b58b8e7eaa9cc9a9efb782fd1027c2558fabf16feed7cb5c6de2947edf11c6313f15993;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8725265e5a271263ccbe7116afe38e45dcc87372d90b3afc34b18544eb66c6e96e19424bb3229df0c51e07031c5e63e15509eb0a1b298ccdfc52476c2e8374d69e8089b1a531386ba0fd167670d0a0369044894c56ea2fe5a59bd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c240c7c479e49d01b2bf34c652ee19b31d0ce30cdd999633ea41e6c45c9ec65b2a104fa59fa4197cb65651a1a79b99e3c4618b8851d14f2509702b2e791f4588211af00ab1b6f1cf40fe791c7b07fb4deb49f0e74494d0f07f78f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104efea5fcad83e8fd1203cca0ae343fe14cbd080254afd1120e046ae291b6001772cbe5a3a4d48229f897e26a6805227ad8a070a538e35555774c0c8a675f71b94af6aa78ba7113665a73d7c83f0910489c603ec574d002619afd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ab36437613438e312197db338623ec85f268ebda4b1674eaf7dd329cbaf2ad6aa71f6753876d7bbcaf5496f2100d8a2952319f8218e900d0a0e34f4308f5238583723d0ee33b0b3fbe7eb1dda4db756d1f18a4a6d21e3f1e709d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h759773a4aab61c32e3e4b588c0cee48f143cd299796ed4bda7efa286b2b4fd54ee995d855afa7b6ba925c423bdd9ab3422274ee9d3a53d1f43ef44aabb0691c06d8e851ef39001e212dff43fa9021d664e253053336d2c54fd5dbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c6c93b14185a4faee30c01f2a889c914d509a6fef048e1b8146f19f4fd15bf1de5fbd120931e2e68b94c3b5c416db6897bc24a97015e9b18c3010a16db16e3a190b9ad9d315e72dd1bb11b4dccaeead3dee985da825ffcde0a33d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112861a47cb87b18f521ab62c400448c4560857b140d91232bc1c8a77f5ebc8d7fce4aa1855e0bb07aaef276aef5632afd86aec6932ed67134416189e38f9520f26e02bd228c618af36db9ea48d2b9f4a136a26df90cd4f03826a2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2f5855257a10b9b3d10b4cc115f33cce0aa425d5ac4ec19195806f7d4af39d0bdc4ffb57ea1910d626a7b23d9314e156d51af185c664b612452ade75f49abe785005719f9e1ffadb039e6c063b6674f7239d0cd5f2f43b3a8ce51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107e77a54551c91515685c773514882d0d0b69749f26b9f5f343964695fe0340f95e49881540926e98a6ed9e805778f3c71a4399a00d0956edf23cd30f73ec2191b03c126811fc325a1b321b4bd1430758b988920711fc460ef134e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10249999e88c1e4669a2bf444f345c398d5942c7b0a6e5ae74e5b36a578342fbfa3aa7c4a9875b6407f2dde7c69b83c73324d790d67343ad3c49557c9e6abc1b8588e3099919c41b9b2014450a06fd4fe362c8cc3a51a5327d1a49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde555fd140a01526989cb6f8c97c748c77022a0a8fe25ae6d52a2b01875760c89ff1e0e6ab584805d485082b2f28d2aebb222f1dff1d0f8767589bcc6e320d307e85d2b49261107770f35364c454a58556350d0872faac415007c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h299712a40460414ba7200a474ef654ef5ee247570975c0a7649c685f641aec31475d9dfe8583d0d072ec8fcb876b5afb2e3b374ae9040ba1edd2ba252ae978d028d5fc8b936d297c0c0e6a25d510f5a8bdbda591ac1a9a6631421c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h835858dcbb470cec2c16084650b26bb28eba7397eb95fbabe86a982501bb22ffa10dc1e6f1545f1f716ca6fcdbaa2a4804602c143b36e0ff8a92a434bb2e0cbdc9a2437b35d013e58f0f7766907ce1c69bcdbda688f767e845512a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5835bd8829b327601911dc85a3a50f55affe11558c1dc6da8ff398232a78af7307029e1ccf6ce29e1ce25c635fa45c8687a0963a4e098ee31c941de68b537a485fc33e85e98965c83d50ede1a22a2b49f56b5a4347d7e5d34e20fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134d998c6651098523e1fc5680906cb3f8953b63b4fa1a2e628cc8dd4379f34c6e5b9ea5edcaa200d8ba76578dfce1203c188638cb9e99e8041d7f3609e07b03d9de4d1ea89cee615bfa8fc6bb52fbbccecb1c46895bf97fdf8aaf9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffc641ddf8bc83a931221885f7f893cc918e354758310bfce477734966e2eb66ea034fa303c62ad50dfd343334932d03adc52743d93836d26ed17428e290cf0818919a3880f0f52f53d6352149f45ecc3ce6585ffaba7cd2e2e9bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19eafeca21632c85a601563b80fb2e0c4873d93c580048d8c9636f6b859aeb80a662c40eb52ed4c40f0d3f83e1088ec6bc1bdf89c1c7a7880f7f500efa30323bca547319aef7ce7eacd18e948dd56cdfc62cc24c5f6285f0398297d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h472e4fdfaa37bcb54746126990897a0e083dc63d04ee5d00570f0e9ae1decfa7abc045c810fb2ee8c499cb415db663e7fe73c3d42221114bed4aa929969697668aa365117c6f4fb27990b955ae36cbf46cd069aaee2eda2eaf10f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47def8c38df2f0a85bb214385861b1437a6663008f02baf0c0413092bdbbcb87919f1ea2f596ab5bf9120845618ce0742d576f07aa3a448cc8fe09cd62988e8f8f0c9ea13cb94e297aa37e7d4d709177d1e070132694f7a6824750;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3cfe09feb1bd555b8e2f45a498a3c7f2f9dd2a98ca56001032c4c3a36a376510b4ade8bba943355ef57075544eff815db2e5f4d8a08e283a81601b4bdeb1f2f8e6ea752ba211f8d3d8ba07bc30379aee08b8ca7c0a40759e542078;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5009abbbf647d23eb11f2f6a8bb676c31cb1c56b206efb57fea0b4aeca339b4b13e5c99f7f4e9e7cdd0c665d4bcaf89f37559e0f1aa0ec07c74748e4ee2238cf6932631f6200facae89d545a9869e2a987d4937561fe30d23f8fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9237d70b279fcba7814534d3911c45308e915543dd3bfd60589cbb3240af3b01c3b13289b16b0a9fdac6215bf8ba0f0e04d8daf476595096d40b0a0b1f4ac871b855b1a7c67f35236a854401e4ce8b5d37a0d30a8cc98ef6d5a745;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d933a2c0f0b63de618944aed125262d4ef26ed10e354af412efe6922bf33840d0f376e1b8d5d072f7e484347e538d9a65ca8fe6e85d9cd2646384f911c875275d27d179fcdbd45a3a5f2375491ed5f5d5e95b7d67890b6630cd176;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29bde2956102779e72529fb6982ffbb51f6501d345cd485deaafbdfc6f9277ebff5bc7522ce627057e4ff1aa256e2a51138747ee1582075ffefdeb92998326ea411f55d57fc3ca203f04f008bf20bee475601eeaf343db0cb5ab2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143b1a42c513844f8bd76f13cb80ff359447152eeaffbe362bf3179b0d126174f3cb15fd18163686dfd1804c2db5135f4817e15b528def0667e415361c49ec17559888091fb62f2e91c15dbf3023f54b4867bb89d1387f73911658e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f3495b406cd93763de1c4393dcc1663e30698607acb800f6e1aaba4cb7dd1f33db7e45242ffff5143858533f8ccd2c77e2bb34aa1554287e6326128329501755a873b7170dd1ba601e3b6e0ee93c5183a38fca450102fc3dcf23c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2bdcceee03d13f9a9a5e1852fb4ead0f5be2c9b16ffa919d3d3fbab34bbd49fa333dd0754c6270812294efb545ecacb18e7e3bdd9efc16221f7a73820d874f7544c8be513e1dbd911d9846838a85f56134126324b79f91d2af3c2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9620b2e9680f3b3920c16ab52df01101edb92648f1ef360552c2c169488a82cecf50765343299caf985ef51f36606b1d916a46be4edc3a32251343d6000108516ae982ead976c6a966a9186d0612c24177dd384526042d06910070;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e74492a2aac5a55b97602b63ead8bb92be8912d28cab7db14595ca2a209e17feeb8417baf40c581221b25a30fb94b9b504c625568bbd15bca37e13cf167d90a1612f9a10b02f44140be2c1da1f6932d2f64d0b37d5d2fe4e8a990;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6bf296f4535365257896daffc271293f1ff83dff17152bf885068081076f3ff5f90a71c67777fa0d7cf824f36d78a2a0589a2f6ff30703054063d85ddfe00f7c1171a69b4bffd0f65d04ac427081bc97b9e00ad62e8b18a01e69d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h275a2545c5a37ac2b4ab509a71bea4ba64eb968b43bebe6cb8ebcd50dd3824d4301a01c97d4c64752da1e7ad97a004afdc4178016d747bbd2880e28b82de2f65c64126d4bb5d47c000f05353d5f5de3b9b6a503d4a96282f7e4d22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35fde1ac46b2cfc5d2f56596cfddfca4716c3e5c582751de34a99e16def6905e95ce872c1d5bf8af0cee3795ec76557eec3ffede2b6e3c7fdc9cdecb9f62205b3e4a273655b18006bc84ea168ecb67296ff9182a08b5f939dde4ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h162770d4832c4b7e09c53d05b2c62a3990fc40e4002d4fa0d5d69f38715c193d6d88d3de67182fcb751a03ad493646affe71127ce7687e72c935053207507d37a28f30b8c4c03dbfc4b673dfa0857fb6b005bdc93371e5dfbdc813;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c62553067f4234fcd28563b56b8da67e1a546720ca84ebe0bb06898cf040eaaf70692d7b6baada75d2e4df37e91a684fd6f9ad5069942b7f6e9283d2a8a4015351fbed407e1dfda874541e9e1c9fc0783e59073dd0d6758e1e3faf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a98fc2d784c2169ee042dc9f2824e3892226c07c97b4cd3a9fdc6d28d4859a4bf6c237ed78200d5086cd176ad67ef9e2e6ec463d90fabc5710c52df08bc4e263d61bb3a44b86ab2147b5455597eca74ff758b41dd64caac7f21f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1436d2b3dca057da5092767d20b4a18020cb412355b6f299df59dfdd6f90507ffb188c8c2756e3375e7d157a1b30f89d2b25dca8933c0ae1e9e01f03ca484cfe557375f710186188ad04902eb24c30f5f218ce4a2a33b3dbbc5c2f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137c38d681599277c8334b3ac4a40c1d6d02d3b242bf21f1acb95249b80952e60a25b244912aa572e65003b918389bf9990e2908bf961a25fec69a2188c17dfa3aece7c41c44057d2649e995d3392899cff97016f877c6467ca1652;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49af5c24e57360b579bc6bc2eaf7af1bc7565e65d5a0bb5e0a1e8ccff883e2e2c1b61aaeeaa2b61ea09cdbbc9e3cd3eb00b16cb6093b3c9fe2c756009f5f99d1300a8eb057b50e41dc20892eb715d15ad5269bbd359a2083f2c3f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4301f645677f54bc1b0f2d343878118409a1f0c4655473c7b2ca89d9610abbe5251fdc5c4e5dcc7e7c6d15e2d06802736f2b7709767ff7e25c1b46ae28cc34bc12dbf9a363970e2846fa3a88ffcb158362a02cbb772b2e417d8e50;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5762f7dfd3f2e218fceda5c5eba184cc9743815d8047eddc963198b86f00ac9535831d6760692c908f372107394cb41ba18733f72cb108f39434e40885c4bcf8387b75082b5ecc899a6d653d38c4ea8376a718f8e77de44d0628b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ede268ff1bdf92ba4b06f8794817a1daaa52bcfeec419bb822baa4004e72767e94c46de16d26d099ee0283559f224e4a9b0f9941296db7eb070424843817ca8b7ff757c45c752aa9f54755c51607d5b1942808ad312fcc45f81c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74fccf072a7e19e3afedf94ec24746eed95786fb732c65154918e246c6690fc41595107adcd654fb0d0994f03e46208e06457f2c124532454ebbd115bcdac5d809ca8deba54d06ac90a18dcc04a74adcf08b9a8c0332b1df9fd0d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62bdb963c95c0310346dafefe2d5f9d8ceeaaf3f2f2b5313c1fcb8cf5410a445d7cc4dc18a44e121a875e4423fc9a0bbd3d3b1d7e303b937100b0ee0720b6b868e7d23f66e7908c56948a07da2e552817bd990c0ff6f2c015f42f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc6b94b83b5e60f4cf9bc3a859d96132c93dfafe6e380bbd39d1e97174e85597442be903577d1ad584759af1b1cdde13664312ea6a0f22a5d5017f423ec4a2410715ab96160b145e72338dafac33eb8fd98e2749bf420ef3e167f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ed16f23f98b3fb45d15a9ca21f01b521a4ee10f9128492cacdfa97ef5ed034f806e60a055eb3a98a0e6314c07879a0ab96bbbb25875b14e47989b78aa5e4ff737006282cdd5b5487bae462a7a81937fb90f95da92c9257d6a6b87;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc9e4bfaed7b03eb8f0c6e4f867b5deca75c5a6a805f0ffd2e6e3b23a83efcaf99243fdcd89bc66ddfb662a2f7f73f87fb5ca7736eedacd3ab442be62df6323ba1bb6ee058c36af5e6ab05ef9217b1efb494454bb58af0f458f40a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127e44dd523c98777bf5223d5612d1261d1534fde8100ccafca2354a8ebdebf19824038c5ca954a3d7315479c4422368109077463e0438cdf802a8c124f0e60dfa7de424a6a8739e24f8849e36532525c7a535c72c4420ae8de93fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfeccb2a5d8c8294eb9a98827b13d0d3c151f94012de1f739f9d2ee7406ef1923e462a8767a747b8dca262c1e293988e0e299a836e689c7d648b023ae7a5b29a3a5d71aadf2ba6f7270e6c3a7deef1a744c1aeab334480b40d23f77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7504324f4724bef413bcb25eba5ee35590e792038e0a4b73edcf954b4904bf90dfa9fce849d95015b40c32732026eec654878265be5dfe1900795f9a21f34e068eafb1fa28875e0b055a93ef462852bfbc9ce80d6e4ab6d7108ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5227a80c806310d300e318417b8f8e7747a850ff683d1c78be3cf442657e361ceb2f8e4117eb787b5c17dee13bbab0c802ebfcd2d0929641a31b3755a6752b7aab4f099a3074dcd6d07713ff77542534acfc674c016491caf691a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6439b068faf4fee2153e76913fca72b786bee44e4f9b44fbc4cceb6443f9c2409fe44f3580a80d6862ec1679b13cd4cce463f8bf36fc73fb9bba0d685aafcb04930382907b39d660c0c12e5631e9565cfe99814305846169623077;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h719dc1fbaf3ea1228bcd9e9c251294da1243ec399194e4ec5d50ab10c40264c9bf13c43463d35aa22039c3264e4ea7335486a1070ca7581afd8629259be5e4555cbe5f1a0f35a06f0ffd741839f5083018176e2313739afd007a93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h730e832d4755a76a5dc08f398f84ad5e401eb2e0b7edefc126b77a4172de94ab988b8d8d128f648c5200f3b2cc0dc0059f97d6434014a994dd942f31a817f7a642719ebc7b9c6f9e705e6836f9264caeb542dea7e36ce24b69016e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1ba8c2bfbc9d4fdd41eaa54ffa485ed4ae2419ba404cde173c22e50096b31c9ffdd5714bce2090ed348c3662c4031ee7c54eb6f5cbc5c477bd637b07e1eb13953026b0f7a6b0e98f05840d29722a6fff79437b78b13b555ab54de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6fee6d69c0beb01971d97f9fa6d3acbb77d8c8cba69aad7cce55134ebb126684874883c83beec4ea6c446d08d907b68bc1136bb009cb42e6ef5dd2baade2948638b47dbb3d6822a28299089f63d682c1474e75abe85ee7a861e9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe1c8625e99100b7dc40f3de2e1f948e830e63fa112634bc49ec5d4e4ae0f9663cca4c9d8953339417b1a851e2793f3439837534ab4c3f5fd806ada4483004d1ffbec52889ec8cf8a0aec7c0fa767a1fb42a978f63fdda0fe03d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13654d95584a53549cdd5fe355cc771e0191821c9dee104211eab6289a74c0fd977f4f2a69536a62860759ba608398ec036d94f310c57fffb0a50b097a0bb6992e3e433a7bcff2fec4b8bc75d25e9c2f7802d3161a07d9ce5dd4517;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea3b3147c107596815ae2d8260e517e6ff24adf06f8d2a678ac254ce4f6593894eba9f8a38850f44d2052287ce8c868ec86c0bad9c974faa81112e45ae1f44749ed057791e905518a204343f556f5e288dd8ebab4dba908a9899e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16779a68457bfc24fc642d11f9fc25e79a5855d116b91e75e089ad78269b6745792344114ba236a5be16c838ab427e6786a0c5b73c235d2e301fa419804368e5dff93e89c95bc79a94b03b9f6ea0b6c6de2555038de001a3e843249;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb967d2362c90447664f418db245b177280486a062d7873c33b891e1204d917070994634d6c8cbe4d9731854d06735ff97e61b4058dbbd6e948b392dfad6026e40f405429dec616a7b7f22a1f88ca6c66d9deac8d89e84c5d52a0bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb7e7b0e4de531b4d076f17b4b20c5569eadcf7e105c5a912e969a85ccdc26744fea673c57999b40a844400cc0340b5998b9b64e85dcf965581f85aba8fb198ced028e92eef3648729807b7e2b79efb436b9e9c38e4478a7e69617;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbec63024914768f67a3417a4612a76f02dd6a24614f37d288724102cb12200105c14128a8aaf329cb7d0d679b05f185f9853f133397de58d75270a973084879f3baee7e133d49d1fdec6a79c6b0cbc183993325a5a1bd45e2ef41c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1568ad1652797bc288b75de66d8978ca5ab0ad86926b5524c7cd4b7b70dbf821ae8c7c803e1b61f997db1afe256b374f7410ca05b8e475b577d1cd34d098b3c4a680c7998e5672b8c7855e0e238b2311b5c89b7a2b6e68eccd456d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he20ecb1b076493de2a7f9822927d8efc09763adf0fc80619999d2c01bf90968dce4b8e223d877449f0ca04924ef5832e40d4d1d9b37170dda80b51db17e1612c3b2e92b5c16d8fde0b85f8e945683d3cd67bc4d33c0937f57e1afb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1315abf4a9a9d7f7a6b0990321bef278ea4a861d9aaa9f6e4b2a910efd94fdb23229c74146fb4d044d9019ec9d9432bc78fdbf42cdf4d4e0d10db4ba4b517f735ab6394270d7bdd561e2d82e51e11658c4c2317d34fc16e1a122958;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131fa06fe0b1a4128a17d26bc1d51271a2bd514e6213473f78b7d7711a2c60e83aeef07becd5268f595785f17ed72c0880cf2fbe9794be471296a61413797551ab9586689eb908546a866df84e8ffa93af5f8132849c153a00091af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193db8920367a66fae8fec81b7e8c5f359fa3162dcbb3cc253dd93751dbee95d65bb3683bdf248d732d025e7cd83f305cfce5b8fe4ea3df76e2cac551c5cbe2a5c87e8d6c450a95911348b13dac9f2128db04802aa57df21406a85f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h689b77a10bca3429e74f691e704bd552b197ce3bfc4769fae76896b468f1096df1194bc6594dedb688e7d9012296b70bc251dcc472702db7dab3932b091faa63d4b7d6e31889c9c59029e751a137ed0c11343f09f68b3024847989;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9739a9053254ec67852539987d580a4ffb17d1c8ecd1c28b982380fb5c18c455073ebb3abdbd912fc535eb5727bdde8e0fc065d9452da07b4fd7ac4c14b891f33d463df3d37c4380311dd22891e7ab0488837b3bc596dda5af45f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34829acd2fd8a8ea6819d50a85a657b9d54015eb29fe997f5643e0b9839fbbcd93a1ca36caddd37af0002bc05362e434d5d203521f34f8ff3030076b0325f622b06ceb5d14b1c2000b4ef46db1df7995ea4ff7002d6b6cd7c55a61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13201782b246067f51798be48a9ee7e9a2914fb3ecf5a81579f6975f063e370c4d07dd9999199b9c57d7af4a01c0f58241681032125847be6daf97bd7cafbd1679a2bcb0f9e5c2c564eb694d22b92a59aa592851dabe96b2310bc5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1414ee74e4db0aa53ce9c7d6b01661e38ba508e06f2ff4d0a027afa0e5abab13f3dfba97fcdef71b135161b8d56275a97653542e32e81bf6dbab52599c8426d8d537b83c9c86d932730c6ab7734f477b4cba0505504c9a2476f77e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cd451c9433089245b7a5a6fa9d9e461c8258094d9d3d522f195c0fc0bdd3f867ec2b7c23059e7256046062e76192ba9d13285855e5482a3cf52c7b8694f85c7901e1b7d21fb73e0db94477cedf47651a1d3b0628504e3e5fbff69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dda235394938bf52e519dcf8162596b700675e84aa6f712ffcc5265e0c8253701029abc2b1530cb72586ef4daf140f6370850e75672d8441ea4feeed18e353c3ed18a01a5d9fb5c38e57cf6bfccc8296ef43cae60fb6369f45deff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2c42cd8c032d501bffe82d4a65d074f405fa21c2eba65b88aae3078056c84e782c16a958dda289267c510e7b33db6f7f4082eef745805a6b677ff61dd352fa404f026d6b79601fddce3f5f408d020138af7d7045da9db7a43c226;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100d46f0634a61379aa117e14b138c991fa74c5a8a401b997b2a8580d064fe983ae4385ff9b1e69f89d5d7ed5d0a2c66b257d432e87e01aab7cd4fbb945c606cedbf22866613f494632a924f45f0f719bdeb47b381a0c8a73d70331;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123c9d214ffa2019452b892ddc09b12f345b8eb4b5fcde91e78c2d1309e1f9cbceb6bf5365946a680d9a97fc8a47bb3f8312511407ce9ff40bd3a1be3f582a210d795f48d356a402f3b46952f0f23111ed80a49edfc7a7afde6f674;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h654561857bdbfd93fa54e8de85ceeacaf4112cc7ee44c1b7b6757bdfef061883344947898ac89f725b46fe67cb9495c7c8c580dc381f8deecc1b693c3fa41f49285c841aca2507048fba88d432265db090dd284767da4270c41bd6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5e1857f71471a03cd91fa3b8211fd5b9dbe41051af731f4b6838282bfa699aa5b422cff82db73185aa1933c4065ba837e2b7b629735f22633be3d9a0d263f2fb6e86c2e464b0ea7f89a9040a2a79f7e9c9ec240048cdc0cd5cf4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65fd7692e9381885192474feb652fd137a4e6bfc0898727ef1f48cb50f5ec5ba1fa858b2fd48023a962631593213ea60ba4398d7f52d383b493ee390d35433abbf9a87e5eb26314b2180269f386acdee2fa562d92d7fb76866fe27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f84c365b0100a3976327820ab8c07e902aba4f7b8b86bc022ab4b7ca0516878f70377f620f7d86833a21bde6fe098e72e2acaea299bd605769f452bf1f463aaac5819d0c3c9451de664d9e47407bd40becd53e9fa9f2fd4ca803b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b51e0cc14507c336b0f029ce823ea0bb38a8d5b4728bcddd0635c30515371ea1b8e6faf66fd8d471926df7a6c0e81ce8bab175ab7058d3537f968e6891c153b40ac185fac08039b3fa589ab4e93a4a427ffa42dc1f16e879b2ee2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1588b75884b3b290894363afa71511f17bbb9d0a8679c4624ca9135325b93153248542035402100ceb07a351484b00346bac8ba8b2a37de7144ddc3c0256b1136d37e137e6cc565d7789174dbf140787036d3128a7d451c2427fc38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f5ed7208082f1af5e56d872458db53e3dda87d48844a5693159782f98d6933cbc1daca1a0ce29f6a9f05bad8854d6bbc0b7ad476ebcc41998f8833af41bcd732062bd84970070f13d6196629e5e9e89dc096024b7d6d5f86f7280;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2626d7b121c3edd2508b3c37ea76675421f53e880062e7a338b57cc49c03980014bca3850c76e32f8ff09e848cb88782e515eb99bc05836732ff36533affd7f37a015f9c7e1af69983f1089ad368fc1489a231c3a280cd42ac2125;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e23bec1a741df741ebc970771cc2f59e324d020817692402e7718e565e9c25eb6c7658839095eaa0985d295c893920d587442b90d45db72b3574a42a0ef622c61dc55948856b51168fce36b9253d5ccaab9359d47dbcb93b9a1c9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef7bebd701adde212b7c5f033130bdfcfdca82db6236df084eee34c72186bc5d4a7f29b2eec07fd3be26e43dd8f865a14d53b3681b33a09722d5f602d63aaac021bf55dc5b3f15a1f4b9316ce282ae325979d8569831cad981008a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe4689ab38b3c0a7915e7d4ca1962e68f26701d396da3724cffa4fdaca671fe63f24e267a11fcde9012fb83564e9886d5bd91302807be3b732fd008c1d6f1a30d105a44b8189b207b689cc3f12a9a246bcd3e6139dace3e0b969;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b56a3c48bd4ad46c521023eb0112c24ba8ec9f0e333da139d4418142e997bf684076d607e913d1e8dda9f2f54f7936bd75d4c4bf75252152c9f821acba8cce12fb06be8e9b6d4f3c14e0acb66e0a961fd74b7357ec8af5848c493c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha719bcedf248a082ea6c7c78d65937ba212685ed40a7474c0faadf62089b94c8d638b901db310c8a5143e847c78ccbd356cc883a82460941f573966616ad093f8fa40c2c4cd593cb05955f57eaa0e6ed4a92adcaee0d4dfef5cfae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75cd3a06f5a8207d1ffe68f805a8f690feb27b77fe8f1e555ad23f19980e2401d80c51c5653b0152a7f0017fa3826c240dba912bf1c46db0a57a7e96030953b38e4ee5b81c05e0f61e0966d664213f5c564e85955d6fdb8b7e7643;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdae68be1dc656fb7002bfae0bd32785dbc92fb10a8997d7277c29b3c18d1d4c4d2f8f931aba60a627bf8fdfe31b5da5adee49f68ca609e1a5ca26a1cc604788f714a228b21d6391a769d889d8eb4ee8f38301d74374f45e3a040b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae5b3bb7d4b92350610ae3653de407789620b9c6db7ebd96892411a984e9b3196432dc13d5f42ddfbdce71023dfb23d23e530282fe4e731985889268392b18bc137755a9cf3ee9d44d344df7ccd64d835972733e9872216d258e28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e2915a070846ba6a6ddd6d65057e1ee90cddef844053c0b325a43ab6f79de9c546baf2aa7f794c6397a93606977baea832f51de7d779b9b53e50e113cedba7e9bd9936427088065131deed6888109087c8c50770b4c3a420d2a27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d737f4cfe9aa746a5fda86f6a20302fde7f6a0a62ba791059aae4bb98dce0fb0b85a1bc0ef75592641dd153c5ca238e598f434b685c110649cd5632b2dfbd5703b75780d4ffafc4fad136c73c3b69c856570ea64553a8da3c7cda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10eab21c8041b5d06033e6569aecdf76b8f85067235378142ab251046f56a780b619261078768ff1136050a563054d1cb20955403847e5cc1f759082eb58ec9e37d95ee9f3da9c92848fef2bf13bb885e6aa52602fb08c495f50dda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11371d4f2b6a8ddaad37fc64bb4c35f8e95e9d1f24cd7fe6a46a16b91358784ff768327df921c31466206cb5892a0b21957774a71d3ee7e53b058bdde100b379e095ce3916ccbaab78fc63738973b0e5d4c3d7f02ff94009402c350;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167eea2f0e4ba671458f0da165523256aa8fb74be5b1facda5c8c38da010092042c58a33a2209b9f6fd0eb7b2c1cb3164e9e51eb96972cbdcc0857376068e890f5cd2c2d448d4c059b2e0279469a35eed519589221ea09937e9262b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174ce43f5cdac75112586eb8172b36cd286d0fcf03380a8021a446456ef9d90cf323e476b08d82a5cfb13e4cfbfeff93e0a9033d57812d32109670e1fdb4ee5223ee9c611f912c9bda91c713bb7f7313f8146d86c8c09e94c2971af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b160cf6a6097b8dc5b32a1254a4854e534dc3656848d03e5872999bc4ac10db6c710a4244561b4a6759baf9f833b0f190c458d59cb545c01c65c14052de90b040073eadf8713468bca5f60b3d4a350c01ed089b80bbfea5de440e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd397224a1d8c0653e572e829a1adab8659fd5567002f1e3fae64c02f0e75382d4a7d390928deccc3e51e2d32ceaefca4d0fcc86e4aa11383864d715c37261a7b24f1c64865c4e1ee90d361bd471d0f25e6350e3bae372f8956486;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hebf83879cc3b2f39ec18d4a49caea05cae2cb8b7e429af8a3d853499d370b4d5d86b7453c86705439d610b712a1b179be1d12207553108a1efb13a0f1b52b23501859e0ea61c9b5876de59940ce06b085a0fd391280cc118800051;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3561bc853a3f182aea842ddd9cede5a3261557bbb27f95d4f31581c523ea482ceed8a1ba4b177583ae1f055a125323738f0b4ad56f8c070c09ecea21e4e36f109b952ab977a8cbce7a06126116d416677a2ae64023398d9c60aadd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc0bebab42bac511d70ecdd7db3631b2c0a642ec3478476a5a733cab325fbde97f89e64e58f8b6852ac1618dd4cdf69080ad6a3a835d9a0da1effd6cf01df779df3bcacb427e4f3fc1db62012cb00d06e31841d3fa8ea9cd015596;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec852c7815411ac2e5d0ce3527df520afe3634917dfa51a8c9cc598cfe00befc05080546eb804c5d62272d1b774fa20339e6a2cca6d16a79506d63bed61d6a31f5709ce5ff724aa550871df703ca2a655ce97772a1cbc46424fc20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15347b96d18719cb18a8e518cb352499f2802f3efe1cc0af97c028c5dd93f353b8021cc07d44c32d34f3c2c568cb6f6db09be3da5ecebf094ccfb50e229965cc0f50d9a93c5435114ecce66c888019bb3f30b3587c0e6019f5340f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125df7cc897e5c39ca91a34dd404951cb6cda0110635739cfb935c7402ce39f8000ae13fffa14b2ed7d417e5e2f28c6cce395b53303f451a9e0a3e2207d49322b7fac4333fa8d6a16c1a9730653c5644cc9b4bb8ee1c2236d98cde6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e737c2b91b34b016156e13a0015c0e7e2b1facaf79c784d1e7f44ab4665f201250cf90042a3c4a405b23d8dd124aba4a4f19ab3c84077a8f8fe256be1adc1946503fe6fbe6876cdeebd8add5da03ad93f4dac595dd0768a40ce094;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26c67f1ad5efd72187b4f97b1fdcbe99f08ef0dddb6db418f006aca0e00044b3a7e628cbb7de5d6699de351487caa878f9042c7367daefa0bb7c87f8689c2a91dea5a643040ff2f44e7c6c4662f51f9c07d5a9543196b062ca3b8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27285736bd4242e26957f564dc72003f55ff86851cff6403012d879bd0710e50c21ba9d1e0d2cfaf0b0758ab79eb8a7af1eaff8b8f2c8209357e63842b142682ef11498d230e5f7bec9fa76ccf9ae0113b7a32de967afdf1115066;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42ba7b5ae03ecfa490a6a278096364d90a02482e7671cf65ff0726796f72bbe1cf35714d31c10060f4daba8fd1940e4ac1049f18e5cd01aa6a98339edab4591adcf9325cf1f94487edbf5cb4696fa20261b5fe69b415422d1d83e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10aed5e787a0d3bf3024fa034409f17d4692a3ab9bb70eade2e3b44554462fc7c8eee6989d292e487c610977de12fa853d134875113dda9feb353eb6453750e1c2cd553d906261ce1c6f030f7d4c40bc958068d8f31ebee44c62256;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef38ebab0d36b56a803e79d1af606d1e237b8397ac293e0904c10f487d02d20ea0798c424b765ea8ecea3dcc6fe348f800b345e1119383ea601c76345bf8b00a82a2936d78b34f1876409c6e4effcf216edefd112eb8c848857b0b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93bbd9f4bfe7bab8297c439caaf7628771c020a001bdafdc8b95430bc7f48cf69ca6bd0711cb66d7b1e0b57ea47ddbc2d69e20e9e4cdf35a36e951d84d4228f6da88d4af984fa2e7ea329d420df41cbec0110e72e6fcd28496628c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb859f8dc88c5225b9faae3f5c7e10078b0a3d940c333215e2b91279aea34a7a03a7e018317469c99a7f907782d7ec2f7afb8ba7f3ad1d97404df42229116dfb6c975284a31414e88c7422fb3a129ffbdd6f1eea3af8eddb4959f9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4cec024a680eed7c1105ba840caf141cf902626735f6f0938fa357946623fa69d41698cb630a8cfc4b2daafc0a3a609e0d7207fb726777251086dc8ff95ae00902641f561c898d5623da1124ed9cd270e9cc6d5de7e84f04f3e26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0dacca35f93b2557c46cf5b8a5b1c4f0e197d841d4e7c6bb222675d6b65bf913c66670f90b296f33af00ae96868aae9ddeddeb09d3554300df22df79d3382fd04917337c89bb88a403269323056d27aac3f939c8b67e5dc839095;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c09119680b8bd2226944fdd161727e27d3b5962dfec92fc4f9c5e040daa9a8379e4eb95e9e0b1e0a543108d6babd9ad859231b4d4e2a5a7ba8adc78d0b6239b2d66a1a6dee985f9f3d7858a77c0d77415a96f7714c939e171287b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b03bf57e1f790aab0e545c03b76661147a41fb0cbff185d53921a86fe8f15dd4fa8a601792a604aa54e94bf56ab3ba24d0e245ff1e2882547131aac75bb70d9fb620d9b9123728fe87222ca7ad752342e1953f870f51a55665226;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186724fe271adbd5f49b1aa97180f7634a5e1c26801f3a08cc5eee1b62bd6b4096b3a8593fc776036967981c5c16cf4080a08211e0a177b0a7e2f7bdc793595d9a89c92dd22ed9526388282c9ace14c5b0585e885a7fa4df4794b66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h585f1eafe27b117b58357ddaf62a9c2d139f95e456ccd0a32ff20892c3a6cc3d6148dba2a285a0047e5102c08f07c5f20840ea42b3fecc534262455a87c836616193eff65d99736a6a72efbaf5940e3d35372664137326dfd51930;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dff172bcc955a3857ba2ba79fb5fcd32537c040234d7d44a8985dec0ae8feeb839640f755929ebcdc6aba29810f084997dc376922b31a825a8fdaa073acbf48c98887850d3bc26749cb61b3d6d13df016d598cb250fa6d047efe49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72ec6ffb53fe933f6eb469ffe4e3322cdd94f0e78675b0f89119a04a2c105e943567014bcdefc217b98a9cbdaf0e35f70922e698765992d667f461de4a139cd92a6fe915782248f467d4aaf6cfd1a16e75f966918cb41cae1b982d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd54f6fff6c6c557960e2aaf7bbbfa90adbe1b657aa40af1a6845316b035da0e4fc8d03f6cb70195562b98e29f9e30a5dd827b95092a6cb90495adf54ed89a1faf6378c7817634f4b2bfc109996074bee85659a4b62af15bc95cc82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h552f05f3294c4beeb2f540f0f091275b3e75e0db862d05c1f4523b28a11b2727ea3a3a5955ce56f059ad65e4162d0be864e796944337f42231818c758296437684456d3613dd0288d95251c47a5f19464591ef8705e5f5aec5c476;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5941b35c13c415ce0de5f41750a41c59add04b6ac7dc666be57cf8f8124412a7db5dd5cc1dc484adcc0c501f9ea3c0529c9c8dd222e0e4e4a27c27e1917d8a4f1bbbcde038848fd461a168b86103fc55296c839fdf689fcf0866f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12563e13c6047d23c2347edb570e12742aa62e869cdeb769ddf4e4bfe9f789ea77a72b34bd3bfc7893b1391803ea7a030a23d699f028072e14a81afe14cc13be54ee94d6f427754fae44b45f7ea30e78467901ce974e38a62bc67b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68986295d37d2cfe900be4f944beffa6b584affb1b401c615405156e5fe36a95ff26afea583ddf7fe000ea2ad5784637aa064db9c8560e397dbd0ed1a0ea920ff682a9ca0d3d5e7170bcf1639a81e27133ac44bfb625979500cb82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31d0ed7e09a1b8dd400f968f616fa225819b67d354b8a114493116a56ec1c2aceb4a85dde341d36f77355885ec0e07cc3019e73881ecb0d0a57ee36c818f6f44657e50a5788bfd47d814850f1cb1a8e5effdec4660f9153c4d4912;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30479f6c8220dc3fc8229c5a9a918f04324bba97f3ea779d2787a140dfe2c12fac6878a35263419195ac42c76d2ab087103f8e692211c82f3a74de4c6053307137ff26eca57d8e804ca8fa265a2900f154bd1b9ddf9bc033c970a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e06e4135f7dbdbcc462337bd54263e9aafaa1ba5a288c2d51b99b79d2b6f51a8ffb15655622032702a54b7814b8e1cf47ccb8e5d97cf0462aa2d44bc21fe97f9c5ddb3ad0abe42dab63cea7ae4d48aa140bbc8adb08d5d1999e86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80a6caa4e18cb68a6d6504a46dc1d89594d8b9f2c53cb65159495daaf6300a687ede891e9366066cd155af1f4a4b9d582f46c6079e20d441f64c6b853d07d42595794c8c23c81330b86513dd6c9e91cc412929f85c6941022553cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e52f227aed70dd77c9c3ac8a5ae84268710a650edee022c137542703588082178adf711c3c255d4e62c8ecda9058215e07653f2d2a86a280bf3a163739cde620bac28e1b04f61eeac15c8112172d860377013686cc7ced5cfcd88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb287dbb89c7f226178de437c6c1b3aed77d55ce1ee267e2d76a8481e68a99d3a6be8ad1806d0bfa1e8bd56323fa17cbdb9d092db4cc2fc4aa6c5614586b2b0475667eb27398c6664e029cc0d3924078fe1212ccdf9929d8a34ed6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea27777763c2f1bd697b6991469b60dd3dcddeb0f3b8be95cc5edd12ef827733bd30ce5e1ccc3b5e58e504c3a27c3a3da3c4ad68587a62486b7b58f6220df7c1bbbcf626e22a5219db12944974d20a55a2b4a11f5b68a87a19f639;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164c7a120e46a5b4a1fcc2e1a83cd2b7e8820a6c8fed5a1b9f5e05137595582480f97473c2bc6321d06e41229d5853016b85654e90167bd182d3616ce6dfef01d011e2a109eb49f1b5115e1e6df5f88f8aec5041fd925092fe9c522;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29780b2cee653561ba70d6a6cc7930561bee37810d272c1240d8a76a12cc7538f407a37a585a1e4bce11f3ad6821862f75df74d724746f508cd22622cee2917aa0f56c37cbe6e4ab204db8e8d4503b38a5f51e953772f1933a5977;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h789d61ce8f6159843930c4fe16595e82e2f6957cfbfc1c0b8ecbf51d262a139f9c15f62e810e4c914f60f8f5f0b1eee2c0b7ad48866f17c9e37891c9c996c07a122577dd820827c9e3946c0a0a164267c31a4968893d394bf3fdd9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe181b2fcd5ddd7f946b12ab081da774f5da864b3b0f3873729dbd2461a54e4bc3545c19e13b64befe1b6c95be0149344d44840a142b7d6e8363354e3e3cfaf4b204d4aab4876ebb4f7429fbf5eab6c7f99e7d7b5fc33ffde7fd4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1679a7f8768b96ed48d1c8d18fe875816e727915e173c83ae79b1f1deb8722340941f415c70e121eac9f23caff95945244e7ff830d36104a27aa84531c9ffa78a776e99b92cc83e5cfb11bf7cc9013dc82dd81110d1b8137bdae1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h735a485d6ddc87a9e908c19791bc6a499685f512ee7696a565f865309b9887f275f6dde296ee852a4461c9753efec16e725eaa5c5230a027a5bbf3fbe0285a5c7b1146a57959dc1f4c5433f245ee7e065545c13994f1aecce601b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180bac92abec1ad5f1529c00a4b573774551e73ab12c07c24802e680e9213a86a228800b8b57e15910b2631a84e96f20c60ce7e3dae66322de3f6d13cce175a0a516ab0e1cd3a9d269b6f6c41716c4723601cf1e48e5fa74cb7b444;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a0c3cd6727b508a5c8efa13bcc0910430b1e351c3c75a1ea1f2b0ec8c4fe8bf10bd803f24638b69a1b07891bbf403cf0a10d6cfc831ac7dd921af676ce7abbe6461b159d437be48e78b1f25db3103b1ec5a64cc41a4e7257cfdfe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h836aa0d3528e5145305d74fe110a201cd3f51c2335e3b6f2446ec0cfe18371f486fef4dac196bc16fcea026e5b02272f26b967191f24d5eda655519878b2bfcb559bdb287dcd04f24cdd814095b0f0c22c4630af86c4c1bb616208;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f6252e2cc20f448609b654ea7ca9a9c4fe19af2d60545f9122c7b64ae22f864bf69d6bc7cb8c8afa209c359f0e118aec19f2c8d8fda5036ad1d57c2d9af7d6c0b6d78f4fde67255977a545267e458f73d72bb40285f8edda196d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd870711574340078becbfee9473ecb5139cab997bc66b2ef308290c18370939b92ef74eff6853e04dedf92e2173d354019bd923aa43496f9065e591b417ee953d306d0378d7c5deeb7505fcd91b9e6c3f21892f2861aa3da18d9df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127816ef652d000397ed193e396c47544c21d82af60837a8e3b3192d6560ee599c254008cd50c52926ef1cb17f4e6dd001c01e93a2cd8cb2ce5dad7b062fca18f34e1517a892f239062986dada34e4e2288e2b9b1132c11c05d658e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he624f9ce07e84b221c830fb5988f099614ab50b7f5d3b80b356ff8f64bf95f1e2eaab29906d1599d9b2be892d3c857798c1ebfb23f733501a3f3ee1cdb03a1ec03ad8bcb9c169c24ec06ab3aaa6b47ef49474ae46581f9fbda32cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6219716a2b738d698cb23d899712f72d8028e4e120979949cbef322a85057078c9f18cd5a72f017054d18965e38e90526f5d4910dd992d99eb20ef6e3829c6f12de336e91dad34230bdb51d3591cc628fd3a8ccb869d7c5435a908;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h946ab703d8bba825365a2750139b6bb59b4684fe226097b81ae5940f0d12f206f7e24600942c72c67b62874e7081c66a725deb267a1278c01656f387d67573a0d796fcc0667d89ebf9001c41f70d5dae12b23d21fb3a55e1c7a68f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b87cf0477bd9980b7a7e47974980cd12d6586c20181cdf502b3c19b36630c61c6b68a8a7fc886f607a9e1955611081031e120bffec5387bc5e7f46313f70fba27db09fe85d53d3b377ff632cd41d44e62661806cb64a1cd3f22585;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2bc82f4bf9d5202b2de06dc17f42f24668c4ee0ad0d2887d136ef3b56f5cc92a547aadbf53af526a0cf0613b3d352b2a6627f36a6bc4273483b85ef2ab0eedd33df288193deb773790a71e72a8850312b929e4484df8d4b1a8ef8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf9c4d6645cb9c0a35ca345b7d284d1c01a2caf8f5a010931c432f46018152263cf8cf5d8418951474468c4f3f12028be20e05a9c09ad399cf99328bfcb7b93ef5d19e4b6f6a246e51954a397587b5e7da1baba028b683fc3eecc6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb56de60413c9e0158211bbe81b81044aacf812b6c0a0e951981bedb153c84178fadaa351324245c42007b3a7c919bfd326b49665cedd0b648354dbeb5e54e79c4ff7945254d0abace4673ce359db6123c7fc8977b855ad4c6d525;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9af38df1646f506e2127a05148080e17ba97421e274ebf6383f13c7758549eb2f6d96b3e144e3aa0b510826ef62f108df94f444c17166803c0eb947bf27a242050f75639f5505f52f63ed3bbb82a1123c9ef836d4ebd49cd2028c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e2c90ecf83fcede33a4084589124fdd6b1df9ed449a09518198ff23c68f69ddeef01a1f6ebcab07ce311193988bb4ffcc930f0b3e2e6e6bd8300ceef8ca9b3ae7c50fcb827bf16e900bb8f25c24e15361fd169991d6a0fa7f5328;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e05f1f8eb1f3bdf6bdf6c0b76d9e40ab5791dc175fe83fc6b7b36b2b7dffd271389bc4cc975377ed151a57e08316998cbfb529b98a78c78bb8821949b08acb9661cb95696e25797b161db2bf873d8551e747823207cafae1d9ed28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68960aeaddbca8a980ee29cf1ba23d926bebff1c52c2e00ea3099092d785304c94b796c197971533dc39bb0dd892b6cc56d2b464d7cdfd13fe90353bb0a55cc30561226a8860c9a6968b7e2d133fbef76602079893a61e8c7be9bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc02b571b190611567c29e140b2d59fc5bc0a635deddc2bbdf093c109a8bb527c9f0c6808b4a2086611a15e3da56d38e39ef66cbb0ef86104ce068cdde5a230899437a16a42934d7cc3329f50bf8da6f9f878ba5a474c7572740697;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c88e389ea6fd6cf56eec04c9426f75fcc278778c607325a2e545991c8fd14233b25b7dde1a7275b0f81ab2d8a240d427e5c1d187bd9bd1f691d70895b69f6d0ea81dabc83a85b2d819a388d3bd55517071bb8d56ad8445177854;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ebc17291640029d3704def2d9d8510fd2583d433e60cfe2c77a50376231775516f01521656f15b501301d9665aff0503b4291478578356f39f8827bb559784e74ec24083d471b85143013dc4c88d7a059ec290b7fec11573dbfab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1241f35815b865176505e114db36d8d80d41ce68dd9492efd04c701e1c89ef58a92f7009aa62bbe262a7dd6398045a3a767103324323f7002e48f74bca36eae6e6f7ed46c80b4f857dfd31e29b7cd46ea523939ac371178e35c26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7033fe7a2da3facb43853bcbbc2dda8efe16b5110659b4d19a3b73f21191d6cf9fff93de721b1436c8ebd9909340e9a6a699a85674d86022aaa788de983f49afe38fd8a0537e615c807fc9b4cc3b09691a76e89ba3adc4b600479;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce329a3ec65cda7bdb55401c85bf6b24a304a70ed636c31d489bf4fa14580c9e45cc499fa1affb0a21ba83354031cad4940ebdc6f9f228e822c304b574e1db498143f2bbde00fba6226af6dbd5bb1808a57e76add8d5a7cea4dca1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c0d7ae1d5bf1b0aae5e1b0a1c389c3fe35b64e17066ab36b8a071cd094d1321c30dd31d003769da048688c6034733ffa050f74c12b61c853dc3ab050181522460a02b9ad77603e049bebdbc2fbd117980cf012e4206df29e6dfb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fb1d37f6df8815dee8a12f537f26123ea17a51f854d13373e3891d1b5def9e3482238d6d1e889d12ac1a4310b2356f7c023f93577aa908867d18c51e2a69b1db339a321495b5d47ed4354fcae218d2798d3452dba38aa225bc0b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h693bdeeafeddee5579d9c40d030c785a4eb8e483871a7ebc0ea5a69c7a5c6fac5f36c0e29137ede2e684a1839fb9a57e7becf8900595ff7c1cefa8c4f39d878c5758beb46cbaac3a60da016d47c9520a6374072c4bb224587612f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h286ade898d72daac124c114dec7b2e815d89c434f8497ecdf9085773e1e014733dac9325696d93c0e0c7d5046202f526afd71c65baf7dbe139799c38254940999edf258187435bd78d548ca22b2a01aa6b1d5b64153d6842055aa3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c2b075141a5f7e2a619631fd0211f0335b966dbe4be7f5fc0a4c6f5704c24c8034d74ba7e72f1565dcf9a9a118924c963f23e9287f88e118c89d3182f7712776674f1c6dc203cb3b668c6cf27397a4b91319d34fc3361f667787d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8f972748f8d72cb63aafcd216c83e7493604ead7f11815a95d3f6fa1a8f2c9281e5be9027455e3e7f1274cece52acff2d6baa056c51573c860ff52e2ae53582876bd8cb1df1882b918e04a077ac1218822ae35d64a9041939db1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc005cb76878539623daf93d5804f6719c96e2cda4bc84414f85910233f1cb91d27414ab055be31ec9383a6280aaa39caeaa30665be899cdb05ef962c44ae6873ab0e55864e2342c829b2efc8a592f9609f9668c9bd099bead67f1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1231dd62326e6fcd8ba1cef673e307c2fce60e1637caa3d669851b1e3457da6b76c18ab12cf26ede69a03c95a3b3f8857e91ab369cf5ab0191f4b5c328629318c0974dfb3422a646525ff830dc254c5ff8bca0c3e03fef4ef6b1d99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb19cba8a7baa8f068d6e93fa6db8b63edc68cbc29e25bf1f9916461a4b0af9f4737acc6f667b3a26622931f229817810d810836db4392dedf7314d2624f7010d1a055b1e718bc7818d0ee666976ca968dbd7b863acb6b95a632a6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6575e6edfc3b70eb8fa9be6be56be596b1bb556ef668ea50b9935ce3ed6172148f44d2798213b0714569ae7e634655f43d2f2c6419e8965b10f3cf6d3cc215e20413b3f5b2dcf94080138f5b0d7cd3c4da5c5c244ea1a9b12b1c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36b2f17f9969fc26e124d1995b0464cb60994715a9e69e270f40bf2655fea9879f0219c623c781ae518b6ebe6d714704f58802f0e915d919191a74217350a31a4427ca951d8375bcc9abe265783a22c8d467034bfb23949b38f825;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fa036d7fc9a3674df1327809a7ed6cdc7ff75d516e9aa2d18a96435fcffadbe078bb07061e1ab9d3e7b3cfa6a25e011081ff0dab1129f423c81a11c23569c44eb049bc36443b98af173254f22942c5cba3971c2f6991ba44d9473;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b6ea4d06f0ec20bfdcdfcdab3fa718a2eabbf4290b311d80e662e72c7432a609dd90231427cf519111a004114749bf71e990ee9bef33229bec176fee02685cfed273934289b59dd89c4c19c001d19b72b3dde427fdb222e0b8869;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54dab548188bdbaaef9b0825fe3156a60b7a2f67a97e60c7b070020bbfc29c1aa7b90201c59bf458b934b07f967acee723f1e5dc0678c802305305ea30e8672056ab365c0d21998d3e698fce1da0eedb4acb4f838dde816eaeca09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc32c34c8e77c2367f976bda46098d01c5f1b2fc90d555c7c0c46f8bcbd50eda93a0fc8208e207220998a3ef40c62b331534d708eb18534325b1eab0987e1794bdc9d2909771e7c9a5cf3aecb0344aaa454dd55e146c05a5d86ba7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc63c33080f7da263ead1ab782f25d286705833c55db42f480c53ab70c8352b88b353cec0e52582f46b9d87f3a28e554d69f3d2dddaaf8c2bb3fc86cb86ac8851432fbddac76a12e65cadbad18683ee9799b8692a82c81e46cd43b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16da15e175123231bc9eab58600391da30a704d0dd4033348f71de7f4e75923b3335249f5a2c3569b60ca51020f78ffbb1d9f9a50b53f362fb71252daba63cfed8aab37cfd23cadd07bde402967a3d5189feb4f1db9b0a9e50b9538;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4e33c0d4e192d5bcdc9b2a99feeb899de1f6ec35170cd3e4dc6579b375febd29eb7f09e6c36bdefc79865c2aea33b55bc1dd481a4c533eaaf40485bcdfc161253b6525d197c5e9ebabbff9229c95892a2cd5c38924cc798b2cbf9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4926b3468738981ba1cb5071942c05ff9c34343eeddd8fa912eac752ff231bb00036ae661acd1712fd40ed025247a6403ab41b09ac5a4782ad4bceec543ecea9ce188e416b6813fa875184fa17156e360cff1c5af9f9fe1cd63010;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94e2e3b447ea5738611b35a687e6d48f43e56ef176bb9441aaa39deb179300fe2ca8f90770c6041f5469a42b0919bfabe3112569b94d03284b971a3c92064604bb024b60d248403bcb7bfe945db408e88a24dddb532cdbdc173a2c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d801f1112491c8a288d86de3a3269d8241655e0a6f1870ef2e692ae3f9b989e312c476f083835d076e0212a5a662bdd055b3445897161be062c1b708797c5cd93f7ceb96ec97d546d8b23512cf68431dc86d72415131440df7157c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec262a31f11b40f8efe3f251f6fd94dad57f66a65d5cfa43ad480423940aea243a826314991e0007cf1299e4babbcdb744dc2cd3ba619ccfe9d78f79b4c52ee368457d5834cbbcb58cc3a6170f81fef50a98394d9b2689c230820e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c9e1fee9a9a84acaf349bb4e5113c1c13701bbf0c6d53f8ff422e2077c79cff7957ab59ef7c020f6d9f8d7bb91150879b9288378cffa51fe7fb1e3e8c514d7a6d6c9a3a07bc1b1f4c1d8075c63d63890af126f4c9cecde17bf24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6254606023de88538f0b44b04a623c296cd83d73c137a0e646f624513fecc83f9b8a1316a1e7ffff04a7cf970351cc76be487a105d8842cd4f6e62ac504044930fb71c0bb6207314c84823b6e94b82fa6ea95d51defc1dbe39b4f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b4fd04c45ad961efd01d70ef3d8e7bec44ca593d552d62e57e0275437821ecd18cbc209d8193a0ff58cf419e47fc858c9e9cf8cf31d53b8b7b2b71b5549e79c2ebdea2d93e69440d24aa84cc9331c7eba8eabf125dcd73bcc16c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e1614790721a69f83f3a14c83a6ca7e5d0b4263c0d4ae9b3651a24b39ac9fe963ca966e8dfa0b15d298c01e4d78c111f9a315d69f2b2d285b84647cd490dc9d70dcc8091589aa9e0eb56dd91eb0109697a7b8b6ceb115d2c3056c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f19d478bd3725b97be9cbee08cfa78efb1e4e886f03ce861117af4f9aa1bc80ed59be116807fada8c59c4d54e08411f87a1ae489d0810aa49349e0940a962538857ccbd42fb47a0c20ef5a30ca55e37b71853cec9ab593431f7a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h889c626852fec53c9164880fe7d5b9ab48bfccea411a0ab68d1ba8e7996dee802dc56a6498abd941fa34be7836d402f13904771a9be44e3cca5ab364885ccfca77537418a387675a6a43046b5143eecb7ab3c978ca1e159baf5b4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe8d3ccbd27a17a6090a99770bf7bc041b9a345f4f1d6c6809c38fa7b9e9c596c0d04bbcebf37679ca370a3a94bca2a2cc8ad160546535c276452961f2cb3f4f30d81643a92c65fefbad95135a25f183e2c9daf59db9bda61559a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13270eeda467827aa3ebf578361d2c4237c94c013ed677a8837b16d4fa21041f585fffe5f0ebb8c3115dd9fcd83c8c9150d688fd091857c273b5aa918ec5ae8b846aaff53484153caa840f17a09e5f794445b3d14eed7a2854a73ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137fe8eaaa854d2d1264f887e9c50d3bf751faaa8cf9addd7c912b32a7c84d02a723086069f6883342870dd2ab89cd60116001cb0f418d5f14bddf3aea57cf01117abb806a803b15311820eb176f65a57b983fd4329cb712262c8cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd65e68afdbdab2420b896a99f1b19bd6ba285df803a089d2a4906cad3e2d9648ea4b396d4a47d13cc915bf4c8e310b5f9a948f4a26abbe301662429bded7265febc29f1b39cac3d70d4f4e6516a99b437318477378d48468b10ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he82f21db7b5fb38ecb28d3b162c8cea7074060b2a4cb669025310e481bbbac101991192a45c43b88bd4da1324353389c52544ca371ab895ab6c35cb38aae68cc765342861bbde3a1968aad85395bd1ac1309f08c460fee6e4e1d30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4165e2db22bd3e9a7c232b7915a1fd3b18e3a009e8d006b48460ae2df22dec2a28aacebf781ac0e8923ec097bc49d44a824202c04f642e2732edc944cce79df2a3330b104464e72ce3af1d91efd476e69d96e819b9c0412e773393;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15720be9c672368d546a1a6a729984d7fcf4ce7681351c4a2426874e5310aee5f45ad87b6f12b5c8cd6d9873c7b8d0a4e69fda4a5264d67e772ab8d5969315ac47336cd3d7f739d9870980f1ae167dcae5179ceef84b67c95d3f9ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d82536953fd85ca7b2fdc810a35cbf817c3aaca4b5668dafea11627c5f9257b70f67672d28db7da468a6de6a88fdf3561ed9c4650ad0b79835099341fd2395349d672c0301e03c17823ddf293fa7fe96750c34f98a0b962e25bbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e93b9796777989a2335bcca428c15c61d29d99cacce950ec03d60b5d3a7cf740096948ebdf0fca7eab60a029ed77e4a10cca3bbd95f750d0d67844c1a65f4843845e6ede33d8d0432574c2e1749dc517a5c6596ca2ad0f491e0b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3aed564a234e0ef283fb56574e5a3b1eb9162a89f3622865cffa2f4184c81a67d912d2283cd1b5b54014e1bc9e84aa8bce7d77f59d80d762207eb08615c64081989ca19618e13743af8f7a0da54d694105957d70e97b30352739ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a08698ce6f23b6b33d933ec782b01a6e03ab744cac508f308698262e24389f2f60861601f59e0b9173e480b4cfad7a6a651133425b05950d3f349eb47d20feb6947522278cb3d9d3052274e0b9359b66e51725adb773855859a16a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ed61d5654f28463ccb975d1705580bfe4fbac26bd066fcab18480d579fd186b236637baf77481232ad4576ce5aa400ce7e0a750f55c93c5672785f055a98a4b329c40c17372d4bed8f0fbc881f26c60fcc7719bf48116f968e04e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea31663bc476affe0da875f4ffd891ee964b4aecd9cd1ca672f5f29dce97419daab503f38e4063de496c33c5c5761e791954fc4f26b081af885014303fa5b56d190267626ef5c04376fee4b4625d2208ecc1daeef4e67a35eda4e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he32f487e40cd201edbc939f7339cb82f9762d9b7bf0455cf82ee4031feaf31fc936c9ab3fde6dcb7fa8d6a53e347eecbbe37d40818cb0f52f46ed3f906fa9ffd97ebc250be26db15253e3dc820dbb0997f8ff2653a2c381ce0561b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6be6477a540d6a0cae4e277db60b200fb18b3007ba36cda22e2eac540b5ee12c50652954c80b47378903304798203a99e97b4ccbc6a686924c478ca45777630649820ac62142b53ff4f8bb6a347c7479b0dc4e346a2ba679059dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1701881916e6da794e1c524a07716d7852ba3f341dd1d6deebca4208c7d3a0801d7b1475c3f38712dff1f928ee46d2342fe7ead1779ddcc4dc4296d41bf9c99d743b174a0d15e55738294bfdc2f015f6edcc7af600b40048b18324d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194267f5c3f3090b2ce300b613b65ac2d4aa9a4ed7f645f624989531fa859875a14cc4934ad33bf4fa542259008da2eafa8641ffffb9fe1306554125e644260115a6b7dfa7f322969cb22dccce2148995f3d0d7cab795b2c04c4012;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cfc7e71fa57646600f11f9be36a5264a058a9afc8de9245e6e0204ee208aa2f6e2bde6d814c07f675ecd9eda7ecdea5c45da660cc81e3649662b062b049f92c4912c248479365f41adb6ac195a64cf0d867711d64b2af2d034ef45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f14990913a567a7d0a1325090b723a0fa8071b131606ed988f5e72fea7c327a14199f2d6c1d4a0e5f9101df3696251c45506f0f2ebea822f76e55330701f069cba412c61a8973c276aa6c53067f6c1deae21cae886e9bda9c87240;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cdab68b558bc064391d4e0ed3a63d821c43079b550ca0b377607e9deddce59ef0f89783661c5355db2113e733f05b0961208c768266a2ece54ae429ececd52e17f4e2396bcc2eebd89a02643cde2f1bdfa040a1192e1b4bbf94a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1490782d3446b8595eaf66c6d31b9ae18d127ebb21b337fbfeab446cced6ae39c412c7e7294a694c7f88862a636153a4b564e846196fb762a6e8befdd680748dc352e9946d5a31d4a208d1b518509c4d87ad54ccf1cb40686e1440d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181d6b8fce0da9f1a66b30d14323085ce443347add7b869f3eadf3b079003fffb8f29e7d5e4d197d89d5f2da917991318eb44b178362684dd36f7a853494e98d369070c0887e5fe312a7f9121a1af055f3d804d61dd27bf48611c37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4b548c897fc1bb4be947ea5cf5641c8f28516cf30f8010a73c566343aadf5121324d3fbd4edfd86928844ab5270c7b696f7918b6ae9ccd111d35b0a06cf32452372b517e3e595b40adfc96ebb442784146548e5b9571c7af2998;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159df8cf99eb804b2d1ce3ff8a26d7ed7b70b0002b9380e5afea3f6380217868f45f841964ea511f2eb9848d65ed4cc5ba8551663864fe4620ae44f1b621285942a2b95e1935c943e8f32be2b08b32e2c49fc0bda98238109efbda5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1097e279f90124ca5a350c1385b8a2acdadc162e0dc28a3532be3019cb03d68a67a195790b3486499696e598dcdb256f48db23239af9167da2bd33406f6b1f68bbceefff3f10e7acecf647eb7fb8b118153e3d6ac63d44ef5cf5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4cb7a8224ad173b1e1a1303427de302f4cf3334c2bfdbf8e8d901ee353b55f2bd75e39c957099d2affb1440954c111665167e3c22de288d0d5ca9cf433b37109b4b335a7e4676d776bbd76678a1ec2884daf180605a20096ddcea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee2ee4d8ec447d5b4327dedc2f50a80a9a142bfe6c3295d25d6cbb52235907f7cccfbedde490c2300cc7d1e093b8fe0ed50092851f3eddd9778541c207f4ca470d7af8e2ada6d6c8f35b8bd230ba30d18af3e64744ce368224fce1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h331453342bfe5616f872ffed3a2db29f07115e85bec1086b338b8ff3cfc557a6e8b33177a3f0b524021109f398a3dc3df239df25b5310f778e976bcc57f274838e4ce92a94f5441e7c90ac8de65d2faa3fd983697cfd9ac18f8ad7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cd9d40d3910dfdc2ab4813f1b0ea411ef500e531e03ef315329f44d5b8da5af2cad2c1eb8161b44bc9ce68ecba0bc384030fc501beab2a75caecaeab1f8146a5e863d9b732b3746673be34507c1a2de10397e40a4d272daae2e11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5102db02dee1d8fadfc1b16fc168997855f057253138e5fac2f149dba08fdafaf61fbdaff0f2bc3b76375a6b957b71653bff998358e8c34c1b2c0778ba510564b3342648a8c1dbf7ff2ab63faab185b28d86d6655541857ab9ed40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bf924593a260b82fa71d0b16bb0329be66bac5fd7d1528e92c35543933addc13a1b37684faec6134f13e862f4a7104c8efab98cffa894188a24f5b21fb734a2609d70606b218b2d36164a43ca7001112e70fa65dd8bf243be120d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fc463c4e936071e983abc9965f3bb0ca12b3a5c065c42e8a26d84a84003f9a3778ec581b067ab5a6edcb62a2a7888cc46c6429e02c472dea843c2a9929fb7d6837c2d9e1c2325bc07846c18c712f1fa70c9f84c422584c9c2f2b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156c867c3410284a8097581d19f482bb039b77c4ff92bc2e9d2d5a16a9fc738fc22278582662b200aebd7798960f43fed4df4319bb6c713fcb44f6acb780a9e6cd95fabb847010443779c0fa49dc838f141ff1098ea8dab266da742;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4667f64dff5768831c2655dc95bb55ac953d25e73b095624e431fac243ec9bd62d5f6ad08a4d4cafe293de46e6a5a296489a3780846f4bd47fd07f0b2f1765540e2d116850edc875a3b7fd13f0997870aa67694303b0da0772df9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1076e17f44cc1ff2349e504003d6fdbd7f8ae07ecba676247eba0c96a2c2f3fee27159958959c00f4cfb43bad7a9fecaa57b8aed3572158da4e861cdb6ccf55c1ce29c1d076af25b0e908bb800f652e8ac10fc2884876172278096a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h213c26023004a1479c80de97c1dc570568e23e2777a8b2cb45f96317a036029baf1fe84f0688741f3444d24bcec8b3994fb836987ac97c3fb69e759ff41f1569e46ff1b009209625debaf12a0b5a638e94a64f36b836f286773bc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5b9b59afdfa313e1b7dfcff28672c3113ff906093d5ba812b3f2a34126ee1f585576ed9ccedf4c9526f71fe5950c3e4b207d9fb98496e65eb87136ed048c82163868713de0f2049cbd9a9b9c05d5016e07a8419b8046228c29f9d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b9aa0d79aa54ef0738cb5635b55d88f97390401cd7e50e7878ce5b435153888245d02dd231b0e42577a60a5c1dd48f413d52f9bfe7ec3e53eab4e2b7b8fe8bac983a2101346e39b5f0844d6e57c7daeeeb82bb4c9e54f18f81247;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec613e2911e7a6401d112b5a6dd15fc5ab3170ca939e60b4065dde508ffe5c7d2710649a0911ef2abaa7e0379c964f007cbfdb7e7315c67082dec731c4813b4425a19d9de50ebc5a0230db5cc423062dedf63673a1dd805a9f85c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9936bd8b0e5396cd6c9cfee0341bd0e4cb464b1794dbdbcbf2496ffdbe07ac8b6df204d2649c79c0089315cafc9ed215aa7551322f531861ae08d67660dd98f7e774f09010ddccd1c927e2e307b4b11fee824e914dd2b3aaca442;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bab3cc0a715ed49b13688b2a6b4edb093430a99a78c674028935f6ad95c1601fa29c881607dc8278dd1fa6bbf1e48a1b25a1099a63693bf30f5cf557049cb9fb384e5b69f1907d0c3cb8e71d2f1d120bd9e76f7b49ecc41a7823;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d387781915d2cd45c2510f800adf565714180bab2cf471159175847eb08c05bf67708fa2ad5ac533295bdc7b15cbbe5608e0a64e90b5e1638d2a6e6eec4a2add0dfbcb2f903e2ac7c4d7608420ad4e67922bc2b1c2cb355d909db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h116357f9dc1a1af495d0c8d9533bd80ccb63562ed7370186578c0395f5298b1a47136f6eddaf95000e45b4027f84a2bf3448ee208156f8b5634ab69a51d71bde1760e8ff85549f1e535dcc35eb405b31e913d585462e36d6ecba12c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a94d3ff42967c6fc7cf710a095f8aceefd653c34cb71a0096a0f3d6933e03dc3feb754766541e2cf3467c33babe0d196fcc82225ea92d790ad00483c9873b914dffb69acbe7b6ebd7e9f9436d8b8796762a242a6e0db687ce3a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77c07f72d2f15b0f96f1a0bdf4b1383914974b6543b0e83f4e5e7e7bd0af3688b2ef29fa5cf3ea235e5b57ba9c542ff0bd25fbca160d9763ebb095bb067fd9dfa570e815b049f0fff90fa2f435a895e6f97ec5e76cb993cfbe4a5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6c4330ab6766c1be2288479900814962cd53acb6ccb137140be84840eeb41c92b3d657171a5f918bae87b6f9a4c1736799a838323973df1df46ba7b001a17ec343aa06880d3cc3f42c1680ad3f77574ccdb105e6e9c969f0e142c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5895ff04b027a5b02a9585732187a34c605ceca313e0a61b9815ea72ddad813dd4c4751161a3b23ec747de4ea3d8d67e011d713b983c0181816c6a9ba616c2c2761cacb543735d730f0f4b8d10485b24bbd72673074d80c0009eb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92fcb384941ae82635fe2c67d5adfe4feffe5a90645d0d50564f0067419b2c2cb3ab78ecb90504ad7c3048134142cc5869fa891d53636b31a312ff12340b8d5c654102c319fcdb0f1d6293f922c5c51219b0252c40dbab87f9a88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c6c8c62972a3daf86c3e2e0612e3f1bedabfba9518cdd35a8abc748d4669d8636202b1b62925c6228a07d51a5fb8bcdceca3eb020ec8a6b5cab58da1ffa6df0f1374842843aa4de1a925c6c1773573d5f83bdefd2a633d4a80622;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eb10ab39d7d80e1d9aafa98f39cd925c521a05bdd8cb71c9ded16bdb70a0f48247ac7581dc9f3ec85d258e4e41927a0a9680a28e51551a14025657b422a87b815a1b3ee62f165b885c5ca2bf096b688b287e5fd4fbe9b3da580f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173806dea439028c462ed4689bf012f4094fad38c9ee0e696ae8cdc7d791a71d2f29541800723cc3bc61113e7d8ba2df8f577577d3ba79c8877d0ec1257d525895aba2178119c0c4266848cd9111fdfa4501370a3743635b0978e76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fc0f0223304747eecf28f84abd836d530113ccc9ae21b94a02a84d0d557c2dcae6dd23b2c0a646db47d28d3af716683b1a53b9c25ce9190dd3de6df096518a3a3ab224be6fa2a7ac15c0549a33e5fbe3ca75d1b474f779a3ad5fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fc82ab10da59d6962e407270ac5a2023dc36526edabb3d2d3b4ef13ba87e189ac18db64e5f77e69ffd5d4aa339b3c3733f37d718be25e57e9fb6c77627a7149484ef5edc0af585c07048fb1a5390f9519ce9994d74875d382e78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142481e0208036133f78947c7e4f15a7f0373b9aa88773a08c7523dab08f9ba0ec86e72ac391cb19c10a6382457c15bf8760c409e8d15c1eb0562ccbd32282abb48ba639ca9936f0a7f179ce30e97074ff6bf89539f9fd176d0ffa9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf21bbdc0031557b69eb8435ea73089d11bb2b76426414ead5953f8792ddb8dc253109dc8b88292b08b49f81867c6b015a807d030b5bb040babebbab72b0c6b5e349427505069337aaceefc29acc22c79a50470b2da934a6f191b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ec07abd712338975dbe15301ad466a86032b380c1e59298e109bc323ba0d4f4b8c06f6396987ea23212b95361312bff46d4cca6cffaf51136d5c74ca62c2f75d1e89b5b128e9160f95e7c40acf88c6b97d53f83460a83dbfdfa91;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189a2b5b4850bc4d38665f61711a9e614109e669df375ee6727873ab49e7f837203544003fccc8ec9e82b08e4c3c11030827f90bfaab3e564f1a7a6ac25dc90e13e16827d0f00e5b778116712091b86729760f4c00735d323b1497;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab5df4cf761e53cadf67bc5955c3ccc85802b17c13ef5a32ad9e51aca842cec38d7a76a873bffa53edf51275fb0d924d4707c7bd7f7b587be41a0b8a70ef85735cd13a8e6989fcde018184bc00e8b019f936bad5a0275ff3576a6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc5d087452040d0f836a7fb15098d615d5bc3313eccce0f9364078e0caa5036c3d63c3c3a65c4a79056e9d54be0ec1fb5dffa4da7e42a65ed54861aeaea067260e0436c56a62fe09e8e6742fa8ac67a51f67c4d3125b1ee756ae3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c77529bed1fe0a61dee8bf2189215950541a2ed22f04f398e9c0426399b3d9d5b64706b9c3d695f559928c667414af3cdd0cf69245030bb2a981b96a0faa56790a4defcc4c59746cf2e5f97ca06181e472476cffab12ff7a40408;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ba7183ca70394152991abade0d2851201499f22920810bdb0370d6eeb9cd775601e4037efce1fefd04467894f2e10331081e93716c468b38ed05239f2973b314ba30b889be3904297dc8ee84f72d53a1809b45955c98f1cbb0c9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129b44f63f40a9e6e95902f3579ea8b815b00effb5ee836f4ebfae4fca2f379fc501bcccd42188989b1d8faa3463a6abcc563c4fc45cb317e2d8c88b9e6baacfd9161c142b07536c351225d75afab1fa236ff568f57905e4028c37e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137f6a632e55e30ae438ac0223d5c2ab06882ece6a962f71b34c4f69228f3f0e28510daca747d8489a2665b2b87f368aac29d5eda1b31699acc1d8a8bc0d8fc010f0948e51eebfaaf2bc64bb0eb9dce2da2b3e24a8ffafd43552d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb81cb1c034f7c9c90bf83f6e9a188be637f4404ff019bfbcf453a28132b809420b045eb986cfb2be0fe9ec795ebd7ebec4fd5ac6d6c60258061be0e44007bfac4a3b17cb0a4bd47ef9218ef856cb63a728db6d2eaf00c65425b2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9202b246c94dc781b52ab6701baf852f8cc69808a11e742e8586e3bae5628fec3cc2ed9764730969653c44a73b4f30167b7ee079d3a14174edc7385bb3c56a190c874dbf5c5b97e0924b2ff29c50ad27aacc933931ccd8e4b29d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e988668a2fcc434e6c82d289fd833b6110c480e7ab43b9dd702306274a447fa1751007f828d9b13f7d95f2df959db0184e52c5809214748ddf85030a61ebb0f36634a865799e87a37d59e1f37eaeb74bc77cab18403fcd16d77a85;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ed8eedc5916e989397dbd0876b7c88b84a9fe00178664099710c99c3ee107fb9a33fce5cda24d25c807a2240520c2a55a1af2234a38d4feacdfb8995a0b3d41cb6d03c3b6cf4333bc4bb7001d303dffaa6af917d696b38f961c17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cba95f9edf2e0ed1255aca6f7f7c302376b850b4e5ab452879a5992cbe5c7e403bd56691d84e00110a10b08ac2f5879dc0ebb73bf7d341692974797292abb2aeab3cf7a976c98b9ccd93d71467cf77567fa462d5fc98d2486a7f3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd70d82ea84589ef5ef80cde91bbba9139c62fb9e1dc48a01573d326c37c06c73726eda7ead5cc238c01cbcab973c0dfc4ee63996a284f70e8b6af022eaacea407acb6c7797a8a1086282eedde82f9add80b18ac76ddb808f096487;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9cee01a7ac72a7ad56f7693ec70a58d3eb64997b9aaec175e33b9745cb3029a85a83836287d141627834209931eb1550abc1d17fce080e5a1008d5b618ff584cc9d03e5dbac1a2651a81e576a1da66456ee928144cdda3032ee7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108dbe6bcc6c487fa51abdf01f8eef4d5f58041d7ae55c29e4045f29e1f283a36b247cf86ef25083cd3b1659f555f5c7637009fe2871d8fb609cc0de95907ada72a70f655d70e222cf360ea4d0987883c8a755ae9e3e87f1850e17e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e7d27f3d9fa160f022cf2f247e4da75c01077daef8fd1dd270595f19a6f57be997ea89fda6e3dc2b3de625e843b34450dd3d4a4e9c93f4414d8c2ccc72fd677d0f90efa0926e1550e718148e7dd3a31c5564c495ad1300cbff19b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13deee0cf1fdb1a2553fed98b59abf9c2e86ca76f803f660d4ae6fd56264b74c502c1e9e9a41c2af98d8b8049b55234529d3799423d4cb8bf2ee3f8581b18506279f084407b1223124e96e332e5d1eaf820fa70a3726d3ac49dcf71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91b41c47ed5d3ae38d452a44d635a88b23c174917e057b289f2c4c08d10a04f7767e00603ed04ef6003571c54d4d861acc964b8d4869ccd8ab6476b90fbffadeede0f036cdff8a4655a9aaf269595e1e16967c289199551697b0f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65b8b2ce7d59e74ebce6fd7853841c3e4368e0d60692ba266db5f816c7bd84bca4fbeaabfe630583410b4823744cb9e26b147af663cef922293af13c0bb59dd7d77789338332277d26e5cc31258d09fda497bc41e4a9b3742f90eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6e6095535b8d6ebe9f21b7d9732c3422d3f4335735c0cc2bc607dfed53d643bf274362e0dc9eab2b807757b0cd9039931ce7ec93debd9b77438991f3800fc9849087e76c2aac596562b630cf4ba51a7cef1751c0a285455e98c139;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109460beaeb8d3210975c6220ac081ad53857b32d99a00e310d5644e18d2f99dad3f4a72dca46028b0b0f37baf777cba5c2c3f3abef46d412778eab4e8ef2f39c2033bc8ea480ebcc7d82d06e826d6c229ba04fd0e438b22df8b8df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8684d7233884e8632285047e623b157ae6fc6e4a7abfb1cf7c13e8402721b52c1022eb5c7e0ee5963d3f8d451ccf3d18492fa82f9c75fb2b2e9af1bc17685f0bcff95ed324958700bacd56d68a4a37502bc75311c25d0c05e4f4d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101425415ab850e3ba85640377b0efa5b6cbea6bb3fa374615b3be7972670df09b03b7c55618a8b4911d0b7cb14e8c3760e099275224d493390916f6341645e994c43cad77ae115e29d778004c9815ad4c24e74aad3b1a67be6ae07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4efd8f527184638e1c6513fde15fbca5d76189a24ed1b4f674886dff7b52a6a1c0531b4a5b32e85d8ce085bde6c37c78c5b4165bad44679e827b5a8e8c69936dc474a72b4e25ce3bcaef7ee82a5efd8ea8636139eb0ab79b13378;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ad3c53971463566584060a0656a0ad3006cb7e84657a7f7e69df5835c17c45913cdf6ea249132d02b877cda15bdc0f2f14d1dabb7b37c146152f82ca14b29f19a7041024c81efe25ca62972e213424bde1120c62ccf4b9aec979f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3b3502d3538b84c552cfb7b640f2a44d2d09920342868df412a6637b912f27ff2a3c8cdfa9c49ec5d55d990f46e0faa6a14a1ed1d735bf10d6914be59578d664e46f472cc67ed56bec76e49b2d3c942c8fd74602c9cae2de1b27e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3660cfdad043307c15e85604dc5689266ecf4a785677ee82a0a99f96ac833f5182ad9ab37e831f4b93bb187abbc37c04d5bc3650592ca935b46bf50b65e1daa9756869bb9a6121f21c3b11b16866e7890a6e35fc719db5836ec01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e42b2d9b75762afefd41fcc8a6df8e8c8d945bf028be6a3bd2278cd9a08a2483480632485f28a408773689f77ed76e061a82161e6fd5defcb4959bfab171828d738550003b1898cfe324747418fc533603261724771a363d19431;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53ae25cfb44d5fadd2cd7cc16d9224134419b0ddbc4b6d4a5546eb3db9c83b79ceba3667e64380655f9aeb8b25da72d8836e2616437a16a7a9dd1fbb3cd5abaf817d9c3aa4ddee039ec2c8de7925da14555d7937f680eb6d1940cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18772be95ac5232f2cc1af5796b4c8367046a664b7223be5222f3198c62e30ef8c8dfc9c29b9958fdee5ad18e0b093806b9b9ecd4b2f41b57040a1c5d55e131de8a8f0458ad518d9bcb4b1940179a76781d71d2464a1e435bd6b1c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10710050774baa2ec0bc785b52c2a771ed2c8b9ce6213a13bf702ff3ed695c8d1742a190fd9a24412f304e064707e3ffda721593897a2d68d69ddbf02c913ab761c40b9f04e46e8ca15beeb545682b1670b9ce0f6429a2c08392f5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf3a098cdfa1e0da1431f8518261e2f3b530e6e32705218a5d9be528b5f72eec74c6925a88a218ac26eb16a109dff0bb520eef7dfc042b6b85d6c46fc16561cd8ed24fb2ed6a24687b5a181ba8a1dc3279edb0cd39e197e925973d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ee2e4fa195a18d2fd0a70264c109c7d145d3a3117c3a14e5027e8e77985968617a9fda7d8df265eb1054e6d45dd8cdbf1146a5a3187a0ad07f861321bd3a7f6f5619e2d553b3471c403565c5c864e2efc8a508e86b4ca58fac8b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h309c3667c045b6bc5e056d02b64f59dc5cb84635dc15e42393262ae3d52d2a70843a3667fc524d8e91c47ff9652feca9fc9b0d1fd2235f623d22a997c91995cffa56ab204835991a87406f078f68f0caadbcc0efedc69e66a55ccc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h554073143ef283591231935e7339675448570d55bdf09c7536cd4fb1903967fc10f7eff8284ebc4962f42b9c57621b9718c8a799ac91faaa936e708cfa3251a9c8ba9b5ef0abdffd0e2d76842b6b320e9ef587c4edfa486b40507e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27ee7773e821280eac93fcd660d017b08a344be674314f7a02dbdeddb8de3a3e3335b549c1b0f8f9e5655a0070c5241687ae2e8c7d945c202eca966ac0922295b25616a730f400d5b4c7ef9dd2d09ef051df69ee5a61d97baad3a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4057dcdb16280dc147d4825e3b8c75a7eb89f9c8d5fb81a4da19c5768591a31203c456e025ff8a2c3342b5cd214cbc38aa4bfb18a71c86f357085d0c679e21ef18c93ac5e7ccb4ca01e233f232e048b975657a3c485fccbcfc0df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a006837a457f625c088bb3a544080391b9e6c0cf15d93649622b0b0b2eecc555747683e045889c440b341799c27f288d5af954af091ab5a29c2a9ac99088c7093ff1a90f15c1fba8f30dff7b9ec0d300ff239cdf67bde30ce4e45a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142e59fbff73eac87fbf570a29f849becd0fdd8d18a61ad651d36c9b4176d7c10381dd40c4019dcc6d420ef4a34c8a17427df935c9c176eefcdc3192aee501f712561f8289a319f4ba0e50b1c63ea399a405be3057c2e053081bb77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4c969772359153d62dc61c0a71c18e27e22cd86dbb321d8a2541c080ff7f79d47b66068a0684c3a05cac5674f7e9f691b38feddee7ae15b3a380b328f8a5219df4398304a05b08ddfd90aa85f116ab2e71985838a9298137d7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d94568cb8d1e9e64a817d964677abf45a81aaa4de89ceab6369b18d317c3be7da644153226e04eaecc2473273d47b1f495958f96183321e70b7fc00cbec08feabaf4cd6266f39646784b26f0a504410aab42657ff6f33365156b1c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f96326feb96d2ce923ffcadf3a640e12c332c39a4186b5f4f7f0c762199d05dbf47fd5f530eec17c8551aac3b6cf7df7ab2f4125379bf79a4b12ceb4bee0b4e610874646b5be1717274ee8d3d68593cd193c08e6bb6889a9cc3d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64407bbcefef29423195cd422bdd88d4bc48556715c600acad4476b630e615e02454758ea7541de5b1c3c3a823199aa86813e34259c9d2544bda9b2104fa74032a3a88fddf75df9c0c054ab5165136c22a5bfb8c2740180391d765;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1253935db654b70d365c00c18aa9e15aa1f59205b9d81ca4dc1dc2e6e321955c5b0c87d554e1f09351235f79e653549db89cb1457eef55a86e94da8ac8324903725901e6667ac18a9dfc5e55c3169b600b2025afba0bc5d8b253786;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcce7c0aac238af92c5064583fc0ed8cd270708800c2a7ff04eedb5fb86d861b647656dc7b2d4f2ccb2744e4de5e0765b854e8e64c9ce745aa332fdabfba262e214cdfcab9321cbfb6ebfe36ba8696dfc5e027ff6cb5e06c15a09ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf662e5f6f0e6304fc9250b08f479ed46b4bb511eebac7e56de6833e8108d9d2183c7976a46f75551ddb55d8fbc67636781131518b4e42117f3fdd4194c8f44c2e62ce028b16efcdfd37e45b80edebec72438af80d21b63df30d817;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf112945bd3535ce98c3b07af18ad83b25d3ef261a7530cb211ecf3d15406476aaaa1d77a85529bd5bd4a3dec15d6ef2d94dd410f167eba298c6a69afd2b27db47747430459f273a4ac1760160ed9fd0071243798aabae7442b6c9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2050130dfc138fcb7e0c405f14ee5700a6d0d2e3982314014f0f07883448c3af58befc9d8f7fb64124ab2984051f5103537b1812fb5475285a91e3a92a171110167ebf18b8691657738bfecbe1796e847bac80a9ce4f46fe23a56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1938d9a0b79aa02bdc04dddfebb6d4b03a97a7492c2b94c49399595c7c1c523a4596c93e023dfe08128c83a0595561122c1af8df1160a50a8965c57db18dd11a5440f0470b7442d7704e64d1093bd6d72cfce020ce745e88f5dc221;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bccaa6d43497b404506bab87be0250f2338e7f6e626deca7d8dc525e8c05cd627ffad80320cf809a59042ef235fb3872bf17224b8473852b70ee74b145e53f08f3468feea74f03c5439dd556745ce7be6490197b642a205d19365;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160d0d36c8e59e7a280a3ba3aa56f06d8552f43c09f2f49bea0d38f84806e0d85ec71d2703b06f0a8167c6b47642cfeaf8a8706ecb3c5fb7af29836ae4a55e7d947abb7d70b3088b81843c53f2bf60c377b37760f7f168df730d5c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a34bc8260cc3b0bf882b7bd70fe66562ea664d59c7d369d72d97484d1da7e0016c20438a77f01d31c1651f46b634a24be54a9acf68574c42efb307be04c090e9e5de9f28817317f231171438f399086fba9f938eac098f2530155;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61e3a2eedb0742abd58b6608b8b87668a9806e7cbb42003142716aa4119f84ce05521b0cf0c3f42823507944aaa64f498b8ac7d06f4b1bb2b795c77c3cf7346e0e33ca14689cb825b47b9dd0f6af3ddcacd7a9c548c8e64ae677cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f3c80222235de080213dfb8812061d81d7c980aeec214cae7b4300b3fd05f1f86f814c73031aef03a5f3970c03719a964c370369eee0cef5a83875a338351d84581d4adf9c6376b6b23ed9b6c9ffba2cb5304eda6a8155a2b5bd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1835bb142a5dda8eed6a65b3386c2452bdd06d665bd5df047a87a26e87cb3da3525b487f823eea404f034cf0b4aca65656f962e10e54a8b079c3a6da16439ef693d804c95706e6bc5b0cc5d602882ef66f30ad390bb4a065f5f9ac2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5160510b0d2b7ef50456da5bfdcb37cfa77e7afab2d6a3d482461f98280827e9c86f32acf59ccda4ba1500f430a6b9a24ed4b0c41885e8f8c810fa669a46ebead3a20edfd696d4f83654bc185de7f6b699a226881ca850dc33412;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef40979cc35d9cdbaa0bf0776f815f87414a1feaedeedf77c5b0bdb50f454e97ad7d0feefdff4d6fec3cd3d68f98f71d855b955ffda4539f792c2b243905a9a0b79be3494e34048209bc13b71126b8b4f96bc6b4f0df651fd89219;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bc1876bd64fc1c70ce469cd8b37c760db7d02b40bcac56751d2c8f6ae0f2ec39530d1b02c1c38a2d382cbce5e317da3ff78da22b0daabf431e74067bda8dcaba85f2bf504e2b98bfe68ebb1498c28cfb55735160b0b5b61e50750;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90c50db3cabe6719d2d2a51805c719483c562d6e8bfb90921ee6d5a8c8d445b015915f00b8bb82303626e40280a27d86c38e3cc646cfd9c4a3c902f69933dfe0f678504b080f7c4a8e5cdb2ee571f5d9f502319e3d04d30302b632;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fd2aeccd35c87b2dff51015086e328fdff6e88f2330dab6c20bd679db1a48d3e273864006709a9f7a9a80e5a059133ee09eddc0b98d0ef16ad882111df1525a828557e4fc0f406aa128090fd5ed6fc501fa58936a3053b44c1f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23c9e9addab10c2f7e366f06ef8ba0ce9bc22728251a003458a8c952e7540c50d0f4cc6b0fec3b0d897a7a2e39a4a876fb91a08c0907e1651a00f748223bd9c7e7a9315ea0649fe76e628025322dac5b92ddfb734582d9082d3d50;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fc4f12031c2ead80d51cca8c3ffd0da3d87266ca10e6a36dfe65436eae641ac73e0c1a9b5431dc12077436bed7128f9a66868a2fca1329816453077f53d3bc49ef5d9531ef22833431da105568aca28977a0cba608203bf4e9f54;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dbfa936ee9dbaf12f1b61e32325ea8947f45836bc55d024f6644c3bb5a47cde1b734ee83355ad244fd71787954e804828ebc3151bde175b9f55a4743274804dbabb8727edb6917de726cbd8e4abc8ab415b73efee71879a5013387;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c594c02855c71f073c92d052d9fce74a34e27491ac139951c69e9680ef7d35e48ec1744d09f123470a0388022e312e6ea6eadd2f0382948fe94a78dc815e23d88519ee8ce0eb78110fbfe749eb8b09383638a2dfa75965218049df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h672130eaaa6fa956ce1b96aeab7ca253fbbc79fbda270ac6ce309152667bf506020dc3c6b8cd748d43b57a0bdcb2fdf2f246999708689825b3df4030f39ceb8ea42f65349c57fc24f8f2c4e2cb6da20436862326ff4c01a7bcd91c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125ad747b902ac9f73573d7792a00a5706d8ef084017012797e40c5510bc4ff709faea79894c0f41f1cdc053c69b0dba65947d2a61aa8e3fae2db45bc97a6d269c83bd7fa50d2ea71f1a719e621704f880cb62b45bd7e6f579040e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1118d62bb5c55326040908729ac94da0c06152303fac2037ea40e47313392ed85e4b22c9dfb0866faafcb5d7992e2d42716afd3fc35aee81b81f9d8dbe8b3736189cc2217de9fb3151afccf0e512496f2b3729e545fa1ab20710af2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a29c08b50f0aae891b2fe8dd7d96ebf0d792b0cd81626d31846c7d93c137cbd48c3e7853cce3888ffcee231c3c48941cfadddf3bb34b87b51d93314fc155d085e737264b5bf6893775eedefd9cdc2eb67f655a85fdd6ef0312fc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf421f45c03a616c8f72cbf0be96e1640b0e7efbbe4974380adfea8b68dceb4a0cfc4a610ce111f94243729c2d52f9b20cb8832fc730bf5afdc3701577b3be0f4d53e7aac6520a862ae11cdd5e93fb719f769f3b149916ea9bf7641;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12cea1c9348e1f806ec79155cd4c7eb78aea688eca83f87552aa27ff473f933e08ad7ad0783cf2955822be1041796760d35c0f07250b5a238dc26e4ff55adfe2f4d6cf2df88f2465ce52055f39ed786e12242b83f1435d579d31ac9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1adcf739c85f94d54e66b22140693da6a9690fad31b012e3056ad67a8c905f11e3dcb6ce3343a4e633eed1c40c54c94d2653deec5e4fcf5fbd1743e9a718f35285bfee30a3fbc5be2be9d5f3bf9157e983a85b2bcefcaadc853387b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152cbc50ef62304c55547503172d274034d3e97c90fc96b4d6cc4af64ff71dbaf0cabfc7f336829d6c00abef0457e184f52dfc30168ce687ddf3a25ba393db1ae991924faf0f2833e593dc86155dd8b15685cc68e8d05a91fc3c95d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f54c954a2f3146afc1d1d35406a9c7bbabc2e629da43df37e9edf862be77c298c866d5b4d753b9acc9d0c59aa4d2ae654ce6e097460b40144bebfc962a10cdf96d49ffa73ce8c295fbd5181344ed6672b915fe4fc783044c019bdc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9a18ff9eafc338b6e0fa3151b118116ab73b60c1ddaad7bf80fa6a9e246d2a6abb77dafe6f89765e0a7e1ee63eebb1b865c267c5419c13834b11c72875477673c968438b401f50790b90ab981d78e478feee00e76b4c48680f82e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f950aa681b7fcd7d254666fabbe0333d694388be1e5755a16ceeab0244d648fe18b4fc5e6175e4996c5dbcdec1487ea67c905fbc5cd7180743be4eb020bd1f3c565ea09a2a31fa29da4518b50f1528faba6d6f9edc2bab9c4de1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa244dea706b9288afc2def4e616f9607b98abcc09065bdc755220553644b9b47d8bbf97fc7b7102496692dda1c1eab038fb29913bae22be0075cb3da291790c473be9de9e309bbd59d69ffe9ccd5603b1ab4b92b8d98140405468;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9848d32e4f9715d3aed3e87e6aa88671c48afb109a5c1e894afc71e7dfa0f22649276e1583d5cd5df0e910b481c4eac29575de5f4e47fb96705afdc192b95828af55707e9b1377775b142201a9920f23a5e57bf3f37a901403fb10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fcee591f692bb536f1a9698411eb1bc1ac61a83bb01db644b66d32818aee1b6808f5c7d917c8be6410df06c4a724deeeb89dd082c89aed5fc5cbbe0103e7f24baadd34e81758d9cfb67e05c63d1d9aa0bb962ace07d65ad50f084;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15802817efdbb117636b85380697429c01a480b4492b958cfbd74e04a76fc4eed2a6303c67e6faf3a7308ff30012cda87df914d355fdba1532022a744c42dafc878a453cdb787f02bf3a3f7fdff53d40bc844c0e4d9ec4f1ed18282;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h435de0eb30d32c5eca83e5eda1b5c235e9fee7c880b950f8b6ec77e5036ca4f95d3436246f97165d7b3a78a1aac78b34238791504d3f4b55c81de21588bb3ed768e4b2378b56b5abf4d8a5f4a5fb4de814251710b6dade3752f09c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ccd8f51829e6ddacc876091d99ce99fe6811f4a47be8b798959b80c9ca0f5a66911401dfe3a4ac8294a7474a9d523dce0a25351b90ebd7cd60f5ae6f779064b0d3efce2a6d06c5dd9aa74f2e1bb990120f6a2766c8ea0650a7692;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195ac304214c765cfad45ef9a926ce236a9e9c549ee9e0a07435cf8006d8a5de61c3b0499d03a03b0d9a76e55dc726990b233081af552ca2a0bb5411fe01e668e2fc7347cdab94cadf64ab7c0dc2db76dba94eb320766c3c4547825;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf143a8f001a9a325b1d640104ed545fb897ce0fab63cb06522825dfe92ce06b756688c76744c1e73e023df2762cb9fe7f013a6c1eb8264d2db51a77bc2303428122b97728443aa03b4cbc50af47f2fa24a4fc5d4a325676112299f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147a553b4e9a48d9fc5eac873041910684a08eae0e3242c678e1da8ce61090825b67a6a570c385a7476ef71359b3e28f4f038061622e62584beb2507da7f12c54ac7743540b7a8eb600552b8208732195c0fbaad1d8870012252457;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h877afad143edadb1e0ef73a6d01254ec9f570facec1be49b82266adc6d2cd19bdb1262ba42ae63d07dbffb7d2d0983dff5f058c8d9d0f0a761fe336fef8d237b64b87a578307a376c2fa5e8ac7c03fdee0c1b6902c6a8b16317321;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd009a27ffe9b33b15afa3f5e33477f44668f7fea8ade7e4891b51d806bcec84b80bb8c1b9487fd322cf711282c053fe370805e4b098e3eb632fd31f1c3455212545a19f3f79eb44b4b2d42e8fb3fedf424fb4ab25d985b09b5cf30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha20d9a6e6fefb4f0afddd98642440d79ff7aa21c2687456d7c6602fa5a767763d62d79581a2048f1069a69d0a2eca98b3c919798287446f5a3f8cb1a8ab7c6772059ee57c0cb24f98e922850a2534706331c809fd05aa948cae9d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e140ad27eb55faf6426de53c88503dca2f2a9cf141f0b667bedf99859c1b9e817b34852b44f602b0e07bd2af04a2bd5d331a5ca092a8fdb639e12437c129834912fa3b25dcef9d5e9c45e08ed4f8ed19591e5a135f26547a15f9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fc67203b4283806e59f691d1c6636c86e2e5d913d30ffe64be726ba1489f904405801b2fb35fa87353985c64142a382504adf844c8fdf7b86ebc344944893d678e2772a50eaf2a0ef99be9f95299a538746ad1b54a179dd4a8a66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11690f7d23aaedf540dc749bec7c2be4bd6394d263065fbd3f87167bc4ae92bf4796f8f69d9bb0b69bb58c0a9600702fdd0b41ee520aa83053247dadfba7fdbd3f20bbad5eaefcdc46ef0c5a907a777c5feb7f276e1bfbb71551e92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9bf8124069b886dff19ba8653b2a5640d76358130c20c995d150a8e4b774f32afff2f3a8983b587d0fc7b4ee6da73b7c2890c812e4fd3e81c9b1f823e31284aaa1d4a4be3b51d91aa36511df57763fe140f7893e7ea54890328f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15250daf2bde92de4c9ba4d6ddaabda92e215e593020ad075e838f3c423f776d69821721ad7aac370375d70b47ccc0ec69fcc8f163aa844f0de75ac29c056203980611d8d978e71c6d6ae5a1f306a33dcac1cf8eadfbd64e3025eac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h762c71bd62513c9c20dea49e15125eee893ce0835dee77ff1f6ef084cdb2f7a8113920ff5a09bff8e7169939ffc5c89c9e6ca88987d79133854c4b94666e736e12e78dbc54d0817f1b6f97797baefba2d4c235c78836105b71a61e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcabde0f699197c4ddb0cf7bf8827f32cb434f6f508c03bf30b41d72fc734af12d4abf457a8bafab12f7fea832aaf20a0a5c6d312bff261bb4c27863c06ba4413d0cb3418834d97b9b38d0a093043596bc2a0c481dbbceab9f08d1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa448b9e7c156960360d53f65dddda3695ea5970b2c8dd20ec8d0d76c50d06f5468e355c28a86a8e42f1ece959a96bfc9c6b5b9bcffb3a977bed795dd244758a7909306051a4b0b561fb2d2be8934c28f1fe2f5f2fd5265a206069;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da1ea2c1266113e2e0bd062532499bf1fa0900fa937be27a49043409d3d688652cafae94390667c8b318fef1f8d5510ed74e333d8e9566b76779d319e9c0a47f21aa597f89e7fbbab9b6bb11e77e7b313f3cdf8a9b9b2ee63ad3a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1596abb8d160f6028bac215330fcf071fc48c1965f3c8fcdd4dbdc201fb8eccfdef9860a72e16d1a6b9c5b15e34c44a6f2d4bde0584d6adf592780b471036e3c52fceccae2fbbe6caf0d618a02ed3423a75431fc3cec9f0c44808ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfff2a27aca68e6a4f0096efcf8d9b2c17a7e11e2b7318c06fcd151c35a0b814358f4e23f8ded252fba9d38ab4776eecf2cf9c56414beb5a3bc7c0acdee3ce5663bc1c11d4a0d6725eb3a978ae7061f6376c084910e1cc31f06f76a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b220f5e525331bf636f7eeaacd4cfb12bde52c54dae2e8c0ddb146adf668f33ea8618b551518ad29be4b3a56e1da50a3390475298faa1b245fec05643e7e0a310cb825d875419b298f1ff4fe0cc043284adc32b51a5c5edb3002f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h991a5cb79cbeccfd779f44d75f4914251eba81c124ca16056e8a6902201a20003200acf5a2ee54327ad1c6f94283d9969092735c29e1d41ce5ea7cfc0b9c0fc362ebf542cb357a076a5535627195a731e2dfe0c8929ccf89f44086;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82e0944affc4b2c6c84be7fbe33d6515dfbbdae4e0d9cd12a96584266704dd77e63612738a826b06801f471b49b006a5f8bf13d330e0189da3b2d9c8406cc1ea6daa990a5b829c97aaaf76b64b909bf394e136af8bfa9d28acadd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1200e980fd9b8fb728a8989f4d883d86371fa43bb61e43af3ad047d722b840a7130049498bf7ea44959db9f68f4b5fdead2ca5f34e12eb0abca8dfe71f53160677c96b5f994343d430841539c29635a34ddb0c48dbfbd80fc859140;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9b3c90b8ef24ae840ff926f5cdd908071baa606f74b88f2b197ab7941f354130c22e5e2d22976dd2663602e69bc6263afeea19d4cf09677a83e2576cb8847538a43c69f841bc2e4c93392385b384f4c7cb1703013f66caa7ed84c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd54d5f2f70c0ebda16e6ca552c372e9203c0671791748f79a467255a3a043c4dcc3bfbef60d97c7274c2a318c1518413cbdd95bcf0cb901fc82a84df09931f34fb97fe6cb06823f10504f8761923b98bd97e4fc94f2ab52a31de68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1851a83fb70cd751a56e4b2df3199516deef93ec7357dde3068810c5b660a0e3a8b364783368da9649c5aca87593a1088fa7d864916c805319c385607b5cee87bf0e202c20fe45d6c4cef7643de03a66ce29d4e76bbbac2bcaa9d92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce49ba5765ab7ea12e184e0a661ed40f84f8123ce23093075835e09e20f641954ef5129411f16365945b77a7a2ad6ca6ace1bb21a3887f99448141f0068d678851ce46c6e104f8de107dae46817cdc07c94e6e6cd3357be5190cd6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14daf8688123c98c75de8413ececdacd25555cab412e8fd45457a4410d03452896a49cf363c91c75070bba2c14d962f06d1b4acc138b047ff24b9172d7ed9af647ceced21f65b63ede1c8acc47a4642d4b41c4594a7c62d088e35d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h751548b2f66c9f589a8c2a46e6ca4ac8ff07804bc2aad662b5c9736304c31cb72f321e699aec5f2071d782ef2bf3c2015d3092374411d1853a1557247b225f84419117eea894fa020e989f7e531456616d674c07359496ec6e337f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83fede4774f1cbfdfa68900b7a53ac5c07ba8b1e933e270f813a160b777dfbd709397b060afd6f3e3f37b0181c1b0244c4358fda52a46195e46bbc8d8407cb0fc8c60069efe1017e8f4f6f599bf52feeb9a3a9d45795000693afe4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e34c64931ed37b04e5ab7a5cfaaea63da4b901f8cdd389fcd88ba3bc3760fc84817d122b7686bc913273ea9cbe1798263f07e2d2282d6b409ea8e7138314ce61c1d005fd29244e4b9e74f82459253d16fa991c0682e34183d33a8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6796f52bb9b37a4115b9260d653a67bb89cdd85321415baaec204f875e0e5749af0dc1a684392d6713b4124ff5d98a4c2fb98312d9949c0c5b57f29188db2137537d7b7bda45f7a01b884022f40b16cf99333fcdf255cafb21c70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a85f88f1d28d361c67f343645b87b50a5aedc6c9c3bf575b60a0c6ad9cc53e8b75b6d4afa34948105a6411a4cf13e34afef5ea5c03e21448544b7605013443ae60be70d3ce2830728420e21c64d70bc5ba74bb3e14b11e8a997088;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6ab906ee56006e55376fc24099f5f1ddf4f33bbeda7317871db2ec8853b25ed2a911e5706935ce54f52a1b4750b71eb3340c232941bb9ada3a77cad2165dc155418924396e18ea082bb74bce1b9c95be603c7120b1d5df298b78b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40e1b513818f546dd54a0f2029b765a31b266d2f55763400e3f4956e7c37ba9879085e33615627f5f200fbdf83e1f153231e312c246787867f0ce0ca6d293a096a7bf5599ec52ab880d16e3576851e5b3b02f79d330a5f6378c0e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h707e531849faf6740f3452e18a14cb51fee8da208c698327f9acb62f9f0de39b54d8d437d24dfd111a068a794bfbf21132308925938e1e05fb080760ad264a239e4fce2b412acfa902cbbab353f794750acc7bd0c4380da9a8e1c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179b0ed17e33ba057f66864dfb5c7231123a16889ebcf1007873e14c8ae8dd9f84a61cd4512b122653629043da0cc88ab3a06b6f0b33986e2b50182d991dabb695d42f52cd27d5d330310170f62cc94bcd7433dc45920d74e3b417;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4b8a838f11009f8e8721785cc2cfbf6b3206f7f65ebe9c397997990b4d59cbf4e47a2f5b05501d30311900763d135945a03b53bc2587eb0f4b43a4bebcc096f87666f694f851fa00950c8bbf64ca7146db30e45d619f034358b5a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16642aa24472a233bcf56d6453a94b2f19db79439a245be0ded81e26a789def8c990042d8b53f64681567a35ba5fdc0ab05f53f2f2bb673f9cc2691d864d9dc9a7d917d1b183a20a6d14be932eba48c8f526da0bc2275570b416e4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13de3011d35138c015b5443909eede55408c51cd9f6f21eeb0e91fc69e79c07069e8055a208b656524175c73d0698e69d3362f3d3987ac3ed0b8bee0cca62b59599399e48c1024a1379eebe44cc93b662fc9aa4dd63c6cb4557f311;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17153cf2a6199b3cf646e51bc7bd3ac933bfcd58ab79ccf063c8c012e2d63e274ca3510e4f05bf72ee2a5d8690970eeb2e14330581cdeaeaf0bd6f3caa5e6c4d853594eede45ea0aa8d6e3baa7e11e6fb1864382210054e73989121;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd00f75cc3a2d4fa9c3bdc01ec51715519ef05abfdced432d73151ef24f51fe0c5431f0db2bd0abea91224bb2930a25f6b4b132805a662778e0af7727e8bd2fd4a0324a7ff94e583fd4a0cf5a9e970436e11612a4d77a41f5e1a918;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10376336a3839618a263b39507cb97b84148f01c74f3c5fede1da1fa484f774e90649119ffec55c10966aa1f2b5f4d8dd59b35dd7bfbc51116ecdf0902ea0ef644521ecf67694a620a1cf154e96f6354feaeb3419c7b9c22c353580;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5720ba0bd42454e8fc210fbc9f4703928389eb3486ac5f3de723fa3d50b280232f8997a20233a1e6c70b1cc8af6c9f6f214758608a4826e57785632e7bcd5fa856ef660e1defb179288b77e307f15ddbe0e55a474e05552146c5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ceb7b9b11986b1f3dca43948dca7195c84820f89ccb36ab658c265378f53ad7a863cd6ef8f97814c422d3e4f195fef49afc21bb44f3b15bcc88524980a06d26a080667951b1a40eba6daf3cf7431ab680d1dfe2510f9628863ebcb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c76107074a1e9a0de2f2223538705331618678b67b0ce633a4e618454b1f5bf13f56adae80c865d9af1e4e578d2ed159245ad971342c3b1b49dec8f6814038c1bbf85cb1b7f478c714406cd6606932925b286a3af687c116af96fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d457f1bb296dc31057ae1d122da95c62f6d7f29c5686644a840664ceca7bfcd7b07da76d5231376b77f01a3db51f3b64b4c928ae4d78e97632cf4a14660edffb02512f2770229b8781deff760baa39feda6f0f4686162502a2f39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26d3df9f42d37e257dc42c0904d32c32aeacdb26ca67a03d2e17f39d55b92cc27d6458bfb187d6443e957c6f4325de87846ad429e9b1f082d63a7c054301d0520afe41b1134d9013fe075e43b1548fa28df859b301f52ff62e2261;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27d95642870a30307c89bc9d0c741f6c62650d5c2abdcf9989ec8d0c564285c6bf516ff5bddb296e39e1554e29b53e8bcd54c4bdac2dd501d59ce1b0785710b99bc1f8d1d5f25512269c94ce6618b1f68527beb63ac14a8f19ebb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ce6d16e4221f58c9bb828dc44dbc5aed21ff60b4940d75da32295f6e6769431a82cc67dd886b61bddbe2eb788453e018fdf45d89b96ca4ae657d35e1ccb24ccb508c3fa6402074254382701dc0af2114ec3fcd87c12131308c678;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee1c920a40301f06810818d467587a5c7a47605aecdfcd13c2b3f28ced5f4756f9f88fc8ab0a12cb8355b102d88d23c70e4ca20114cc100679a3c64ae94e9f27555fa92eb799d331d38aac1398e4e2ff98396188e5a9b534321fe1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1670e335289120baa64d08f30582d65c94a7b766b94fcee9b485cbac12becc453937778eb477559a3ed58ec9fa1955f7bcfdc14c8ceda74217f78cfad39e9b202ea8ea8ccbca5ca64d7ea62e0abe653fadbc82d3012f843e9b136e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126ad44562253585eb2ab08973e82c8a05e4d4e8e572caee2b930bb185edf3777b8953824337098be298d6f41c94008bfb102d2af6d2e21f03c547484f83100cdcf58f4dcac3b8fb49a90cd69097084fb47820307472a710d58c0fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182951e5584d8ef0f5f71b2d720ada26aca1e2da030c3ee3e9a63ad9666813bcc4e992572e672cd5f7b11a84695723696df3da7a32dbabcdaaaf032a351aac8d048d098c8304af20927ee2d0cb9be969e128eceb77e68898289c1ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6598d474dab43fd2eff7a729afbed6f0fc82aa76168dfaaa3e754ef396f52a61108a68189a48c06909d5015f6e8e711923e8647d293b821b4d54efdddc7a7c614d90a58e8b84634a81d557b70827a890381fe010b0ba4960bfbc1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f629c55e673da3ac6734d717f96073addaaef03df0708ce007bc9dd0d3cd8a440410b9ede27448125e46c66f5fe216cbbeca6d968cfe154a2c1956e9b09fac87264dccc68236e825840552b0a0ab98a6f0a405f4f63f44af07fba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7e2db02ff1b63881e0061f0c46557781ae97ed13d4dfa49af766396f39a5cae7821ecee24ff10364424c5225047cd54cbb5c9615d040362e8fe2b1b4f960a0d07e922bf106b5e4ac0060e9f4ac52b634be8024514226acd610512;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111605fbdf8c8e44db7f27df275497f4d0f4024624e27fef88b1b88aead2771726ea8a875dc38c63ee5e05612b27974c6c4218e0dcb54ef0ddec16449be4721d2e1d6f3b4c9eabff5ad32e7118b84392172f1f58dfb37e8ac5dcba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb441c218f6082c2f3cbe699f69b5936bdd77df06e33eacd0a34eb4d84979b2393b249b71f61de77b1143f1b976b45510cfc3dd24b2a7b2b41d09c20cf36f112d28d9b916f237ad796498e68ae55552cda8769b1dfbc235a5e0b1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dcb765c3e7e4d3fdbd6ac19939a58900d8151a6d5fc3313a3b87858a3f6754d4d2ac69b7951cb1c9a5fe78469507a2da16cff76720d5c9cd764742f729a71ae770b47cec95c58e56e2bf9a388bfc24fcc4edd107177af92065b544;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h88c0480c58b56f3cebc659008f38e82b9483b1df98fe30f8209cbe245749c650af090078b83310094f4ad4d8c4c1a86ad0312ac4331cf2d1144bdb1392091fbd35ad780e73fc08be0789f6423363049b3dced920f9fb9740a94e2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11fd8e014d7e6d9605a35fdc5c1b2eb99721280ec4ffaba114b1d2fed17850ec18543e96f57ab60af524b3d679e77fd111ac7502da7db5faa29be3685e319a3ce6fff36a476ba6a474bef5e35ca41e9b73f70b3126b23e14f1932c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97873941dea3a01f1a5baf84e1b444b82350e17cfc2c2db00bcf61e0246986cf7fdf3c373ab2541fb976ddd22ad3dcc5050d0acaf9567ff6079842742ac4ca0a6b3088da70fa037bfe35d0aab1aa3eea9273060248be19fa62c6dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183d64ec5addc745b5374617d7496abf8f39163a0944ae0a684789adbdc058c7a86d97c96e1237f412fe7ebe0d8bea4c623d2eda07a9215c8b6bbfa1bd6000dc580c219ad84f52f622ed917da7279fca530b6f9f6fdb43911382f15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb17a872d3cd426c86194f342cf092ce7929fcfed4c92563fcd4a9569445dc0485cbe6da50bc151b3a05e5ce7ff9a89b1207f5d545ab5b65bd6c1f03a82d27345d367ade8332bd5a848ef2b88ed20cef25d554a3ab811424a60a14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4555119d101482fb05d251c6720a0a2da952c006e7fbacd805150f641440d92c8b376a6130a127311067bd1506b0084bf4e047b4651f3404c8ca8d29d86e99070a8e125935219fafad40866d45cf3419443b63f1156e5cb6d87ded;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a4d95b33d59475d16e3518966b072bafdddc7f852518e627304fd3676ee4f70163dfea983ca9bc485de2d1d16f77cec293e70f1792f9235d0f623911b40708446c34c50ae77fb1c532893aea0965fc2c5def637f40f75c9ae9efaf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2041c4cdf4f7ea64f1d6458e75d3a7bf94ff66d93a0077f250806806b520fda8548fd828a85eb7495190b8b1bcfa6b616f2444246a9e4b50c1f31575057dd791a0d760cb98a28408f0424bd92f0e3a02202a78eb941213114773ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3912fc3d3963b3053ec917a69f50cc9e774f521a591049267a007a478d17c047a753d89bb2ea2e3d2951637a6b60b3320ea2e4032b3e2478bf77390caf3513b8217125e1e229faaab9538b6c77dfa0482ab3f4647ef4fdc3b22384;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haed5ffaf17ea5c9569eda5e4e7ed94d5fc5e5697464485f08fce15d1bdae901ede26e4c3ac366cfd04e17dda1e1f4a2cd528dc25737185e0dd1798446d5dde156f2f2287bfa30291b72505269e2f86783a0d62a0d9f94e5bd0d7f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad5fed756a41ebe8dcc06df88a9be6b0f26dd34f91747e1b15e7fbc3f93b4b65396d0a6dc1ec12a64f3e08832e0a32f6956076d07d0014dc19d4a7f5211ec5d959ce1c1ee594d6a268bdd2acf797bbf64569a4902033884bbca8f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4e318b53d3676752c5231f25d4e03f90a6fac0184ab3e5d87c67ae2c40fe3af2b3507a5a99632617165fe14dafdef903d42d320f25bb397b41d365dd01f59fe54fa8d46b2e2e46064e8be69ed2129ccf59a645cceab031dd45154;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d91dd6f41db31459689a92c86249c1931b247519c34e5ab0e02a90a923d571013825fb4de185e68f59628e5fc6b757d487f590f37adef3b6fe3835337e6b740fd1223f099ac1ddf8620000032d729f0d06a9b9f704d2959560b445;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d94c0d9e73182216ec024428c3a96b0747c869795acec18f87984396e8234dc7966f124e313e40bbb304ca026bb8a6a6ba452f4fd3042fc2aa437e51923f29b5b4b9b9e1672172242370eaeb7d93036600d0e6612c6c7b5a4356e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he19a39971e40a4da6dc5fa20e127f661e935bcd5c72daf68713ba6597e82a164e7f557558651460efb2bc1c954a616605244b9e75f477109979a567081c45bc95268bd52c9d08960b4f3854a2198b004d2ba55546436144404e5de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32949662ab3827d23656bfba970771bd4f20c13100bcd0922a4e939d9625660ec27b5d30c568595c1e14d736b2f5e9de42fe35f54c9bd6d37f03859744d402fc50a0d0288cf7972ba59012e2e6b69a76da72b33cc8d05fee4195b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1890ce483b497f26ffbee4b504d11f4fab2e3a53c33cfa9a964dca048e81206eae088cce37028dd46a9b09c02ab16098c006d8ae2b4cfac39c96e3c609bac1f00b69515c942585c0776e30fc6ae86b29fd3f51d681a4ad232d3475c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1318d887b21f78cc5d410fed9f69b40e16748baeac013075878554ffe98d9b35ac8177374e75674bf431d729a002320dce2ea23b943a79f2fc126afc1ca19228767523e777a5c6ab48ea68cb554afe863c3d8ff9cfe1b1011074ab7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6879949e7ebfa5fbfb914aa3ec32a5115990149ab4844c9a7d7856257532231177eaa4f70fd42017d4cd9a9f450112ba5adc59f0992f691db3a4cb17dbcfe2e4fafb5d9f7ec672ea97174439f6fda4380a57a3d05cd279e9e04256;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e4113f9debd7c41c0300f013bdd4575d2d9ea2082fb0c813edcdf43b3864f79f895deb123d9d0a8b58aa2f954243d883f798926498ae5c25282fffe25a991517628bb3ff2e74332121268717699a6b8dd8efae156080a7ae84766;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34c355899d01d9bce907b25ce8ea84dea28c032f8e48bf0dd844548fdeb27ed22d5c981bb156c22d4319950d41a850f4f04cfc2458ce91194baf4b25e42cfb9cbd46cf30a82fe0c8d9c19166bf78704541aa51f0e4476fed1a954e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0c89da73ebc3a3cb659cbdd4fd84e2f091be9d91a027a683b23b87ee56a960ccf9d345891107a17ed5b3481628f12448f04f56c23a45611ff1a5b431242010ded43d57200272e35550715755beb1a3dfa67c7b72d7ed0cae8ef45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6916da7678f8adac996162ea89277bec1bca99ce7a62b1a2259803ca91e53fd7395d4d7b87dbb7c4ee7ad9bafe903034ef995c6ce19e57dc8346d4dba2010d0cace8ab964f88706e295960d2cc9da249c54ed03a4bb061f77edad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7559bb0cd0161436a512326ea7bd42c335b4be30cbdab192ecd4fd3e76aadc4714d447fb9fbd8913e5b0bdbb1d2071f8e8986b58f0448eed21a8c0f67bbd120995ec83d38d84bd539d8639fd2f9ae33184e0caa5267b068c29a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ab75dd52efa1a63134105ee8dcde5ad2551f34250a27ced498d83d0cfd17d58c3567491230b467d72ddf20b3ad7937f92922e2f27e113eac06275a019706237a46eb45bfb76ceca3f62a8aa7c1967ff4a1f485144006a134d894f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fdeea330d1fc4e814b8f21c9aecac28f302f180a07861809b6733b171ad1dc6ccd1d150eae6c210c76059c1afe74611b75d9e268faf15853ae93060a58e41dab83c30c88bd406001f8b0b0ea221713ef093ba10af17120ad31524;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6ed2a793853317fa7cf79b1eb406a444ff88b7b7cfc9598336cb6eecb65867881c8c8f3d2b3075432540826a1162ce2e097b946f61cb17b2043a5da8e1929b21fc4df808384f024d53c0f1f97c7baefa147a4c443c751b407b4b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17884d87a29a231d17cf6afb700ea17ec4ce67d9221e70ffb7fe5fcbf9654821b1edf4db7d1873b9a71d125af62884ca496293584bcf7bc530694858914360152c45c183ea44386466c880970180ad1c2f4b150b5b55b2e4667db5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf8c4a1f404f5b055fdd02667503295f4380b31414dd1627fa9badaf46a913e9b323b0661a755258bbe26773c7e9954bcf4b2dc203680b0c39ca978a6caa5e242001c5317efa485da34af1cedd8e40bb967f91c456a269b18f9f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1feac157efc4c8b18930e55df1e0dbda2482a1af45ceaf787e665684156ebcb950dbda30e48b9c359a4789a0b9c62b8c5c65febeb3d2dc641a817105ff82dc57000eb46914c3a1589b29955c42ad0a2a584ebbeb6d5719bc77d1a4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38fe88bb53dc07ca151315f8a651e5c0bdee32129fa9ee395fdd2789c027b72b7c189621b3f3df4c75dbc1d3f3f3f3b0cf19597d13248aa09616d307db9fe65b24f8e7f3d6dea84a60c977bd7c8fbdc87e783294d9d466037212d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16958207f93e7df7ff48889437f559f0f34a2bfe5f263dcc5584baf8b5b025b8991e7365326d04d37138b407621336375c89b64d7a97297a750f8657d8d729676f8fee1b2460e6ac84380055e8fd51e55dffbee98693a1aa45e9ac8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e415fba32976f3c6be2cc0d12e929f2124ac50a66e24b1edce3f30eda4c35c9f82f516e2fa7974f3383617f2b121b54f92318c59df3c97c4c3f7f5b26d6a93c54a9724bf61a15236fb57fe83965a1a4334a9902c63d5c48a73970;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a983a0960a02a3ce867d3ff1f9299c408418e95edd184082726112d694fa0c4b091c13ff8786641861ef7879e54cfce70a7a6883b6794819184038c68240fa007976c6eb6f2fb22ea41515abfe604c61fc52237df710a1098557b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111e4f06b8ab79a25fd36999318cf3463e8878a2da4f06ea244f6c89d437f072c139e87bf6d882b936b8ab1eeb0f27e6eab72e1d6132b7c851b680587792003ca6a5119838db922d1c7c24d3d4344475fad99e943a183974df5b6a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b807d7bf04412d683cdf221272976664369361ac92f63d374988532429cb5bbc8688c9077cc901536ed1d8ecaf86938db80ea823d50106c4791e9275ce3981e8a125a82bab35726c1ded6f58605b050293465af53a7b7dda7f144b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d56c41a799ca62e79e053a9ac6e5fb9d7bca56da517619337edaf8d7d9fbed3d6381f5df533d8d6ac2167a479e3c94cedd0739a09e387a6d5575a850f74f2bc8a4bf023615d6e9fab9bef7e674f3e91a75d4568c5d17092f2da26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d50416f3b12d1a26f23a5f9aa32b1a3316aeaacba8e9ccb3152d35c14da47426d960f1f3b57f59627bc922f96cf9ddd43c094cb6947b74dd03dec884b53be0e995b84c4023281ddfbb35c96745f693086f2f62a0950501c406f9bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13711c73484c294e452822233496e81bc6eaef5d7c5a9abf0576cceec4c35498ae3b4b5e11db00286efd775e75a9a5cb6d854b8c98a34b4b6c681ecd0cff47a062e8fabd6834ce95afd47996352ff5a95d68f448a0a4ce6b8ae28e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf465bd020af18dc9b662eca76ca00ed9d6c188c08f5df5a767afc862aeb06fba09b828685d17310a9c8305aafb09d6915e494039285bc08aca0e3d3df7a803bda0cb72c73102bb76ea3b176a106ea4a2f723659db95671ecb2e300;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8ad970cc04458d47e6feda694f149edd33ab0a1c5084f546eeed8c3d8ca13a46a62c7da6b880f63e3c94d3eb69e3cbc640698f4f901c24f054a131989bf94f0d5a586e879231a0ada36de28f50b1c45fdf3a29c186c0a57b4cfc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11032fa36a933df4922221952a2f787df8e9de20b5109a03e0d7d512e741e2a3a14d903fb1a64ea4740c0d1a311e0201dea93852c8c7f104deddaa681ad55ef31986b5cf603e02dd7d562e7ba7d7080242b212aaf78ca89ddf3415;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11699f1640b4d78bc7a4941e336be067aecada98d5cab5a79712725a4c075a82c94f3331737ad6dd7e3b12f8191ddb612d8fe07ed08f7894f16032fa1e0e525a0978bb5fe284c685068198b95e83eda68f7cebc4298bd595bbc6d5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea1400bbfbba253cfa2e822460b606afe5de0e99080275a3c43a0b93ad18abd8c4ab6e0af8f694ff07056a82adabcb94b9339515f608980b7704972f3d8b4c8fdbaa4535e5fa3a8707539cf6d166360ff3514ee7b4a9d3cc0983f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bbaa378734a78e0a71f2f5362414f8a08510d0dacf041a6dc773bef207f022b3c704fb69fd8a63a7d7d82603551cef220ddc3b5ed05c6a7715ff1b19004bd2b956ddcd54f86fc6a69557d42a72d693a3ebde381a83ca52f5df77a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17b3a07354fdf73899266b0e30c09a8fcf476b0af4a91e3291cc1ed2055803a82d918280d0856a58cac9a3643727f49a3f8adf89ab784b148ff82899b5a96298fcae6cb3486e19ca8711c81ae29e3d25000c81a38c33d70ed8ae59c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6397438a23b5298384c4bb21418fb7286e0d35cb35a0b77bc9d3bd0c5e6af547bd3ff4cfc0d9367b7e1f14bc04fcb4215475b44e498779fabcbe0982cbf9ee23792188481567a34a2f58067ede05564e47cd6bd32491b48d15515;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17dc7f908c21bec6f6ec0bb80960bc7c8054d7803498aeeb94db0c28c6a03c1a61dd86d6e288b73fea02d6faf93d14ce469a59358585a44f62b5df15f47966d847ae6d9a3488c7cfe437bc49265de967767f61f77c8fe104feb684a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb09b6f2e34e12c17010b925c94c472a0ba9f5f2e2eb4076ea0843938ab4d059dcb02bf6dae44b4b385860c95b309c32253c5146dd1208f9e48010ef906d32b27ad2e33674f139506520a780cec60cab9190bcbe3db3ac605f9ef52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe74a98f1417c51687c3422de6938e011fd1add4ff23d7801ea6e41e791deaab294a57e6236b7d94e34b94a7d0772cfa104bf76669e482ae071254a459f9b0edf8d28e390b14656243a0cd43a8ec919e1086695bd1d95fdeaa4f3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha28aade7730afd1281b2636cf6c58fafa2d4e9bf650f3f8d8662a49e46b416d2b1fe4e47c3d6d2564dc93c06054f2886e4ac37713f04295956f9d926c74135b6c558d02f9d7381d326b5518d4257a64b7fba3069ac9d71ac5a2f40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cff8f7f3a559864a81556ab330cb473be23c3a077f9bda078cccf1b3588868af759e045d4795e6656c25a7ac524740de84cba3c55f0302f5d05775ec9f734f5a544a9dcb885286f8be3e99c06070f4ce311e7a5c5cfd5e121d4809;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1298be38e627e7cd814af1b8db115673327c8c4eca8a90fc3e82b17daf5346bbaa32acd25f571945ba26f227a7620b466325d26e819baa1c9e567284f85399b6ecbeb49702223e793c32635a81534fcc45cde4109f422f5c571bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bcfe36ce7c7fd0de5db7b7a448fdd828cf4700920d47e8c51e6e6402fb3eed1db6942306a34c89134c91baa4a941030c0256f4094530b8e00906bb091531d6173f857029a1dfe57c6b58b8bb61426579b054405b5d5184cabb716f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7216a88dc9b55e7b6ddf6326067298e1bd6d17d6f21d1279108ec8dc1a9a220637b2d3547139bd16ff44d2dbdd528a1783150e5292a481f2855b031035796f75d9951a064db7b7f9fc68ddc201c0c1f9fdbcab8c84d9a0907fdcaa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1915210efa9e4292a3a2faf94ec6ef638e508e5a1c2c5da877411491f395f13639b78dcde653ea5017e144572e189e8642f98c59293388a2226ce397b76183218ae476a6bc3ed7433d2c1a987721122a35261022a137a473e2c9dc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1b9484b02765124f8093a424533953eaa51154a314a433204c036cbb070805f4c4e97deed7716fa32120abb51c1b92c123c2c373de1832f3c4fa811820dffb629b0c1ab969e169386319eed5d7382ea25a7dc40a079e40f068fb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195f711bb09cb2529bd6d892f2f23d582295de79080c51a9648472770a330b4c88135ac3c4d51c4c32a0502a8b3fb0f246de3072545e098422ef9be952b4360febf4c60ec037894e85cad981b3d0b90abe62d223445121ceaa16d15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h252e293214feea45f2373b40548bc0c629118e750307def792c46c75d5c5d884c494145c0c71ee150478c3c3a194adc26c221a3c368c653771e0726bb4f93c89562abacbc0d395a728e49a0da217238497bd4de87ba8778232db95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b8a7857cbe8cc81556f10b2ad75811220e8e462725473287af0adf71583e9c2f67f91782fd63c7503283582afa6c22d1b65ab17c24c5af1aa5100bf1e951edf9e515a12237a2fb389a10f61f44b60afc135adb632ed5598e17edc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bad9f518943e521bd6cfbabdf9c7b1a94279f9169a320d74d105526195e9a0d2033aa3fb281829648ab542ffa2640080e9df3db987f5539acfe0097513b4fd2387ab28cae8d3f23a180b59eabb9d4934972b2a4570e2a2cd5d9766;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db8be64d660b6123aa8feb9ab1ad2cbb6d89baf7de4ad933d5ddd91cadb4547b84ca3bcb81c90e26e7c56e82a59d409fe8b54d5c27edf0f6a28ac1174cfb080513213c8114df86dd69a6033cfb9a746a1d6446a180ce1f78a7650e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10aefb102f5bedeecec718d2bb71a9ec1caad9948a59dd10623835d8d179dc7beb4a9bf2efd1e7944d9a576854f9d60de48b364df00bb3d7f9ff6cb1cf83a7bc8520047216ba0cc29d145d1a072397c973842d7de6d920d4c75cdf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e6c0fec574aff965edee15e6168cfc03217372be3729ce2c3c3c54500bb27e4f1b0f05a4cc81dd6e7f6b294a3efe5a4940ba5a631dc9681b6a7d1226a0151d35d2b5206cb580f6b0739ac45e46422ee75cf1a3eba72652adda87a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6e3a9582c3bb6423d8d63a33c0fb4396154ad5312123c70f69f571a4998cfb71697ad874714c7f2fa047dab55a48668e31d3a4600882014bbe22325ed1f3c5dd6fa2bbd6a77076cafaf0b7745bb9961809b4aadcf5a8dbf745718;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1056929a39aab848958fde70b838b3ab7dda64febb0e2ead8f2bdbe670753adb6df6619f5758e2bc12180c8ce5584543159c565a8e701f113ef13eb870c918e3001c38b0a21cbc3ad914c9a8d569cdee309e0704bf231f5a60e7f8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb55b0077481110bd8ed8c3b4bd031beb47c73d1fc8c706a5f537ef089ab8c51fdf428df7d15de3e5a1811a5ea49f577e4b96777b551a12eaeccf5dca18a5d2455ce47055917b671234067da95494a6a1b646b5aa07b7bd8dfcb0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha19c585facc9343544f16f59cc8c19935ac20d5af5f0a64ae2d8a3dcffb8041f9951e040e4c9a13a9e3f5f00492f1c7f0b0ef1cc43439beef780a57a8395f8ad20dd091ea6a24e069d12f1d7f68755e27bd699a74df0aee65c6337;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d016c9a37b9786a321e3ca5b3641b60529e2a397f7138d7545d479490e1d8d777cb8d6fb818db3f076174b6484e95b1a52e5d0d69ab99ace9b0d536f7c94cbe26623879e4ef028402c4bb54e4ab4fe26b65e3ec721370748edf583;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c47ba2b150bce62b6a389fdab212dc9805a62dd60b046380c26a008141615fa626fdbe81a68abe68d55bdc0fe6a8a239322777a91b6ac0c8505856943719cde979681d92753fa81aef2c7e57e2a96dd4626c969063ebea1fd374c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed45078fe80e47a56380693d95408bd0c80925999f7023c05d3ede63054ac6a2413b5882f5ce92122944e2768291bfaaf0d679dfe0b14feaaf0c018e19df2e85865361bd5cd66e9de43636e3f2c9430b7b3b251d4dda1cd9c2ffc1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153c6febc1c471f39e2049494ae17f9c4500ca4b391cb63483ee677720deb648f52cc11d9eee646188e1fdb84e558f8c5354c81019824a0f93b37eab756a25f716695a7b97e88651a290d2db472a771815493e7f86fedb10881e8ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haead7ca469facc2674bd8372de6f142c06ed1842723c35f16a2315e182e0df0816541a323a35f8c8d701009baa338c38ac7d0166b89681c6de4af0afe97be88cc1c11b9495946472562c05e9b78c6c9183b86e53a121d9678c778b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1c599505ec535a53f3551bbf7107c7a98d4e7df9974eca9ff8112c5a97692676b503ca9fe5ecd0b72eb375e7e1afa9fccb5db5518efb25f7518ef743825737d869116a03f56298552ead84aabbf0eb91280455b055123f4483ef2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ecd7ea78f32e7a03f10c2c71e4949eddfd22e4b8e39a77ebac39ed016e0b130d7f091652c2c05ee68bad6277c8b0ad35982dd476095059386a4580ad5c7e0781fa97ba13083914910b44c9badc542c8f1879792e2c41f3781202a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69a501e1c548df02271a33b3429064e391d4ebc9f7503a0a9de880bd9d1a82d754bbc238a243c444097c369abc7840bf7854d81bc3a382e372ead41d16aa7e34e016c2de859028c0adcfa9c6b36131c2a5a12c718029054d580725;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1754bbd8f9ab925d0336d649455b8795550235476d73e0ae0f48919f266dd9c1d7c95ad9c1080c4667fb40354ab4df0f9cb805c6e6d26242cafceb1bda031de1cef993ae8413dfcaf04f3ca0d45008943d148db0f43298a9d0bf23f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112007ee0d44a62874c0778be10f2ddb22f605aac29c6de0b6efbaf63916e43363c733993e525607e31c3a835f31f1afba58ae9d4851c2f0953833ef4f5c0ed336a358c1130b09516623161d874cb5348bfdd76944cf18f7e67b40f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122efee14c7542a97cdc2d2c817ef2a43fb8f32783a8cc4fbf1e3f5263881e6b05d71068a49930e04d0a5308bdcdf560f29d1851c95ac3e7907694fa7b6e6c676a13a8c4795bc15ce8ba9b4d52559e696e6ceb6bc4dbd451c8ab13f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181336c37e9fb570145c5bd4c548da57e6b2ca7c9e224db4c8abfd32250617be19cf5cf56124a81a4bfce79cbf066bdadd34b460d9d9d2f262fea3c3e4fcebf98b5a76d79bbc657463dce8a4dd9ca6d472877d23698d0deae58ddb5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5f6ef01682a1dba0290e720e2f932fbe35cd8c8a2031c86dcd5877d9369cf1f5cf333405bfd2814cbb8acc60d4d1ef660c7f4091a6b4e9353d1616d953c759327f91be34b889b4cac358c1e53136df0eca6a3d261c623c99fcd58;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76d977f7a027f4bf745e3154cbb9e0ddc18ba22fab3e7717fc29366360fe95f16052beffdef37003b323414146ba9637c107934ba6c53e13a0792855dda25626347eef7267d8fc4ebeb78116eadb3f9304ae6a4fa42262007890f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d7096a29e52214b438ff016485510c70757b625b9271879ce46f4e5febe3fb3849014176f503107c1973a4122e0d5f3b2ad032b1804a0176a3f60315f0109823f9ae71a09f066308161e9a85e0376add89e878b3edada746007f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1758aaea7c8a8db18811f52b8d58a64edc899fbf0191c015069a2b687204443e5dc8851ad211d705cf2108a53a9b41bd9f3f4cd59f54b95ccccca8261cc32b242b2c13a30aa70c512620e3abb9fbbc8f4a851aa7691a0ca5bd811ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfd513f3f9265e70e0982ca708ec9474441713c0d6c32c4471c8e500d0a0d522033da4c5a25ed6de63a8407907242b72b7fe993c695a8323962c1f79e50bf6dcd3e917a126ba22c764819f58882f2f40c66014169fbbd7866a7332;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h60c79b54b55dbfcd85492d272eb09a4ecb71834b34170c594eb2a9dde9bf8639ad77ec2f423a4426c2ac8aa1b0df484f142f856daea2de39c91ccce3894cd29b09c9d1967b230c845ec2ed0812983e8d585ec8f01ffe71e1766b7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb43886fd16c335ad58adb46a480e66a7940a7da39850549dabe025d405c4dc316664d2cbcc3633157905172e14f479a672eef272eec170f0c1f8decbfa949cce4ed2ece3c0fc7c8e89c1f664c0a74a3c16f15b86eec8a200bb247;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141576ac022bb547e1ac8003fac94a04fffd3445331a9755dd1b1533c0ae0d8767bdcc8d00338b1429d482e4f1674c9e3f10905224873f07002934ae2e5e3f21b5ba46fd1b3c572894934142673c8d89da5825630e00dc9a65133c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc43bdaee9f218f305adcbbb2f18e6edd311d4b940888a6d6844a76eb850c1aafe7ff243775e842a1263cd772f383cd941a8a1437c573871ea97e8e0a1ebd9f29626bf80d38d4f651712453fbe9ccfde8e1bcaa15bf2bac40140684;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e02a3e0ff913c9eda87a2eb6992d66c2a781543879e40d3c1f99c795f028cf3b5e3c1ed42481227813d5ccd80463ede5e93306468a7bc8f3b635f02e48157b0d4a8237f5084fc28de68f864aec930f33ad7553f094520f4f1985a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9eca55a7bc92fc8a034acb7f4a4b0c11c4f7819c9fdbdbf9c8f497a84bd853a6015644849fd545eeceeb7bbc15bfbedfb5f182eb1dafc97f1be52282dbb24a1e32a5a1e6910647588fb3d1080315c297b262ba3bd214e0e5a47da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hecbd2abcc6ba18ddb7dbea9f07115a705f251502788a2c969bfc1f4feb9f7922a2336c64645d9c0410bc19066c1b8623a353e5f1cdafbb6b49be01b0a7f35779272297212e8eecb8e1a39953ab687833aeb60f87accf2a79f41c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda5ff04f30f94dd0e3dc1a1eb9c916f3ee0ae53123d63cffa781efc4b4fccb9871e7bc4a0a9078001cdb32e24fabed27c48cea720b8c30a41585b49f6e8285a7430d7337e918c28129944c629dc805ec30f85054941f3f5bf6a359;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f62c9f91e81f7ccf283aec50e58936fa32d9abd81e2433aada87334a020f5a42d0181fc39e80219f57376c6c6e4f05580da39268841c1ecf2dec276257972b35d1cb3352610dc386cb8f9693979ad6614d17ce709cfcd8e093fd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0d9d944aa745f5c8b379582cacdee88fa0c71593e55044fd297b8fcc29ed53b57a6dd13bc16b134f0d706335e8a449fca44c939c593c2889b5df757963a07b0557b83bb94083e42b55f9ac5433e9a60afc4c3d61285346773a754;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0ed2fcfd0312fd32fdadd2e009972ee0de4e4a458ca3fec20ef5d3a3997485f578cd2e4d1533b3b0c0ac2b96b33482a74df8f8f316442fe57ab054f8a83f7c26113c5aed15dadb8d99514b18e95dd5c6b12cd8cf187ccb47ae536;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13fe5c27586bea3c261a2877a558b852c1513d2be03b5a769a1108a6e7aba9cbfa79bc644776323c646c426f336fed0547aa77c32d0d2a19d446c2d47fd661ac65759bf61bcc2c02a18b99886f757602b1178300388b7cabf31e3ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haef72e2b156e5a3356a9446eab9624543dfb0c861817ba0f960f5383345b9d83604196d75dbe44b5583c82021802c392da949aa1364efe6fe5953aaa2ad381ea8e28608edc492a2e4963f3555043e618dc00b0a02a74f8db4ae363;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa1f9e34d980e91b53f42a0973894b467dd6093ee771546a7874fa8181ec281de4250ffdf5e8bca37224808af062e6856999170542a178fff2c84fa3aa8f32efee0f0e3e77c994330073b21a02fbb6e20bcffef76a3618543eef51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a54aaf9228fa6da7e0a8f68d4601ba8092836c1d7ce5a16466671cb4c6115e05e193fc9aafa96a681f56a78411ce3870e9f1a2223785c0fa31c8557ae6a6e8f1fc2ac99bd2f7c305928a884a0a8d8d10ec5611c3f9eb3bb27d396a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dee0cfeef0c89b25574f63838c0e650a5cf61dbaca0ba7dcba80f31851900933810ec18637a623a15c9c316da8e147c8632ffa204badaa5e445d52cd032774e558da2e4a2a720e276342d8c461b13d6498e8d1b62572d84105f36b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27f80d5590d44f6a656f3dbcfe753e0999424345855e6c5ec1feddd1f282187f369f38f10280d7e882c1e61bd23d7e8d2cf7831fbbe051860d1a2ddbe57b65e6b41d93d08068ec0b27b9449632dc2a14e732417b9cd2a5dbbdad9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0c5ee5fcf6ab8439181bfe4e96998a475de03a8272262b1a5f731e110484b653e5b038cad6722cbd25ae78e040277b0c1d67d3999ac23162b5da17fc0b5d13eabf5eaeef61ad2f9b02f689140bfb79b4cdfd73cd1f5a2feecd7de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136f650c01448660178c3faeabffc99486aaa92549d2639cc63423df075f6568648e12948b2cfd9e750e02de47a08faf16b4a5ade18166d691845d7b03be11967224cf56eac4be0aceefd3894db2d8d6a25b1c24067ce2f5629a8bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3717a8e7791dd9e273ea4b26890ffaec27ffa2feba60a61effb632429e4b1bfbbf55cc2a056a58375d66b2dd40375fca16335a9bd18a047411757e544e87594fb455695b5d0929292d7b3bb1577d2e0fa99a2c409c803ad2a1083f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7732c51051f2933e6ce158ceb0216e956a667c5a8a11627cc9fea412bdbbe700838685d3f532495b59da6a5d106966d6f63605ba67612dba3fa6ea61ddae0a2f8accb071183e4c7ab35f678908460aa1431cc78e6857523923f7fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70bd26ec223c448ba5a395ace247240cd11e7a0f0d69d1b7d8f337d6e750b36e5955aa888b43313be14835eb0dfc253ffa63bf9605449f00109f2e1be1c219c19032d8e7f3e3b09ce0e8988d33c119c1d85e249bb2e5c6b40541ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e514a1ed50c7303121bfc71651d29cdb761416c937d6f2d24ae244767333d62b2fa113c1a909916e85c1b63c1849f2834edaa9f12e41679e1e4c7a808661110c4755e5a0f1195335440c8e46e78d5f23b9d782f5beaa5d2a4d1db8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bc5540a54f7c2db052d4662fee1d12b28e62b7399f1596b07751fe7e34857e2adddd2d01ed0b6ea3d7b083e7c47459bbf4a09202b533db4a0bb87c0df816f451d5a15a36c516d59db0ebb4d4d8f80031559604d4c06f99e030328;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb2fa0a040225fc7f88dbc4dc75c07aeca504f639f47bc759c381a935136cad670dc689e65d7662bef25f57948e84eed33e3fa013a5c62e5a353e60583f608732ae8203560325e173526bfd15fbd54f71eac1b0724166af09c22d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c8a8fd3cb54715bce300e94f6aaf69ce33f6e465ff9e7a7549b73f02f30f4f167e233a85133475c1429b611bd0c92c317dac0e27d4af2583ea96c6796a9ca027f98de72f2ebd3faec066389cf28a453bc4e794d19fd82eafb2b29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e394ecc1d9e3e94154c5041ce25747d8ccfc2c23f3af378bf845fadda1b6dd7b4bf9140542d4556a031ab193cbb891fcec5ee901ae52bc8d881ae11b0b51c346a9099c837e947c24d81a018f97aa05555e4d1985263bacd89b1c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85acf4e6587beb85bb39c1232b5fb33c80824fabe216e78b2537df4c6d4fdbeb04a7dad8ab22e258368847363754bf363482d6640ee7cdfd281d42219efb6af10bc84d6100b63527aecf6803f4ec39797ca807eba4d5a90ac49f38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d282f8976fe11df434d91d1354b7dc6697b13e78c6ad89203d7d40021917d1ede15702cf707aa92271c3ce3ede98056145fac1aad64b0cda89f9ebf12cc6cd7076ba67048314698d949bce5f887db05e088441fbc6a6d1ff23d1a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac0459b4301d799e31e7661a5cf829732fe00e6ff6b7b6e08954125b567bc85ef9ae97af4cf40e3ab1a6fef14fc4a36a4e93b32d16be5074a37e2f44e5d6e6d1fa64e7c75d374b742cbea1c22731fee2d6930756fb06115caafc6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed6bdf09a2689bb525985e74252a13e1fc06cd23953fc52b8df4ec0ace5afece531f0e12b8313e6b86336046b4d77ccd49251eff3d6c6c7ae9646e7f348aaf568f1c7031de317f25145d6f7d824e5609611b4ba136fc3563812269;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18dfa01fc46fa6e0d51eab5fceb28d308b00e4a0a90e8d7bcf890d3f22a73d192e709496bbc107bd4f320ecd105df00f586a0e74651873ee1c508e502b583df78ac25c4b9d58525020b8d2f3fc79a32f33053987d1219e37708189b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15491c152a6f953d442cee43a1615ffe0ef166fe8946b3a61ade400b29e25ee3a183888b657c0869c0e19135e2a3232c6cda7edf901a0ce6ffe8aa84cf3607f28a91511fbf956e002b611880cb66ef1b73931e5a44767d7b056152f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6663c6ff05137a49f5b06f837d6adbc3a270942b460cc44c8f0f22ab2f8acd559e2515b462590d29b155a85c851158e3b7f457e436d1b8ecfe65fd6466eebdce157a4b1b0f989b5125f18df787b4eb5d8f0c1a69d1aba52e75f66a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ae2394441269584523a605332500a3e20e699d306377aa89f384f295a2a3682a03cebf9cf6206d2603e4f9dc9ee317bb2f6515450d20f131128e9d6208a1276191c8de99953924264a1e968312f0a7353e5918c95e2e7cbe41180;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15faa6811170b77aaa0db9986eeedb5f1d774737e3a1f3c2d489ff5bc37cc40b042ce29cc833bedcb754a316646e79bc6e6c87835aad19416692d1dc215a5f04de6d15cbced5ed83b67217a91a6df426d28d08d3c3cf28b1619e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b28950845aab1562d4914ebe0f2d7e78502bd219aa28defad9f40e7dab579b7107cd93f4e9ce39af3cc071175fc85db18a18616b261fd5c147433a85b603bb9e647fb4a86e2ccd27d68e9977f4c634ecb2375b3738fb3ca057ef70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1734f7f5b02b1682a737c58334944407c095a22a4d42274e746bde667e55a750d4b9d0065778e5d561cfb617be450eee4d7b1280f67ab28532b4e620576edc02dab01c0e77cf600933301930eef96c8d073d87fc85ae4475a424fb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149db6206eeec8172342a6a76a7d2c929741229e6eb4f26aabf5f93d38f2b41f4a15dde3824a0368609184119c035b2b3a416025a245369c47ccf4d13ee983323cb0ae63ab3b69053c588bc5adeb5222f9933e5de4057c4ea34161c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d8caca91c207bfa9754e877772fc3559edbe3fc2452fe99a9de0fc9fa824815f1fb9e745577653b5700907a749defe7086c55107c4a5b1f4822b9db3684c311e5fc05073e7fa906a8b37fefe12d84617809b18138a04b4c476b79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197ccb62f62dd067f07edd803297f315ab251fad93d63cd227bbbede9c1fe41ddf5f21685f97f61d07ac03cf597a150b72256cc97cd8bba7edbffdc2722e30210873e1f1b19ba40f9918935139ec38e849e50919e11502d6f18dd26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1084d3061b6ec2a946cdd092d761731452bebe84ba083bf0ae9b52cc4264bf711771cea124cacc79786293eae0735291841e6a1bedf695ca0f7ff2639f283ca52fe71c662b8b543200e780c47af6a38b22249fb311f7d32e19ea27d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4e22ab63087163c43e78939f813c381458a36d1d8e131802561e3e58ebfb6fc52c5cff7298b8ceb6c37b95d38a9cf3c2fd6f692f778a2d3d412deb5ad508d4f3dae8dedad35b0ded56a160289d0e022caf83e45030870ada371c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc2ea6f2b5920c218f7af7bae5062eae6bd54ea0842fd9c2d0226c179382fc897f517ef7d1cce009f8abf31efa51ac2c22c3103374121835127cc321be901c24cd1c37e2a208e48c9859fbdefe121d16cab998b80526e5505b8d1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164112cefa4f075036ac543c0292b697612e518cfcf9f9fb83f7dbe47f95eb33ca0036bb061e0afaf9b1294319c919dc74345aa3d15ec1e4b529317bd71489ba37b03a7f1365008253c8d230ef20aab3bd1b8df967d5dd92a3e6c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2798670847aab56d0f3b333fa9e69965b1cd97ccec9159603f4d959869431f4bd2fecaf1e7b3344cc0ec6989173db6a4991e752da5171dd742b3c282652b8ad6a65978135444a5144f8a1d5fca99b2524322bb627df11ae09869ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb48687af763e75900f2d51c8047d79bb68674ed8518da0710b8abb762f0ac9b6d8259d60bc560ef342f46136fdf6bb9effb95e81a115b2b37dc2e20a0665d63ab54511f5a5524fb1f80ef212dc1585133d5a50ad577f2d1cbfc637;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb4db0205dfb63888dc54994245cd041108776ef042c6c604e1983df884ea37b6a186a5dddc41d132cc1eaddff1ad358967aa219d8906cbb27ce4666e4353c9c76e91a8c239afa3d28d0f8382cdddff1f3ee5d733404b81052eebf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7eb7cec70e0d4b1f1a7e96b2b28975092ae3c64fc6a834f1ce72d217bd86655dd09903d36d063c3b766fa1c280f082a3c698dbe00ed4420f90d7eda74a86860861236de0953373e94f26edbd1dd884422db316c94fc134827903c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104a3e54c6fb2d3285bfcf1459684bb169d579a605bc5d2da0502ab01014969c20d89a8168916e491d1ace0c8eededffeb8c8488a68384a4f2be56be1e4edc7ef999d0244dd21d82268c9cdf99358428be517092a9d967bd8aa815a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152b707df0a363ad2a31f20173166b8db302a60d7c625fc02487dd76407e41fd3e2e43d0076d8dee268944af472eb4e08cae219b8400cdcb6adb9e678b8deeed2d8811fbe99038bce5fd7cc5c18b12155e161ed317ec4c3cd7eb678;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h66235b4c4a619edee7cc2841f124b682bcc2990f3aedcdcca624e3aa0519cad4a897f61b9bf97e0008c7bc4a7d950dc0fc15b7c9b851f2490ab805f39ea651cde72c8ccd001cbed490eeb2ad17909a200ea064fccc1c177a5ae139;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d13ca85e6a94b82d05796156c20df44c686ab79b9156bea6f4b054b46c8c4bb9683dc290a45b8b12fb6810b6dbf98eed31c321268599d77e8d982d2f20044e2126b522ccb0c8a19d7c9b1da83e89ee182eb072e224b2b90adcde2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18eb42fc1faf92b5de097a1368775076c96b5c59e2a58dffc3be4801f5073f4090de654a79b8873b787bf5ee09a89e0b9a9ffae660e047bbb2e486d9a559d6d69af016179fea8757d24c677b87987ecb78ef9662156537a01aec586;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7af29a828f74d6e36188e0bc6b435e0b20057faba07675bb482db0d8557094c4dd6f80a5d38a04ec718a3abfb2db768c71982ef553bc964a53703c8b2b14c209fa3188a92d76b69dfb11f9ab54efc37f4f986267c556bfb36985f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e641527dc3627d5a77ec0b0b29aec6f18a8cc365cb1b26916bbb0a613264c1e6c4b3a099765afd5133f6d63ac01165c8d3d74d5b532f5e6971d1914746307b00f65ad6f7a66816f66affb30999650248f159817d4cad59e436c181;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170368908a822fd2e16748bc9d50441c0654a5d35e39651e19e41ef5e38dd13cfd978582276c7f7f8f45ff6c20a1cbd1c2f4105051c620032f27f05ae542f97d1e0a2f09ef63b9b46718013bdb86f1d3299fd1960c2c7e74eabcd59;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eb90f2ea2d855d7c86bd3742cdf31c5cb5acedbe462c95d64913d2ba565562a3b22226f143aa8552989783fc9c9c2ba10855b04b96efbf6875485fe9f6bc234bc640b9852a5bae3b581f8fb4f70fa91203f8cd95cf723663fc68b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94f4a852f11781f8e3ee4b1d0dccb298a7599935a5a0d2af0676a67d4937c706ceb181c1afade8231a5f7a268bf5f82821ce457cb51fe0f31ee03dd1db571ad6a8b027943677eb3f7acc2ef27f36bb9f328ce58cf38ee1525a62e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149ce24364bc736bf8bf52c19a54caf2dbabe302eb5fb03fa53cac0e984c538d74e2b50dd59bc087176730d680fa9181d7231a52d06e172d295972d1c0b29a26c84bb41b1679270077d63b26023f6ac704d962d4acd39d85bc5b902;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd39235d11b3a05ad73fae070f9b6d88dd633f13dfba1d9a46bc1c67f5bfb80619fcd80977b5b5c83b364d96e857f715c429ea17eb0f7b15d1a36041834dc6a6dcd1ecebf7ce53e4c341f997087f4355d1aec069450ed261bebbc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d6ef98bcaefe225c272b6160d40ad74da648055ac549c09047c58ef5a92b522e29c06cf1135e0ded6c4a54e7da9fb038103353beaaca16a5dae6488c348c5b216fcc26fc1714d7dcf2125538679b93a61dea867499fdabe413635;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1328e80fdcfb246393e72e8ed8a61c9c38619a2c8385c4d85b8642cc00074059659cdf112a6ceeedb1f307cf7e8ff7b690d40e08cb2cc2d58e89e38310dd65c0c2e7d177b20fe6153c8d8b8588d65c04ca587916b2a8883fb980402;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha31ffb434961f098a76c5944303e5b5ccabd03c8a0139f3a805b3015d6ba8409fc6833e6261a5be4c7928ca9ff9b4af1704febd96a47e202bdd7a476c5d392c8963be92bcc506e733842a2a65e10094d45e222d18717af14ef2624;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h847ae208ef7eaae0d3e0299ba6d10e9d336353f4d00eda32d415d93e6c11a3b7c26940d8456506041f2950eaceebd9b73c132247a56720f64d8226e9e8dc0dbece4fad3f7eb5c55605d0d3e66d9e69080563b2cdf256b14eb3310b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3719616e87d418da24cfa8127dc2e62b62838ee71973f2841094ab1f7e6779acd86ab60bdb5594f873f6e45b1ea46d7a1861d7a4eebe1ae7ce20725fdf00055880fd36d3bf6338eb1083f51aa06e7215e46cab7a8d897d9ffe764d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f34d3942bcce175dd093b13327779f63ab89d5e156b1e0bd6b657f578e404dac0893fe21f3fbfcabdb83fdcad89079e7d06855ee3131c2cd8cefa7c1e898e4904cd4337f26271881d72917c7f81baeb1b4b6f98ee07c1edb36870;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75f07d4fc436627aa20bdda4ae08699834585636b7df54c7d380f28ce7ee5eecd127024a76ae6c140abc7ff6c5aa62250234d05b80fa0ab5213c1046dea1138476e952da13e81f4afc0c4b9406a360f0e326d4202e1f5d715bb976;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72b80eea0af5f6a94c2e1ab1d9b628e3772f43085d10f6e475cfdd196f53b94685c8c309e2edda098d1eb34b40dad13b5eeabf57dc96654f1b169afa5adb636f793232c0021798fd578f09ff89d5f9ac66e0e32f6f619766e4db67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fa33f6a7ad5b610905a18f4b09e32e17de751d16a420605e69f09bb891f1f1176fefc3ae2fc619b98ebd37a9af56d855066654dd7d81361ab7be5a7873029566d6c689b6eacb62631aa5cf56eb94c2c3267865173bd0e4cf08317;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19398aca97d9d1270d4e848c685f93920b76cd49ecfca5b79caa418b2961665dd1cbce59519dfd6bd08f9e2e132e619d4a0c35ef5396d36fbc195630eb2e2ec3e80a479cb8148787d41c2f54230a16e7af1a65fae958bff618cb829;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf885bcae17029a84cd4fcf49a07aecd2a94dfdef369bff0dbe3b3362f559d38422469dec01b1d914296aeaa789a0fed62c29afacf745881d25fbde3ab234afe56e89ff4b2eca2376c7180a4dc0e1148e07dbeafb1f3451befba350;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170e0207c1d2f24bf1443a946e386d705329917a71be6f010a426e74fff97b91bd5e33e3acaaf26082f35d9b30547468aa3828c287bfad4e2cfd0fe38358c862ceedda5881fcd9a86a405b5f693c7f9b286a0375b3b9b910daab3c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ed784ce28854c013da1e28bc63ccc2cb12d66654f59359b1b6eab6db6eced832edcc56973459774213737658c2d3f5a543fb9299acd755b07f776931db917e3cfb19a0bdb1a5e6af91fd7ace443cbc7f2a689869791c84f03b2eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1359dad69aea3fafa880d7cb0aa08c3c7a9305cbeb7ea12eebb5855b87eb1ed45e44849bfbebf5dfde1f45c0511ee3f2ae4957acf26f8afd06f36b841b0d0e172df13a7ae87df5a669be49c7cd8c357100fad4fdf6f3f7ce26babf0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b0a5c85854e70a15598553db5b78d1b3290b7b768c7b76d9fd552da563f956db00d229c5cd8391ffc7de6c0aa354c1cf2ee8392c91edc92585606d068ccf8ecfd58cc1f7691ba2f8744be94e9c8414c3cd14c4bb72aaa2ce5eea9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b6c5ae81cb6ff83235534d0a6aaae7ae50a34c94d138156c3d28a828a507fccc7f90bcb5a216d78e1a18a9124d7eb85ef3c7af2c494877d932612bc4c807ab7f14112fcf0b19de4e3defabaa0fb508c46736f246a8e2c0a6260e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ddef70504b8d96cbbeecd8ad19e5b0ae10e67e7879fbe7fba8a096d150fc3252490008cc4467feeacaac1528c0c402b30120dd8e50663cc78da1ef0eccc4e3f5b136599637fad949f13c0736dd1a38dedc0051df7ae92e31a583f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1495a8e99d30d266d666262b5ea4207e2050344dd56d214b79c1282608f2ede4590ec3609c6d39d894b79283a637b6feb89d33e099abf1725ca28dfd4445fb6f780a1f9634c6147980643b2e4c5379f0f94a364eb8d2baa4bdd3791;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb586cbf1de6781a3ec23cad306c6d38f689d100691eba32e94cca3e12ce4c0a3f2daa890b2012df9a63a8d96c6def46fedafb6b28d3a6a6b3a4107007bb1e5fd8efe9ea05b310235eb25a14266d2ecf433097106c9523c1d362e92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5a46d340f34ea59904e93602ec638edfd97e11b5e9c3b7e19c69a2471ee0f59f2a555563db35ef8a328236f9687e07da6f00ef924e30ed8e389ebebde04fee946cfd4d2f88279d4e65752fc0d5fd4653d0cd0ffd134e745893712;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105b6c2925379d53dc29adf95d156623f222d9cf850bc203861780d0470ec7656905929c42f3c590b884c1a5155378eb0ed2e8a7d4533325360979826bbfb10d51d4e4aa0d16ed13c91c24e6a4dfbd112ead32fcf3d08b63d7ac7e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca2cbb120250bfd0498c0916b8ddb66f8a3146eaa4a7c923619d691eb8489d917b582a84a1b577a67b46250e30a1fe0efa6d99681d40be977bf45db5145db6dd72aaa0bd87a8c92c5237477dd3b82a29d0dcb653e5b2cfe12fb0da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf74b6aa204bf742a924dd51339d85db84106ed84a7d3f9473f48a278fcf7320de21f91114f753cc1b21740050298dc9c529375d2b32848de2a4a5905099d603692c206b9b5e339d3e8015302da4ee7259e283ea187bfc9eaa38c88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h587f2e48952997eed9d472c84e490744fda42bb6caa1d8b3fdca1dbbd0d4d0ea560cc5a2e9f1e320a9247ff36a2c7b376c7970328039e54ccd62be97b469a78007caf1d850e56dd5221218c7499392a356bf790fa3c11161213b7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17193a72fcff759151a45bedfeb39585bd3f1c19891c3840b189efe27e62c605e7cd58c02648977531f7806716ddaee9e9b6c267b02089eb19326325b29d7813552aa5994c938eb01098292b652af6d9f7de581467da222e6213873;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fb3716c5d6c5956c3744bde67d04bf6cba1cda42720857d531914b7b828efbcba0046ab8bfa1e4e3293ed193daca7e0cbcbe4b285366113fba8ca77d4449d8df6be0c825463d433bd0b6c02e26f3576a074fd9c76f4c3d81cc16f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbb944e12d222bff556015955aab7f5fe15dc23f3b5008edfd86b25a9f8d6733c6fbe6c5f89bd44a5bcbfae64ef16c94576ff9a36d4717feaafc988970a7a0c955425666afdf36a91b72c7d2bcd6c6089a4d4316f1a64d7d39d73c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d810a8f40f1b171cf7ce4eac1c31aa27e504913b032cc7c4d8d8a9dced355d8495eff601e73b5711d559b7eb97bfe57a886945ede5910aa8f7d394928b499450abab8b23b1ab694f84fa524b51d3005b48a6ef4df0a8317c13497c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef3bbeae141de7ad71f281ddbecaf009892ae335b59c23f5e67a89d859356c2bf496a2be46088bcff500b02cf76489abe7c720d9fa5f5169218870046a840beb2e8d3d5e45dca08da01654ad3f4c88ea69c5df09dfcdb100b55a97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0d1c7de31877f448e9d8e576fe9cf921abedeb5f8ebb8f2cacd7023b1fe2f30e218a59a4b88d8722db8fc3b07ee2a83bf25dee34e68814a9bbe5f6b85dde25afd7ef87e1d6e4f85ebb03156139f24faf93d1da7dfb5e72f97f499;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf7f7ce80194576165559dcc0b3ebf0c46fcae36597a5e7ad5d0b687cb0e1a5e4927e0389bb2cde576441d31b2a39d603b109e17d060db3a74fb8875585591271570689939902909c3ebbc5923c060dbd2ad8f37204f1629a15fe8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156cafb3200eca8fc0fd1f71f47627ddff13c75ea9fcc154b2ec4cd8cd9786161396f4e4c237a0a7b881590be431f9be63462581cd06d582c984f05f76951e65e3e04baac8022bf33279aaefbd79784269cc5de8846b081b87dc4a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31032d7b6c78604d7f68a76474cdc9b118a86c1f1f763280b65c4befaf76b170d1588e19acabc2ff52fc4525a985c5aaff44fc2e54d36f31c3184960913db3fdc03bc0966393c2480f6c3c4fdd82082fc5a4f7c7b6c23ec186c3f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25e4a69d24ac37b54f429a893170767d201e909b929e6cf4de06e94d3557a252ac6790eb67e795d20d5c2e18fe1451611adf0802c0bfd0781f5f29f2462c0e3afe8b45ef438ac47885449fb5e1890c386e2c17dbadedfe2ce92b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h678b41df0cf359d261a447895e054c396df127c6c2cee2638a877c1897aaf6cca043c62929a80ed1ed5487971a170c458ae3bd69be4e8f57c5123f8296262faeaf6503849e63cafa202fb3313615c3d542938110109599b54f0ed9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcbb07a71e2ef2cc43170b686e327a1dc8952deb24b1209b002bfca0ff9166dabc9c1fe684b77333897f994ffd7f07b88951fc26595159961c9fdcd440673480e487a53bd613c2f62bbdd2657570d1fa1afd447e5836bc1db5fb81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha79c4d51596da8b2d487e5a1280a8517192649e7737ea37dba04826f5103d97c9f4d6492e26e62baf4fc650917a4f87125d9a75c538ba6e1a406d071af2af0dbc14c5016fa4669618be4360ed7b8a0b6e2efc61537b31ab62161f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14db1d71ae1b482839ac295dfc6d8252746c7a82e448cff7fe206b0828335d3ff3dcf14f8c84da02cccacb5356ddaa79f1876d995c7df75a1ba67b1bf4fece86f7e24299a65831cc614fefd634bbd095eda1a316c90d98463e9ebee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e004bcdbb349480aa416cdf62dd50b964ad9f522da6a776c00238a4a0916fecf9ccb762398aacbc0988b0a2d6052627a9aef17592e75aeaa44b7c8f6891d6d581064519b7c9f17699ab2a4090f56c346533474afb81bac976fd060;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9c175c25b7448c9ec809a91609d576bd491915f4017b82afc081dd7097aa9b864c12fa45bc50a0390843a07bbb6b7e273736df51680315bd33fb7ae686a75112891b6ff4bdcaf4527fae49e2b64b21c57da2aeecdded0cf0f50b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f504640884bf762d159848dad77833f7a52595459313fb6cee5eb66eeba00792fb56d09e7075abe087d2ad98f483e0695acd7ab9cb1417bcd62ee25cbe46aa9e81988e20a9048e1c8c131c2bfca06ed6eb28ce2afe429ab269ae5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf4f2562d10aa440e2fff3384eddd12ca798ca63b439c911cffee6eba310bb17791a48317b9c92d04403d7dbddf9d6815d14504111e7b6754e48550ae1c6d5da4add518860ebc487662e0226379a5780b9a8cdca235d61257a245f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f149b0d2ac2badd3e7ac612088422004c28eff15069a176c9b1beab6baadd03523d4619252c5f978a4878c3a91b208ce8f43a547a03ea42469031332c4fbfe55437890c8dff78069ae0ad68462bdc4b6f05b2c068a710db9bef358;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf3f9b7b5479e8d8da6487b0011fd0216a983a623ab9a45dd6f79afe906d3ad88bb4c37adaf37b40759428f8bb3c6ebc08d02fd1c3ada3976ba7177a0368c24d9a2c4355cf82bdd27e0db6470e4546621bc7d629e19af05112542e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e4349a577fad65a94dda80f9d108786d15842df6019959f7ff93ed123a87f6390525a7fbf5af93289663f659da980fc2a26256c2775286214740236e033afbf6ab92c4f0d5973a933919def5a47ffc0afdc8287c1d88cdcbf0098;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11556cb4d4de7ca54c7c0ad5beec1950e7f39f3d905532a63a3df8298fe175f4e39452153811099cf7155e4c533d0ddc4c273fc5dbd67716e094485bd27605855ea38523193ec08b65762d018d6f9d024019c87111975a2301b9d6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae5ba5529346967ede7b3238f3edd2e9726ef8f82ed0fc2b95bc6d6f9a489d42107a59a0f1fc6edd11af70b704827761a1cb183980796d08493d9ed9b42b948374a67a4d5c73c88e8ca6047c085a8c1308d9e36be91003fd68d874;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fcdea1f7422e3ca118ecd4e22cb14a69b6a25ba181671389020791369c8ea440b7653aa27d31f2611248cd7c49cd44a8dec14f155c14852b7209c90179d3309eef7747c530e3a72d2dcae2401c81f2be3f03511df52e687e7e7486;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c93d26bda75c64cf893b19c17c5077bd1d959362a5ee4e960f03a1a08855ed544dd199b6ad57ea936f08bd95a0873ed8109e0f1a4f4964c89a947b84e4ae987d7923a9e032c52bda2b7c1c540d505801997a6c651abc2ee3c9be14;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cced3982ade253d83d86dd7c4233fd13e80a6c2fdc4c42c1393f0def7a3233c511edf0092e223da9cce10e4640874fa64c5aa7a05a3d7f1edb1f327f058a7a9d23beb022bf644791327eb649a308d6ac0a225e10111620cd71b1f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29fd168dd4bf0f21985a566a675cf36d33f517bc10ea05bbf34557bf63f3d7e8c05afe87247f0daf2d838ac7e1d883001a609a375ef2e853ac038d6301a07c55013cb9cb10677d911c41ef18a4e82fd840779c95c46def2be0af1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6fac62475a2dc2dfec539d09b00ee9bd202247c51f54f392dcd9a966070bdce8b0d3673235fe75f815bd4f0adeb0159f6854bd034d37e7f844928e9e6b95177fa81bf9d66f8aa502f088c83d3005d44790b02f687feb49e3d2b40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec736d4c559a817ed2263f2937cbeb69eca9a0cdda61ae268f1558d30fa705bf79d7d57e2e5edb6a468d141cba8d962bfb88be8be1aa36e705bb1f68038039977fac6e053ce254f8630f909b8f53f48ad3d6b8567e86a7861bd6c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79a53bc3927b34299b43ce37a87a1bcd85d7dd408eb2799b9854a215e04941ccfdbccea8b5027e990a3a26cae1e6c1b4f1295fbdc7e8ff84420e92de6952f325fc07a3ceb5152b0e1ee7bcc8438a48d4e419e157c84195e6ab81b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14010ef112c5307578dda43672bb78e740e92fbba0a20095da098632fb06098b2c5b4c8f879d7830264f81d51e58e187a88885a0255a5d09475a7ea748fef7af5b7062f07afe4bc1242fe84fd37aa062e3f41ab184d4e1841341f19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c1a7a38cf72f824fe667280bc98859ee3b9f7ed747ffc157fff57731a2b988418d706d6d836522f2896167cf01b00acca1bcf40dab678aa73d5e576929cc153e78bdda5612003e2f23c36e7a7f168f4539eecb8740f40ac1b456e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1774eb8b93b4546de3886667e282925dd7849fad1b4ee3d1890cf5d63ee4c2b22363f128308fd8a8bc9d46397e042a33dc0acea52f66cba4fdaefb58a5b298ed061e037e0b579eeff518eb0b6a805a5968e10a3d97bd40c08ab0639;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h282a86aa59998f721720acb47830d216d7e305e1a1b6e97f8689b0888f3c7b7ddee2dcc1f34f4a7c3b3641ed1306e2a408f9041e447e381900200d109f3ec715a24dbcfcd8140ce57f355dbac8c183c0f0b347cabb2204a18ccbe0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37fa8f407bc72c16b698465053840de069415ba71b6652ba8b75815295b0bdad323194be759acd2154d6992b9b1d106ef9d9ac6f0f64b229890fd93acc788df45a9340378719180a29f6030a6da0e5eaf530b49d0bc9a4cb9e1d0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8b13b6c0f82e1151327dd2fd8ad7827dc577b191fccaa6bddd4d348d0d18d60eca7dedd9bbbca1fd57369fefae210f5685cfe6657ee83c0720f3721983cddef65bebf4020127efc5c964954154a63419a795ec78ccbd3d1840e7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4693f561d3156130f68bca340364f8da078de8e7edfc2ba96bd5651018c374d5dda2d0a9b314c3adbc83d97693a7ad96274fcca2eeea6a0de3716fe71529dfb04159540f62b5dca32f1a0cc75fb5d67c191a9706490cca5bd8684;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b633f1a8a7e4b04afa378dbe886f814ee229db225793d0e7bd8b470a51bc641a456a345fb9c40480cb3ed0a1caa21b71f47b533e72f73eeb2aab88870a608a7654134f3370e61f7c7a3d945d9dacc0094f8f8d0f72d5e0b55511f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b41b48bc181c4bd0ff4d23e939d604f0c7734b2de14a08ad185ddea657a778cb30da156dc86a7bfe72c47ec3343ff1b0cd85c744298d25ec3d7ebf7d43acd3c6677922acc9652f8914b598c7f72ffb78104e5bdf7d33861d84f25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63135f82bfaa895d78f39cd0537dd1662b7aaf79c61f24ca012593cb231dd662433b06225df238e0cba42cba61c74cdddb253acc6414cefa50a9ac590f94e35da733802c4b1e314e3650c31a08fd034dc476b8bbf13e3fbe456271;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bca8776c354cc62c1227b31275d2123041b4e890e26ed6fefe6c5f9c16f3874deb64bf3bc266bfa6f1c00c94c8689cf9b86c83b7fe6b456e257ddf8e494784df02ccf1add89d284cba6a9cb2f180412e31d5f986bd319233fc7eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144d93b4563005a3b8e9d57cb733913fdd770dee1f22b85a72fc800f428ff0e740521c83a02487e39eebf7abbef4490ae7b183741e72f3ab611dacd44bbf174243b0763a2c69a9dcf1481db33da3a0eb366deab9c00e4b00a5c1866;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171e46a6991f684b25357918b73fedd806aa980632797933a3cf6d85ef457a62c826ef4edeaf935b28304eea731d2202cf00217da3cc96c3d3f2bf04f7841008e6cb7e1d55de89485e089862efc4b21c65c19a0788aff6575573281;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d902c4d5465bcdcda88d249cd85a848c44c01a74fbc6de0afd1ef4c590f135b55152c1f3b7af0473a8157c5a888095bdcd3529080cb25f163c2398975d9e6c4cb9635d315c5d72861a0dc924139f596ccc32f11c7588ae07f0f2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90745a58bc7fc1588076d7f6144913b195180adbdf8b89903ea1ba9d6e67360f833746914741511d8bd12c74092888774b475c724e96eecfd546e4c2d830e94c3e6ed122c38a36d4aac2fc63c8b241d892ed14c0cbd3441acaf954;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1e3c13816e991a8372632d2b74917b2d1be6eb323d662fdad28a1a10aa08a9ca10c3ce6b569d3fe9f25f43f64e4c57acd7fb4d16869c8d3381ecd84f1c35179726d70eb5f9828bfc8f7d24b7906d7d2555236117da7b8b281aa06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9062e2a29329ea2e444f5709bfa5553a2bedd7d397404b30126b79a82acb9e95c8c4bba09522487bb4262682ceff5b40b2fd87649a9ecdcc3296bccfb9dfdd5b02782a9a3faa7ba1e0bf4481ca6a5d6143a634e34bca7993bf2eed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171cd0863ecafbcd987497939e1203daf19b6d9080481ca3827801b6e8977fb8e712c34c4de96803e0dfaaa943d06118c621f7c836642d80180eb37e1fa8ec08a54607e6259fe7f0704b439d585a290d4f501081ce0d13fa45ffe13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1739bbbcaa2eeadd334b668d94804e55ab7597476032be8186f6be78f2d533b8504d9990cb9e3b121ecb312839d6818c8029cbc313e8a06462909fc08fd4bfeeacc35d4782111dd63e66f994cd6f519968ea54762a9c84519b86346;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcce96b15012bad6f63ae35a6b67f35e054575607b91cbdedc1f7e72c706bd164ff295d6677460e46d8a40e731bbad424e758c3f2feff60f6b5c1dd33e94cb2545d791df7188e79a92bb393a501ac47b538d5c5d549f85ec6ba057;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5f28e35de030105198dea91e50bd2096379aadde6676764d297bd69a5077e6d3263d4f88420d8c641ed08c00c2cd85144cc951ee28720872700057b92b3301ff006941a3fba75f7297fee6d577cfe40e5c56cb15e44b65e0a51f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3437ba1cd4f854741ce975e44e90bf1f18c6c1cdc70ead9ca67c0a54992c5459d7cb8c66abec12995f59d8e6f86e32195b1faea0587ec5123ad6d45fe4a5a6ec92fd5c44ef3226c641c403450edf0f68f88f87f75581d4e39d381;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e20140c84a2f6acb36842ef3450a192bd70c59610404d5ddfbd5db4e1073763068d1421ef137dc8bd3a89f266754b119888d28094c910fe00b047ccebc4e5b44f2a9c70581e3de300d0b9a83665b9f8305753c6368167ed2f6a29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had10ee094b92b3fa944946661d5297d61a4d44f874c2d5fea11e3fcaedc6b24c9966e7d4ef596f5098752a0e652638dd37380f7fc5c695528e4b18f649d5413a016e06902b716ab761a3f59164fcde88abd8dd9ad2c2fa1da22b98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b539c3b4ef25f69f89699e37a63a40b3a7ae830eb3ca28545f7720050f37b59843fc08231636a9cf103d497d55cb811f2b906359e65707a858e973d6e4df606a4b39e07ae1143c39950cbd9eca8a2a548baeeea4a744f76e9c53e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a82fdd8ca50de6371e73957063590e929bc6bdddec2f8fd884eefe1278bd963c5a3a458fae3a65d5fe46c00aa64ab274065efe9b02dbf6ba8d3b7039c31d8b0c406e0c340f8d387267e40721836c3992a0ce10e930017139b5df8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ecd864157fa2ea2bb4605c09cbd9bf406c871f2b5b736edf2369693f036ca03c75f413f17cceff869047e28b4d5c464b4a06b40ed9443157985c633e718ae2e14f607bc23c1bbc50ba5090283325c3cfb66b5f745fc96eebba992;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1105c289172ca7aa0cc3b5e16e959cb133becd773e9fedea7d82aae1faab5d7c446bec73af70316c10cd048d79241b23613958a343db416a4c0bb2973b69172d71d1442cad932d00e8a36e7a9f1adb742c6cc295336566eceb58150;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0ed0da519ae4b0f6c5b06472e4e69b6d58584bb7294309c692e82d92d740042b6ffa588b4821560ee9763a9e6a22a17a19bc7057c1dc118a82b40d2bc87c425a7e6f71654d29f290776c15088e3d8a27577c02f49db71c7e2ad3c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf198afeb8e3c621cfed04df4ed14e3fb7fe98f46e90d8c6cb7f7c9f8ac02f0e46abf942933170b8b97fecab26288d5579aadfd4abdf678732db8d54cdb7a201908f5365b20be0fb911c787c8a65f3d9fcf1e5802a19da72f51cbb2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102ea2b15c26ad3cf94113bebaa1cfc59371fd5910ff2158827fa43cd4f8df64b2005d8c463404e0352ee293195541ba535d16aa28d2c14035668291e6ec7659311614be12d503c94867e631b0a90cd9183dd7d15f6715959067557;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a9cc47fbe502c74f08641e46c251000cb2287da9a5148aa203cbfcc7d531a6e1a6df5b28406d9b635d25bb7f4315e1dd0473ea7b44b4da59fee15c2c311d72596695aa789a9cd64b05337f256c5a40da2dfe5ca268b3672c86067;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd18bdad20d014ddb33724318b089bb2521b7ada0f39a6889ab030d4320c7f069027ec10b08ce68c2b5a66fbaa788007c301b0935665d76ee5d31e4dc083e3e543f554a5c5e333bdb07a54e74071ee316c12d98163e5636100e4c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h349bf616b35aad8993ed3518e8e693bf4837ff6ceac98eb4d2d20b166d1faa502ada2b2e5e71fc4265f4f613ef8fa36c31fe2799a5e59321edf31f582c307f96652d60fbc4c75bf8a6e3a976d821192a61c76ade265be95cfe95df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90807c225c8e58081a127b7167c0c26c16fb0c82cf865f485bf0f61c8cd599760068658c33cce14288783d4334d001ab916442794f94210c8e12a0dda9a5fb46cbe64a671648a1c042b10ef9662eb539ee6620c2b79e79ba3e5ba0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee1e1266e33425b0e1ed9efb7cfce7572dc14f50f7f9a39e7e78c744bdb5b68219e8a6f7342a9de7d8011a4b26d1d2b50cac1e02c91dbb96a5ac04653fe3ff3878d5645533145f30fa355d992338e4b31b932d0cb6c89c2bb0999a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fd53c214752be10bec9a4deef7523d171a88c68dad510f09f55572ea61ebea5aa51aa22a4ef396c7203105622ca625479aaeeb6f4348de157129f87c131c65fff981a821580cdef9d394dbbf7142a2b2ceb6a66bd3474438b6ead;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b51b3eef32b69679917bf8a8c9f7ae60de60836a38e6ac165cdfd216759d269705a8fa3dacc0ff4b71f31d0074ddace45b337b5a50f83f5dca2272fcc160e5ed1238ddfa88ac920c93300edce6e70d6100bd988c3f10f393188a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142b2f64dfc92f514075948e321e2fdec8e92174db72c91ae335eb3d7225fc7f496a77f1061a240b7276570ed3edec269a171a3eabe22461d0a628d0bd58ed9e248b298d584e31172afdffd07bb36922bf075991d30610e90a547d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3afbe0861236877ffd8e0634c4d8c585f1a177e873f362935bf022b59c485baf65bf406cb799dfd00e286ae94096d4412dfec1c50f94e4fe4e4b04ff6d4c8e49c3d9c9cbe9342291815488e3cca046e53eeb2a5306cf805727aa3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2722099d037cc6057b16765d3f26e8dd5ea63dd37f6360ab6ffb5f6105b57abc09dcc1f716cf07855071c7e7182af6dbbe8f72319ae3c1f3d382814466cbb8825a61f0400c9881ef8827e8ca0c84e17201886b7c2559c0bcfa470f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dee012da3e0c1f2583a40fa5185d24ff84068204790668200a9bc10c43deb0f2af73e6936500cf6008716e0157b8359849f31d178085f7fbf226701f501ce4cda9e703db8b74c6459bce308baf43b29d2b0aa86eea8f5a6af580b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a774d147ff961ec3d082b4f0ccdcf8477a7bc51cb0406f2aee8023e567204ffc0565c99a19bcd6a1b667586d4e2e0bc9cdc3ba7feaef87666c0c31854a998972b176fbeced72981b82edb2eb341b5a3c3edfd4824d4d520ef1ce1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156135f32926be698abb17336860632912a145df7294aad277fd7704d6cca250015ed2436fcd4559cddc78ecff9972d19cb9efeb29c0753b861fe69c60f1884abac593aea990b409f347749801a2bbcb12b48edef71bcaef38ac9cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1414a76381122f5439e5f7500b6484d72c7c1f6b90c1e19927b13c070f53a5526ea4ec9aa6edc8e90c9dde86f65bcb93d768eef276184e263e8b5b1835950d88137c8ac1edec2b9c5013f5dfd653c444a6d5aa3e326823f7f8c29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49ebc0ac1832488b52b58e1b012ed112d7b44025f25a214944cf79947dd75bdfd2177f16a3eab4dba00e102d24d7adbc887f14f228d9b971ce3824e60c3f3e4a3af3154599e5a37e074a84f27e80673f8a5db2b943b9f54101f831;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c79d28aca6f4c5b547046536e4f5610dd4ec41d0343d64e7ad407c02124b04e7dc67454abe4afeaba8a262d9a48a711a4b244d916059aff97f4a0ae624c0b72fcac87978c4c4c203e44499ae949a8e739582fce592fe4751706d4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h431af5663a462e83efc279984fcd6169845b63a3786b985adc050828c1571e9f4f0c421bc04cbecccc82c8b515052772f5270b1c9ca9f2752583f82efe9c5c325adfc483ed2a09d7df0e93aed4ed3ccfec09326faeadab9d3b47c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ad04b093870bc5d5b26e5ec537a5a9e7db351ec1af551603c5f568c99051fa947cc5c2c1107654484e42700df82cb19713c9636eb7374f75995bdf7dd4743144959e83d0bed3d70d560b3b51041d5b295c2eda9d40f393805fbac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0d217f8e9ea04cfa1f451fb26908e10a5577101a873c146676172a10baf2d4e7f83abe099544ad038d310df8da5420d2074b2b9f34462e04bda070063504143426b597a7fccac5794f712b0ef2d80298faeec76716a72bc32eb4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1146368b4d2eb139d72034b0b63f7396f50c83431681fa5783b28feb559169d54c3a285936b1acd90e4f5c94eb9cda636985401c545598a10759df033e93d5fe2ee380081d9393ad7ee9cf6ad5fb061eb83c8890b249ee7b71be0b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da70fd470e36a20c37d02a0cb2202094576ebc488abfd26b5eb1036ad87383d3e91dfb9f2a0f7f158158a97c9f8ab00e7d73ca108f4a6ba390203bd2a951f32818b4e25cd3bc4700beec2cc4444298831877fe27ee441aa4fae168;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18730f10e6515c230cf10773652d1d1f4b61d9d52bb0186f14b576335fb1fa2db850c4be5141c5543b013287fbac0a1c17fda301d3023ffb8539db4cb3a5f537769a90ae68ec913e38db2d557a55f227922c19bf3f866526697612c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h322d838080cbea8f5b449fa382240ddecd333dc5b16bbcade5c974b142f4758bc82f38d70341b3181d6e11a347fe0ac8640171b6008fd6a9d4c835831ed32b23a53357f47775aaf42c1f16cc37f3b2d2564736249fb789bba57996;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefe06d716ef6bf52ee7c4109e87c6fc29631507daff127d02cd2cb1b2e2aa5f364b15571cfe0d5a4c1659e6a06f890761012daf0a26fff305ead8d2ca8905da6927967a5ae9681d3f06c8d2eafe294297d695469549fc2fe2586a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he62a26ea77a15b8d5d2fbebf75806d3a0d17d2a5be0bd5b59422f3fbab0448436fb7e043ad5fc29bc2a5dfce7beb87a74aab55b8ea469915f73a02b41a57c3e3ffdcb6062063e0ab10b0c083fb5df0d1e6d4405f199478a676e79f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3b35e0933b9a796bd0f8a0b9d3a25099f6179552625a3b48bd6ddab25d638004950c2b15728d395cb79a6904b77cb4462254f093ce18a1b65c47df6262b04c628710bd80b76f6bfb20385ca57f4dec1705a897f202162d2afc181;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17bc7dbb5689fe1c4da15747db7ee841e9cea0a95eb7bc211cb7e00c165a4f79415fa987273cccd5feff1fbcffc3555753adbd9425768ae64275fbcd7a0a9fb9ca23969d32fdc39cf0f69f5a6b4a253f2750cae2414151931e35490;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbfe6141d0c2124786f7f9976ccceae2768e84e23c0a3500df6e48c42600b95fcc272091c9f139fa52fab383278727c142b37bec6463ba464d4dfec10fd3156da24764f4c1474d822717ff997ad9ad8aaad2b8d20aaa76069d8c0f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5b76975dd17f53e14348d9264b4b8b5c058c524b39c61913dde2de4e5b7c4a6ce4548e650c05203360aefada0eea10958809003bc5384ec825bed2cb4c3c038f98f845e0ab3dde97f234d37cdd7f89f1ac82830ad6bf9edf7972c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49a09a345abd7c24dd7d7e07cde37a12be9d54f59d970b99f9694036386682f6cf739b6014c04533ea6485fe1c92e07632fc49955f499a6a43159f308be2ecd8db74ef8f9441be19e8e1ab19cbaf126b923c259343cab27f4b53ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe98f4e5e8c5b93722b6414d54b1ebdced5e5dd709215e3dccd8ad3368491d4e0149e54645918be6dc6b4b6971606a10e91d796c53f235a0d153bda8fb431c3609b85a80accaa16e3253a7dae90dc741183eafdc248599cf93b676;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ea7471e978165b143a5a4c7fbda13967ecb7ce92117d4bc6f5e7bb91ecd3269713d4fa9e189e388d64ec1ba9b6577f001c4a1fb692579ce4a2f130176c3109298eaae8e999c00e24188f71a91e667ba1e6fe556bd24741b0e0309;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1266190d0a44e0fb684a5fa687d2d6188ea386407634a2ec5bdc03711ed65c3259b9554c0cd392ff83a18955df9df2a30d72d47d36a3a9b368729024fbc5fa14113dca86027e5dfa0567d83eaa1e4186a4437d3f637f1e51d31d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6e377e651ac02ba8c60e606cf10456631979f37dbce368c606e92950557e046f6d6eedcb67d7518bf94788ea8248ace42689b10c92cdaea1658222f61935502cfd5b8ca715b09988b198eb6d4bdfbb1ff29d9c8dc6bd9e19edd9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e405441989e900167e3615a12f048e54c728969535c80025774e0935e6ae70eb7310aeebaf834900a17e156e993d4ccba474dd6f5e615d4dd7d9ea4b9f4f57e81004ffc832da87ce8e89d08e597d1b303700e8e060f8afce8ab73;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha312918f9c6a76bcc30b1f5c007ce119ad56d70ff04151c773533a9cf611edb59db788209783eb0d67cb69badde803aaa2340891a1cb79702d277f60bb0ef884ec884a0d55336df3748d80359ac342f082f12bc48047d6c187b4f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aef1155641b5e7a05a2c12154fec32b895b4f8f2d1a5f74238b4f06aa6298118c900b36d6cc41a6dfc0e541372eed7fcc49ed84d202b0f09f54411a353ecf6f607c42a27c205dc4ca83e06e4baec97439e5df1e9dde7fb8243eb53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h208845ab9f5c8bb0a8deb36e1bce65ecaf4a910342046ebf131df411144d62ce65f8422367d11a551028d77fb994b082a7984abd09ab47af83c6e0f2ee9660d8c68cbbf5f92c2eb1ec0d2426d2006cdec97278889c4cf4670125c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0e10355cde0626fbffa005d71437bd0421e519fce0fe0bdaad11ea471e513e8c6fa2c7a8933e8ba3002f68894dfd36ac4ceb9fe9a7855ff4d87729463a3c81881ce5441f09db2311a3975cc7494b94c68a3bdc140bc19402cf1d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a656f044872c8ada403e1902606670c554d4073f28b6724211d0f193253ce3f8715e2654c3fcb81d428eae1040a32cfad424fb540ec8d804c3789c94c44982088f7ec7ea3218a93291d4768d03e285a3d149a77435aee21a60b1bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h951d28520316f0c617d573083f9909b0177ef980752b1859f994e5b7bc92f108cf8c6dd73170774a17faa1a0ec378cf2266b640d975c563c1cdb0632369ee98259eabbde318d7584374d1ad06e1ca52932700196a0ddd20c86d5d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114f4123843eaa0688ea50713215c86ee8ebef31b3b50bc89a0a5f3d152f5bf3c2168ba4e6d0a92a03d3fefcaba1642e1d8b3a87bc4914d8065a0d5d5e24e125241b62ed21b683ed0507182bcefb15b964c772b985db4eb9f302d31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cb43850fc349738361bdd0cd6e5fc6b9219fe5db3d284741b548d75f5cf04289f40bab2153650e7f05f306deaf00379d40fe438aa39bfda959dfb5a98e6762042a26142482e7741699aabbf24a296265eaad246c415ddb4807b39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7aef3ee7628c606a25c5298f43ff098f672950b5c00efc8fb19dea1dfde5ec11e3e1d9a2cf32a1e39ad0a78b49ba48d2fa01bd49e7394895fe0c1059d1d96b7551ff4d548b58c360d3f8ab51b3b757f3cd33c1e3a5230c2b0c774;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf500d5631c5943f024a4c33a60486b7db07d71fd709644107dbb1764d0660300e8f251cbcc8db8407c2160de3973254671ba2b08302fd94e9d4ed4bc24607036d816563da055fd8b6d32e17815109bdc6ebbeabfc573cb60645908;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8ec24d322bd80679964a6769208b72a800b5df4d754f323c03fbffc67cc9ab3635b6e6160b853c0599376bd3dd33fd638767f3b028d9326b6888bd322d64284459f79be0c74e780756184bc070dcb1b3e595575b4800e33c858d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6794e10b333c8604dd647bc75314b8029e10312c1098d47fe8a8076c3973871a4aa3a386ec19328d4cffb1feaa17beccaa0c839caf094dcf9b4320505be3617aa4ccb69b2df05d56ba77ca64a209b30be79f31ba9805be13dfbdbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7bd65d4485595e087cf6ba0fcb00c781d1dcff9167971ab032769385b124b6eb62caca893b6b25bc724c317bc7b734ef0f60e5e163a4acabe3fcc9dc7f7117a21e4be8aea72309c56542931a43b188a2d2a709977734bd4a38d61;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c33b5ed4d3a67701d7d24826b6573334cc34a01870b1319ab7b71177eb937fa1c8f245e048404564874dec14305b25d53841c6abedc15dacbd7af14d14721853818a973eedd485b648fb88c56a24f92276d4b8960628bf733fb21b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0fd61a191c32ec6007206f8f2369efc29b693ff6fa8dce865e536c38c627bdfc4452df40c14709feab7c06dc8316fcaad9adf0678158d4d97644fc230dc9e1ff2e06392e6f834bd396da11657677ab2dcd0cc9dc8fea484b7d689;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1128020d4b1007453738cab5b9f1c95b65f8bb3a3932ed94dd5e2518da094eed08eccdb982726ed5947402d346c58bd8459ec912feae2911848470f1655b7a7053ac2b0a144ada38ab49dd469a3e927bb2ee8b117a965bb6fae3b41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ce1de96508dc98e09dc7d17f938049cf1d0ec987e2ee7f0c0d009eee03deb66e2bfa4c92fc86b00fda6a33931358dc60d75f41b440ee5adf1596f6eac97db60191f469838ace43386f477cf7ba531fc125b18976b519714268408;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1606207aca2d7eea91d72c031bb67ac8145d5ce1a46bc883c982638537cab36906fec6f46275946975d2872cc94322ffc77c042237e7b400e92d5b4b09fc074b6bd650f09feaab9c9c3307500860cf7b638c3c5f524fdae0af1d836;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f7bbe8fd8f154bffe2b3bd74cce9f13619fa837988e07a9451d1b5cb86f30c0996b3d15255f2211c296521e8e32f0201570cdb29b42f2d2d4edeed427ac9a3be33db782adc0d7feb09a9899da3836cbecdb17047a84e804a08a43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ca248e531cee621428329ea21a32e4ca68b9899b8fc1010b54b27fbd7511b2c07b0d2ae344b04f66bd4420a62730fb431846fea565f7db5c739e11df0fa284e097414f998381e8a23f859a0482cc7ac65b09e301d7152f3615d6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb9b10a1342cc325122b30934791a4386ccab7152d0182cd6487034c2ef96bc9fdb8bbdaad50ba996c908744cdb414535727935bfbf0daa6a2e3f8f698db08c3ac090a3b2fe5e923e6c7b2f4ec1155bcc1f80b7f12373e9b04bb1d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2b909d455713f6075a9c50e162b3a439635791d555064c217e858b8b36615e6b417cb7dccac4c9802e330a0831381ad96b488c9f53433cbfc7e4687d0f806b336566dc51f9ccc544fab4726837faa2c9af8eedbac342919de1021;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc96c774b76ef46aec61ae1b679e55f61c4b721e3ef2a785f1a202cf442f34dc9c71c303abb1ca8ccc4d044408049ab05040a07cadef11e1d4cc04d2faecdc001094f3ded249e6af1aeb547a022db3631184bdbc03c8b48b1ee04aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1828e2b61e72b57fc277b3ec978213e39115afbdd2549a378fc8fc980a7777fde5c1a26a79b5ff65db8dd6a9dbfe1861ab524a2e056f7fe9256078b486e3e58a1b10574f6278345702c82fd3efcda872645d72252ed3af4f2536298;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1894e8ca323f0981c7b8e21d8459b56c7a787bd2e5c863e80ee3f47604bb38a4968abcc17eb00f22281ae75fc9b4d70e188ae7001c937f130da7a03f24202439f29bbcb8c0f6e27dfee3d55fc17601f267dc5d34ae795627cf343c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83d9f6ac7ab0c10ef2791dbf4d502512cae2f492e37bcfd42d5343a45a6d8d2b5f5884dbe31b5cef76ebd929b0b643b33640bab508eb4ed8704a45119107e714ff67415c1562aa4f41980f52f0618145cf5834dc99d48699e68fab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9aee4d0a565998f353026a73dc341acb5a7430b4fb15b2a6c18f375576b85b5674ae2e64c5b5a4ac3304f74c01213051b2e5c9a3a36be4613c72cd28067ab8aba81e9a657fe2c252d7a8f1f63442392b71fc909bd74281259731b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e703e8ff53982ad121c0cb8ff3615a8aadc3d7959d9b18056696430992c5a1d7b890b7da816f8dabb3c6d5a13f222cb4af1fd04efd3c625fc0911b4227d0bf5590a6d2e643efdfc74e4ed936fd85320d9787d33868ff16263a26f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2aa2551b9a6bb461b21d21e6940cbe82dcde6e355433f681952f97f104e144e7f198fd07c6abcc1df5582e73343e2e08d393781efed29af62273f7d38b9f90b2ce0ea9e0e2bc8206dab7f8b1508d6c198d0e0e6c437684f1853a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdec03110d0dd005febf88ae2e06fc520949c7fa9393e2737ec49e1d24ee611c8244819554f8a6c1a87c90aaca675d55928e83e29176eb4389685ca5dab5a277fa67cb911759ae160a8e2178be314a7d82246a84a004a1853ff8c63;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9a8c2fbeb75462a3b98b0fa949391b29dcc537b4060f45780166381992b1e3ec1b983f7b750f86af3158699ba4ac895be27cbd0b354a575180d571cdd9fc6dce59918d1789ee53d16ed276854745e00923991b561d1775fa6bfe3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce344f4869b2eb476908fb0b588881d3d514d69de637f571cf34bdada0e67026f2eb6c2bbd532174d4dee964c0dd357ed13df4b4280754ee23436ab50550558aa077d623cba19e2f7998aaeadb901d7b516c780acc2b7eebf6eeeb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184f38c7169c083f65e66238ef4fa2ee0e627a000467d04bdc5a9bd02b5860539669ebc922702c481113bf97e8ae4b7081640a9a3df3a1ab2c41cce4f8dcf3ec178561042c45f035cef535da534328031b0614fd6c4fd361361fe72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c5dbf382b5a556c70a13bb1bfd0df08644e163ce91d35bf71df4f8b3f8acce105a4bedb424a82eff8327cfece6968d1ef61b1ccd6bc109c09b2b6bb8f376182cc8d3a5ab2a1775804e8ad3f66e800ab8ac377a870d073925c03c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf856563072eb0b88cecd63a9765c32b71a11dcd9137abedf89546f0468a2679b36f6dc1e712bd56d67c1f6086b88186cf1e670e7295a6dc854a98f6f5d41740c73eeed34f58461bf2b68a13aef95f056def816d4de151553b2da7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8608aaee7868db4035e898953a7ee6f9c55531a3f5b45e84973c3a08d586bb77ebed07a4e9d9fe206ea88e7eaa5f6720c8c9e274b89dfdfe5ba5c376289fb2f7431bc945d17d3cca51fab8ae3f30d2c334ebbcd5dd185192258f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9f33055c93708dd5b3c1a671778bebe20fd53d6215a0bf544053d6f0be307f254da9406c8a4c8f642a8e5f02d12e5e09f2c37509ddf25f4a79aaf15c8c8a1f25a112a3bbe3d7610e771459c37913cf530af8f3658e49504d878c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1208213899488cbaae9795deeba69291bdf2ac2c271a710919d6c71a4eef8bcf1989ea47a4f6769d48e61b0277e380fc94ae4b46a382b9007e932e48cce77aeb75bfb89ab42f9e48af90a61ce3dcd02115ee91214cb7332b54f2a24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166775f528a867449695a1dd88a93cf6ecc7e3954f10bddd1934d86cd9832dc636736b63ba5b7d6e28634fa51eef70d5e930c997812b3fcfff885af6d286c6dd21e622dc2936b893ebfe798cac3c3a3f8f8fa29644d0b2f90e29565;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1beb264bf766ee09bc07acf7ebc8934be7c7af9c660a233e3bc42e02746cb002488c90c96a78ca22afb199422c8f5a805c94dc19a8d953247ee98e48edb42ba3de051c63ea216946909c04f289713023f7430e04ce646a4e59f0965;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9fe0b983c40cf267743916c5d178e99a92f7d8f7577449e58948379ee1673cedfeb70c720f62e908aa150b081e1ed2efc7ded0d99fe691cfa5de7eb6512f45ec433d36b849ec4a14872fb7a9fdf77121e4ef8c0ea36297e8d97fc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4662ed48b45dedb9504e4560d435a59b39de56ab83fc8e4f2a354d814521d13702c12cba3f3549e9d95397d2944370ce03f4e647dc26f5f082645c84c1ddf3e4ea2762d5fbb64710371e52c42d6ef7097e26b80d007d62e6d2c3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3cb5061be0d59c1a96d18872ec78b421f2fb8882deb729f0901fd6e4d105f5f5b567ea03d4e7674f28c8a9ef8a4a14124d27206e4ed594e58470807b6a53723a14416c226ef3d7f553dd469d3e948608e94979d1c58262bba07c39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbe1b09803d3e0ac29c25c097a07de6a354f7bc1e100b1e353f860caef77281f6fd3c774a54faab4543a3763c362659de0050bbab8bc47d579ca658778beb06ac0dba85018c75bccee227d3627fd3e07c04b20492188fb8b890644;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b4cd175f778ee51a1bfe28d4cf479b9d6aaaf8092081d5b66d54f88be487800876555d685a48b918676460aee6b474150d8af7cef861e5546db9d685076d6b5a63016d0c4efccb2588873b572a2a8e125bbbd65336a85b619e41c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b09452e8d3667a77e5ad0b6e0f6536c8d28a479467763521f0f8d2bedfca0f95fa1b0ae8c14b06853e2edb8a77f36244cc4606146f5cf4999c99d11eb97519d34dc15b10632ef19254dbc523dfd7ab24118ccf6db9bd978140e82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5913e0e076a711b3aec7ac68583668bf1ee8e26d20cc1f47d2efa1236cb171ee4bbbd046adfadafd97dec8222fe7d4c6935f5869ed10c18d3474aea790ae559587e78d3f574304c5363fcf1eb91deddb6a3e2bac850892dd6acd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78e0e4f15da6b8a3893401479165c1415c60bd06b160e95ec5b6934694f8464f0e5e1349d8e7912e5d5fad33c16c9ce070cf1a6068a1120d7cd39db5822161e045760a5f94e1fde54f575cbcc115a021074407a47429a8f69d9982;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7e584eb6d05ca7933823b036f6be09e6b845040e730d137112ca3594738c246b992dec6d95106b12e44e3d179bb3f75277e2ad322c168558f13aaf70393c5fb40b1249c23b37c5fe3ca0618510c5be8f77bb3954ca0ef9b01ac67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d34fc3b42dffe64d7b65f5f241c483337c4cef545f0b6213dfb0c62386ee3a08c3b64dab71d3dd4221057734a34ab784e48d1d86e49be2ac46e360d0fc1dfde39f9e1a4f63a043ecbcef97779ce477d541e67e56b04c070b6b90b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b31bb574dbdf6bf63bf703a5faafcb1a84603528824bfe539d46aa0e92bfd25d18ca68d1a47e556df53f214ebb0f9f63b346dcb89c3494066dacd452577e13caab81ed76e8d35267f3b0eed7db89c4b4c528af20ec64d818e5055;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a106dcfc12b584245a64526b4e7be62eb5c5a599c5cc3daf144764d8340d383c401c08f66090a2baf7f6f07d1b18d7707ba8b8d7f870a95c2b3c35c79e7ea32b867e3046ded70660b9fcebcc0f9c85c83f7b6bdff878c855a8dc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h470a150f98f7d834e83b1089c2d21dfc609514ed10da2e88dd5ea1c94a13359eb9291c1c1580d2187d97a5f9381e43ac2c6ed1097e0cc2e5e34be8107f10c2c317985d131877482bf13a94e008dfec672c8f73755f132d4a8d4abf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h653af9b03907ef2ee08b4509c01ee6f1638307012acd1f85d58ecc7d1bdf20b4a99925167574d719f9c99d910d10f1546c889807b8de0cecb36316e0cf806c1ca055738a02fce3a04997aeb389682d30be54a7cf7a08a201e1df8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1499f9f75fa59c5859c291228cf3e1c39be5099ab4d90ae50c9b956446fcde94060f0a98fba0ce2eaeb966b697a4f085aa4a9ddc1689aff97b31a1858e13cc8b66b26280181af0a12a3e16aed50064ff10d2a2fe5c0609843b06643;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172dc190044dbebfacc2c16a6a1dc4241bd9e88a5bbdfed992245d0362ee97f25c25d0965cb0d0f47573235957f3f85614647ac0c206830205fcba5ba389e0a6f5c989ec6f6ad50cbc440d6d1b54863e003f07ef71452042df78d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9f225db1c8384cf76e5910c343a8dd8b0f806fbdbe83c35749cd911d5f000cc7d393628c5840db21c60c5be890657c3ee3dfc144a3422c6aba1a3c3a5081a264b7f8f9cde0a158ac6ace48bce3ec9f06c17019da4a7db7a9b4e94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5738c02928433777a684c9705f76df2d1bbbc0a03239e6acc120eba5ea31ef8edaa532850602063caa963dbe44aaf1fa083c63394408754a9cf8be59b43feb9b3567ad71e379abde5daacc78a1a10a23a09af508a0688b124bca8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fda795146db44d2c4903c3cf916421211a45daf05bbcce95e83bc758200a7ff2185fa45c6ab52e58b44625ddcca7fadc8344f0d62df3a07875a1d6b85c7d84a4d2a7ba3d34aac1495ed94dd0a03414be623921220101921fe73289;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5f7284655c0910939f3043278a3fafd3b734081a298628bf4ab5ac6c68cf475e6e962e562d5fc959f0c5051e28940fe7211b22bf500da7597979518a86f5607bc2eb25bf46dc981de348276814af182f46e1bb4ff7ef07177ab84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5289ee97763e16101c587314a88d8b94d90c8901149ec9ce89c29f601a2b7d9871655fb6ccecade8a6eb7ef74875e383f6aa832813681b55fff4087269c8d25407632d016b442fdf9bafa08c1464f27cb0005cf78c2955bab1311;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11064eaa07ecf6b61baff569599a5302e4f24397e789f88f816cd297a4921d8e6b721628d92106a01e5b8a206f2c5285bc2e495422c0cc060015fcdc7119cf920024999e50a8ecbd7d7e419cd81889f3540537e39db551065970a13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139cd7606ea6d6788978c897bcf87cf0959f0f6e8fac5c7eb1790f7a5021a1490c77f2da2abc59dae6273550f98394126709aee16ee070248d8021ab53b44c468fa73e2809fe813fc1ecf0a0752915408dc37022c0449979afe20ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h554869159c88bcb7cca6a0fc4e2b252f1c6554e2f3bf60a3cbabda5f697e09631e7a5fc5f59b431a4b008de5661b37dbba011ee83692c886aecc9f08d8fd6b33f3993cb56458f59a0845ebd39d686a23943614e5a33c7169c13496;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d382246f8294764daec7bbb7695a416ecef823142c6737187091792571108895b14d795504f281cd13e1d308fec85cc5fbf323493fcbf3187c0b2aaa44192523910b7621ee5efb84823b54be574e9ea95585b48518e75e3e3c54a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178cd9e470b0aeb9e499259d4dbb3555fc00a617b939650fa68ecbf47fde6c18150afd2fae2449229bcb40e38439f5dc7c0dccf8a3b1cf564895f8af36dafd283f0370e75c31d7c7517eeaf0833064ebe0e4a6b783e8987ac7d6089;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d5403e1fa6fb66a8364c9f03533e34f2153cfdd46c225ee47506e5a7f1e56b53cf14804328c2eb60d4efc6df96763c4cab6142d3639696ebd45b5e07b772006469aa8184d761ae0b6966843548b58660ebc1b3fa4dbd19e1b9396;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e688c05c68a7a01b898f73d2811be48fc165f4e5c098c70b1cfd5b4ec334da4c5af0135690784745932faed2a67e3bddfc412b191637c08ba1177df514acc0d2a2375b7cddab2c848288d3bfd3725f6d698145f1dbc825f72df8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fed56ce3e3eabf2adbc9e2631e4d98ec6263e3d98dce44678c3d7299d2c9d33e1b6c18d92d786860769b9018102004879e1c026be3635443e843a4d2d8866cd7f5b82d9f64baedf1d99afeeb027b5f8cb576e511c0f18aa63a7c05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170dfbca0e36c57cbd248148946a7e7b00c92b2a9124ee565c2b4b7ddf7998fe6a625b6dfc5649406ec2f1b3f7c44ff0b100626a4bacc3650e3a1d59961ca25bc4afb18ca9868f798c3901822d696623b2fa4eeb3fa7d2ab9a25b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6d0bb10314170b2317da899e743429a91c892242ae1c5556cc80444119c71380ec55295ee2615e18233d94e1cd19838f403c78c5d634fa990c0e4150b4cff9b63fbb83a73a56ba73597ba9c50375c759f159ae98864bfc8d7279a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ced2ea820dc28e57452ed10b7ebb181f01eb25f1d25e757158cf75ecf95c71e1ccdb2896ff6a30a4ad563eeb29425cc2c1bb6cdad0aeaa2d3ce84fc29f35122d20d5aca2ec3408a542566f9c3b2f51db8719ac97fc6e1b8ae3651;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc7f37413e95ce781c6ae37356e60edf42151666f46f38676f8705b98abd65ce4a29519283080e799353fa1ecf8e4628bab6ff0d8486d9ab455b17b4733d0cbdd812f3d3b3fda23e3a7775b1489a9164d9fa728af83f88c00a0f9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98f61cca5926780b2e4de36aa91473e50e5cc84ecb8733f6fd5479ded15eb43d6b0892c269aac21908a982f3aaa556aa6daf00985cb574f7f3ac24c50466288e7c7ad1e0d62e8cf50e5992a0fb0e10a935fcfaf05c07b08fe123fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1674e389d6594ffdd74f14a3b59d6af2420b5a7eb9d90384318dedbb0c5359c9cb1cc6f4e3322cee2dee90efcac1296f4a6d9553722697746dea7cf4d5b00053f12a42c6018aa838572081002072b233ef061729e36003a53d9bce2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h850c0a633dcf4a5fc7657c8770e3301c59791c6544a0423d8e78904e649980608d0ebf7cb36820f3c48632bd027296d840863fbb2e18443551ef07f66fe4ac887db718fa946222e1032673e3571a7c71d4c8e5ee20e84622e39f7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha56e3900daa5e116f97cbf48ec83e67dc8455410ea95a97cdc63819139950437f63eadaa2c368b51c0133611f15d178d0178d2a4f073935fa0b3f10d4ddb561b5e26eb631f49c67123d857fc9ff7c000d8e07081a0b5198d94e597;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90b4cc3e03a4f6498824888a04921da938fa170d94f3caa24204de2665d831e7c7e9d2b7fd9423eda0cc6ebbf253fe065dc091b1bb17a3743d88811b82dd8aeab2620daab574edf4da5db99b24be599d84a9a4316539a541910805;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b45334fde32e2fce40d5fce8449fa03a627b16e7906f7cc53684e8014db670312c4974730c371e851ad33eca070df03db84b6939ca4a5567050e0c045343d52bc80d6f71440b10e47fed28501437ffe3c94c0db99aa2538885e32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1667b78e9871e57d8f815990eec13a60811d1b1ed94174e14fd50b8bbab6dc2a69b09acbdafc1c55dc3712305b8fa507a9060612017bc7cf3a8a7c191743012e03b78551c8de641ab6f425139e43f5a072118ed572f857d98b76eec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h831fca765f359be83af528f03b4178c3ac717fc1c31557e0c3559040ca4139720f33d526b9cbc5345dedb9a30d0d2336b1937911ba8970713fdd2d2dad5e78ececa8fb2fb9d6a684734b99a1d0dbc6f7f602604d1df08ca6d3c517;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e40d5cef15a81ecc2937e9c15c00fa92475566bbeb2ff9544c1cc6d6954b1ba237ec6e2b4418fcba8a6458bdec6807f508dc5eee3bc8d74be4b4d1c3ea19359b5d46f3c91d97d3137e30049997e45c7843d8e378bdd3efafc04be0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9cb5aa8e3b58449cf032c72b6ec323d4d7440f931148aeb56cd3601176a908888b1edd379405dc660d5f5035571e0335b84bde57b00d97a676aee80dc4b859d0024dff8454b9746b0c8ad3ca9327f94dc498c9de8ffb0a1ad50c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c73d2b51732fcea00ed9f38262ffb63d0a637a1a01ae3aa8686511dd18d5bfc0672105233e16edf0351d4885f5a789bf1408c948a881f17a6ed00eb8996b1c50b38e4844a975fa571fb8c7495fbb46dfad84b95b76c01ea5a987aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2f9904ccd46a306158681cf9385a5a11099201bcf3abaac1e0aff431906c42bafa047e585774fb6583532dac916b51f10485f6ca8bd7da61ac1a7ba0ab9b1a0e4dc5560d4a998672440b7160ede027b1638a57cc69fbfc9b2a76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159bf81b5196101afc4779f0c261c73f20fcadb452771fbe1303bb5d8aeb3d64d99d3c1601c64b6808c8dbb9eb2f9a06b34c5e2def58265daf256574ac8147921cd72a743b5f527ba3f5f59ab52416091889dee6b0c1f7288733057;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5c7fb5e2f3744a719fb416447037ae8a66d2cc30272c03645fb3fa86c4f76d7946936dd2d23f31a32736f9fba540f4964944331ba74542bed19f4ba58e13152cdf50b06a01393013a38a247f93a5c94c57e9bcaa9a982868bdb8c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac2b2508aa7662cf6a681c8848fcf3da1254f6ef6c44cf09527c8571cff38304925e33e81d2b404ba660caa2fc3fb0130c3eb6237eb7eec44930d1eb2c45bf0d65ceb2b105b745c311279232c0a1cb6f75f9f451002fbc1f99763a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb15b96b71e9db393ad7e5b567b08ba78901e98137e7cedfc918510f6eadbc7555b33366083273a17b8076f34240417ebe639035e6722ef9fb29af0b0d39785272e72e5f1d121d43e2beed5e5e13777d55a758e0614398afaa99de0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha99371a389a5af0ba83ca7d899cb3e1b170bed0096a382850e85ba9b79376bd9fd5f444927de5e0b9a04dea9e431713d9b92030f0ebd89e55451ebe685c100863a9c1dc6a12f5f821d71e4c92c01dc060195a0e867e5ee93cf6867;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b72b2912611ab87dac56d35557caf1479c05541599d72566068a9f54ab332182719a7f1401a6e000b43a078bdbe2355f74a8dec511fcbf482bc809c2167497cc671fc3ca09beabe654213950eebf8223df086c459054af0a917f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h403075265d0419a1fdc920f7492235af73008a22b4926fc3183dcfd80d6dba416d8b8cec6cf20cd4a45f27c139badb1c4aab9b01376eae80dc6a369c15caf22a38c6b645491704e80caf2a561b551bce1bdf2cfb5b0d2517becc80;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf84ca0b1cdd43e65b7940c679d34e9846ffcf8865fcceb0ce3254229d2515725ba6fe9ded634ccaa553894ce8fb43bb0ddf02ee515a0d0170e00eb699e685b47d15cc21eba1aaf3d7fe130be9bca61f38ec7b9667d4e645936a25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb827c3cfa8f4bcd3dc55d660ef8fbc35ae81d0ef4ba013c0fe6c05cc2a666f04236d1a3ea53c4e72f8ec558a50aa90d8078c367120fccd81029a0f419d4beb8008aaac5b3ca3d8b66bd71e4a9982d2b96c58308d20f0d774066cd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h217ce7c0e3219b90cbed432bfa5a3b10b48ea43a7a05728f90cd0eda02b7596b06870233c68400458b57f8bbfc62886d8dc97149530c6445997902d0e3e07415861f45d48483fc66ae2fdcb7f241734c63863256fe015a0c511d32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a32a1cc8af6c53d7abba6c35acb5fff3450cd9d43eaedf7c1b144f7aab841539163cd737292f886d6b9f4138c5db40dde9b54cfbf7b0740b9695811ef9b0eea04e331c0ec41bc174ab3df7e5d14e17ea4a7e741767749ccb8c75a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9ef5792ed1d726ce8cc12c55ad0f82ab4952f8c65af7a1d60007886b9d8204520bf2188ffd14c2b8603de1e7d8165c5c49a6c3fbc8bfc1e5c8c7940a5ef817e85328ba652061414a765f766cc7b638487c017efd7f74528729e67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c2621fad3d6a5034614a3d4dc1d7702c2d54962234bddc8a23c8a4635197dad5971045d65493e7ddf762aabc5906bf2530d36e784500f9f2511c2385df246fa672738c8c51c355727c4c6827cdd7a0bb0faef7601d8b87e8c9945;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b9f58796a31d77086dc9e0d6d50c2314894fdc34124928838233b5a512e62ff578403106eaaf5b12647fea917125ad3b049724edf438e874f1fd52b5af6461bfb824bcf3c7d2b975193c4a83584c25b18dadb929830b08b3949c0;
        #1
        $finish();
    end
endmodule
