module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [11:0] src13;
    reg [10:0] src14;
    reg [9:0] src15;
    reg [8:0] src16;
    reg [7:0] src17;
    reg [6:0] src18;
    reg [5:0] src19;
    reg [4:0] src20;
    reg [3:0] src21;
    reg [2:0] src22;
    reg [1:0] src23;
    reg [0:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3])<<21) + ((src22[0] + src22[1] + src22[2])<<22) + ((src23[0] + src23[1])<<23) + ((src24[0])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0bdedb54c00914a8dd82e253fb1abf2830d2bf404;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b7c6b44cb5c8ff9a8ae647a9fde4c747faacfb972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba50d32669013df6b7d3f41a3ab15fabf341030fb3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef89ae54cbfc45e989146edaaeb6a6cbe4ea37169b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h884357dd0a49e28ff9d8d95c611a519743ea9953cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c01cf573931db7a421f0aea18dceaa704b3cd2fef0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9cdb00b001614b1c4da059ebe4791542e8539ec17e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a6ee759bb9a6a8105115d433b6cd0f8739547a2ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd54c2cc5f1b50863924148c6208d6ceccf354f0b62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192cec789a74312c774c607a3363c0a7de9a408fafa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe2085122d55843c04887adbe12039dcf658558fa0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3be05d02e4a060f509b6ac71e532715506b6985d00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h542c35330746370c4501f00f52f3b53dbc30902469;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3628338b039b12799c71c66b4e0fe919a49bed9b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a6381a263841a2d53a5e8fd3ddee83c4586aa428c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb0ce2d8adeff6fcb7e01aebe4597808e2ec7a7f66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a206afb487f93263c2e943765011c1b15917926c35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153aaf1acf3ba3f95140eb3a62baa37e15b13c10563;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42c38fd3ddcd2e3f5dd17f451ae71ac735f19fe104;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133405e2ebb5df8665cba7d0a49a4eee4ada9a506fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95e7096862c3860fc3b96ea5569e3aee2a43518cd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9a83cc84d7b2a204fd0f08beda851d19d2b3ae01b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1d425283774fde3c546913a010508df69f118ddb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b05fe0abcb9ebe7edfb21574750f7a44e2965148f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aacc05a9d6cc05af3f66a156539f0c920147d14acd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4cb9a298f7850a3850e96269c3bb9e48ef055e2eaf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f591185ceac7875c4d7584e08103b3d29ef050c9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10587fcc6bec6fbc3c4f0ef752e7314bc37074050d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169f95947a7bcd75a72ce6e7c05bbf6f233535a517f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd85d02ec047d8339ed8680ef8cc45915a9e1d682d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f7b89684941b090fd18f6b0575198474a13ba19b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d3820a10f04b93b54013255dd779acaa62fe76993;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h885518a599e41a43df6d9dde746b924c13a935f6b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4915e1632526694b4618c01fb8159cd9755d800c63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cc014e519cb7944929eeaa569309c443574dc82f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a406aad9dd2566dcc9ca4a3c8db23202fc3ff1147;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d25b230858bea15c2c41c751ac398aa96e241767cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c171964906e766c6c80a48b8da4bb9bd96e9ca92b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c71acf01d96cd19c4e8469e1edd08a575fecf68743;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4886c83d4b813d1df3c1313654ad5c9e779275c73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17614cf0761c9477e32043a0c1483f42bf95326ea7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h713bee5404bcd9a47dea53f48670a19cb0359fa704;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10363aac58847cb37dcdc1759422d2a88a3a1be2a4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1dff1eec5eafc5f05249efbc62ed65d33acf24ba5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4b3cda869e4f84ff84a3ca71ad735d2449effe667;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93ee83c7f30f0306faf86b3cc6602164ca54af67b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h752d5123c6d6f14a705f4e44f4dede8cf520ac817a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da6824eb8247cb2fc2f522fc11f6fed43cc8e46a38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1154d6b35ea988bc8ec516e1adc600bf1d3cd234515;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e54579fd6e20d5747ee3d396617f7bd600ce30ec7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d14744c2e11109e088930c129ab3a10656d3565c09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab2d501d72e9e83789f24fbeb47a8f09eb7fdecc82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12af70d73043f662f3b12736c32e9cc020cc2520700;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5e9b2f5cdc848524b64d4c4e5912a3e7922b1f288;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6e3933169667b13099fbbe8f50a781bc75482adc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edae1e46e4a60bb635a922ee9ac0311e9d2defd697;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197c655fffd4f76d25c882557e363542828bc74fb03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2627e9d925b7a9182def73d8f49c4eb9425229d24a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110a12bb3fd63eb62099cde5c4e367d622ff244f24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161a3d142643a11e85eb693d60fc955a5e20cdf2e52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164d818b79c4d69d30d4e3996d90af593bc84c7863f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a370b651a18de50c1ac2e4f094e820dbbdc37dea7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8ff03d57aebc91aca7131914416dbbd953179b318;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15acdf8af907fc4698c38b634af75ac3bfd2ce17cda;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9c176ef3231b94c2213ccd70bb555e66b28e5c00b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff07afb1c9b29bd1d12e0a680797169f61e2ad9a50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha02889e6d762502bbdaf1d4751c0fdcf378a95c6a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183b5e032ca4beac69eadc7d59f8236f8cc66707b88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1250220dbdb76de2e4a10ea0aa5a8c9a485b34e31d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1341e378ea346750d26f7f1c4b3282109848872b2fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c281e299faafcb7319b2d2306dc0a1758c2df3000;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2617fcb602fe8f97af4ce51594e17cb979042fe1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175e71f3293e8b43106350ab5a166eb721c2578974c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165b21b199f9b4c8c6ba590be19391bee10365eacc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6cff6f19ccd3d379d3a77039caf01c402abf85ae2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10007634819ca01f226b27585ef1a2f80690ed6a020;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3692c0b12f1a4e616beba3a80d990f48c4f4734d15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a6245b094aa9697b0da22f65aee1ecbca4aa90710;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19633c8a7fe04e0be9b2df7dac506215fac8443c164;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a99d8730f9f4e940c779a29be12a29e99cbc897f49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9abe11311bcdcc4539730e929868850f130f3c231a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe8de8e04d38173c20169e13d0ea4a482fee167ade;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd8ff1b1dcbb1069359b2a6302fc92e56a796d8597;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171f2e3be66c29cde06e25075029189502444201d6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdabdf9207db7da2b6dac973c7caf1a09e9fd8d2a08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e2b1965546598144f10ac8ba44ca5a49f4f9bd34db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30230f1a8b95a6d35baeb3d8dea57ecde8d8fe2587;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd04dc7dd4d93fac11700ece548c214f07bcd6540b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173180141534e71efdb7d6d4ee4aa2cbc054930d624;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19edc828651754bcc1c7767b8e7389a89b1d768107f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194fd099baf99d05df8300a68510a6885ecad94e28b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192bee8299fd439bdde211298413fec2ad12f6e3907;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97e6b3784943ac59b335b9be58abcfab6dc6a7a12f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he70ab03087477eb7349463878bdf118542a0450904;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1751eb634635119b2944e4d9ce70ce3deeac5e81af0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1dbeb6544997113002bc5e27caf9af61b3721f42c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha9a7cf28f592432c5f74d67994edae0715f962300c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha93f80187d7994ad0ad99da035f6f6d43d69db5526;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193c1153643ec89d5f1aed0ec4600412b9440278ee0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1674c4b3cd6295e529e19558fb9aeaada0c0be05657;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1c0877b4f2b45b60c5219e23dabf9a5f74c1a5a8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4c4f0ed756ad15b090fe5dc4ff271c4b9fb0965b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9dfceb14efdcaa70bd1d7bf5f24abfe7ce0ac5296;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fe7d64a0479056c572704068bce561c503562b8d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc377a1fe30786a429ccd06f4cd2c6987202b58e50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h865b3eacb68fd7aa1950d6bf40e680ee56f783f75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14704633ac0e077a89491eb8204d1bb8d027be353d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1fc4ebaf1173cf933f519b1fa55e94adef6a7395a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1883ea1d6c1f4a62fc1ae390af2feba95ce248d744a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b50618a0e446b6694ddd82f736052ac110cb3a7287;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c989cb165156c279252eb666edd5b2446ffe77f18b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4cac32e463b4d70217104210098c623a8a889f8295;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23b68dd156939e61e0329016cfb9da2a8b10d66b19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18808825fb0db257720bc115fcff13959b8ef3ee263;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha35173fcd2b399d8223951cc3f34c678d8c6c68522;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a1bf1905eebb26e589ade92052b5a608f67ce30d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h303527042f0eff7ce998c6c94de27e899064afdc5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f8dd49a88f53cb466a337aa6a0608bc5c12f74073;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae0c3a02147f84f31bee9bd249e8bfa63f557f4ce6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14adf51ab3688b0b9d303ef3f5dafa5add07ce9e461;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0359393b2fdd9a2422e6a61e4a96dd3a4c3c9320e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1803ff4c131fa06d705850f5f5ab9e27229d75c203;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6027300373316630be9dbea0428cf3a7c2da44a9e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8344cce95e2bc71ca4ae4e7a4b0ff7d2f1f3da9e0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb8f5e71d5d49d72a114c19e79f1953a8b0a8994fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59d63bd8b5a55dbe135277409832d0d476d2647c53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16fc5a45019deadead7e93eb57f110291e15847d95e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc8712274fed27c22bcd5a1a743373ac00e78b0fad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2af24f7f065d7ac91a98c45927dfd5bf529b6b96c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hffcd0497d2fc3b54eb4eeb81c3dec7291c02bcb7b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124cf2be3f20ca3c01c5fda5dcfec47ccbada6dce5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a00062bf1c547214b5ae82eb1ad6f120620bfba702;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95562cf10b4886de3f7de743393514ebae88a85721;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4050ded160e01dc5021c4e22e728d5dd796ebff02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2de73cc2ea1c5ad403916f21721950e54ea30a7819;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27ef919ec5cda71c525f85170f33010fa6c59e2cd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h525c1efdb9360a2900d7116a77ea2995f4e6e5f5b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5a468c24d43f97f99501ae55cd3ab14c245e5ee8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19304ab04159b16a86283343d5700480d500975caa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ac76bb0e02e09aea40c4754a9eef6f325fc0309f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd98b02460f9187924d381ee17bf5b80f1902b64eb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1168ed6c1f513a726175f14adaa3567138b743d87d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbab5bad87db67aec199f3cd263a9dd1f3b29a637a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87f1a2c9453b1c82419749def20b93eebb4cf3a573;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde3bbdc2d1358ec5c7003b037bf1b7073712c4a2b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18926556327846d598c500881268283d28f607e632b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h395dfb68e0bd540159736d0b3714af52d7f9853d1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bada6bc139a95ac91430c859e7682471f663924e11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h446a34194abf39ed666ac58df41db726d206f4cb93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4117d05fdf45174af3eff11564c9e7f2335485c21f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h65bda7ab978731aec092f954df9f3f9ea66f474340;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd1ad5ec0e132c9735e7772c9d3eef94cdadd61745;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a9149fa6712eb989fedf015772efd88ae69033031;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134af85750d95dec79246c472ebb686c94a1a00acce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c696e4c2b1643d2529698c8cae5202f0bd85aa2ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h722aac1b5294db579f8c86a8e7c33571e2ee8d5bde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10265c36eac877177b493935f83fb845487f1f38d24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a477f87473c3b4d8f6b3c07f22010674275cc77ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1755674bbd83f7df2b6d3da1f5a72e8c3a8601b140d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bf6707da5544fe18024b0a97e151b36f5fac8f982;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125196e2234c84db3e1b87e742ddfbd1d7b9dbe0027;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f952c8e55a41eb7a877ed3938ea9450e5986d0983;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc0d03bddd9aeda3ceb2978133e68f06f0b14eda90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca5f8e0b27716120f23a323ceea348e6b522fcaefa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b259ddf75bf803266b7a074d741958a5e7609f950b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1ac204ac087add9e5b8af99aef52b5159ae3f1472;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h562fabecd202a919d781874521af02d74573fd0817;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e27b063702b666930d69a0346ec0897d952bf900d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145f7baa79eff72d2c1ee0320cff21161083aa6d97d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ef0bcd12da67d3d5ecf4f02b5bf7a035384e2e49e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143e7fb8b53e23d2efca494add12dba7683e6c3cd78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f36ce31c0a69ebe4c1dcf0b4dadfdf0614e10793b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db2f979a1004ba4546c7f3e2328342859916480f2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36c8ddecf4a02826e4fc62e2a44c362b845cdda941;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc9b6dc83bc1d8abda82c8256c2503620886a514d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8926cb540c9bd03b2600b25357c37bd482f66f22a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16402505b8399d6ac1b5ef9869ca358e40a02f9c1ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdcec838daf989b44da5029ea5b369e7b318c26a39d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d31f74ddd066f8dafff10f0417238e4ae609a007e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd14e01451cf91fc4863a29298a57bd3148487063e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe876af73e9e97035f561d2abdd033ae2765f28761;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef1e7eb42d22495f16b1f7d34fdec981ebc35687e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b44ea168a85e8cbdbaf57b48f4fafa6c13c27fdca3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c275d8c4ed9e7e4cd65e572d6d8aeb9ad2a878658;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6df5605854049927f490b6835d0ade5a98182e9e4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d6efe07dfbbcd1bfdfd11700f1f83a373c73a4ca8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b06eab64cd04a2366f6b8a82fd6fa082f0e085c73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f9df7ca4bc43e26ebfc4d7a1c8d9dcdec22afa4b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1451ee1dd2e879110551cbb5bbd540248df196e461a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef617aaa5d5c4d10b5b3fad40dca275f98108734dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0dd132968590cb59910c5ad22fda96e23a2e90815;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2ebdf473aaa9bb58ab6e9308fd5ed9e8056cb77bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75235172749a31f933e9461e28e0dcb55356a96fc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c547d8ea2d2bf703e35794340dc4b50df0dd38ba32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176de0a2b02006f30e261e9a59a5b910a03ee26337e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1586a8ec1a970ad095a662f4538f2bfa8bba16cb946;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1875d5e8875399a7957c35b0b12bb6c0e48ca81759c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf61aa4af242b4b69fc622d8f5432a6959e8855b1a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a8f1ba3630e510a4b6f39ddbefd816721a6f8b3fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141fdf21eecbd1e26235de32f082bb114d30143251f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1749ca223f2a481e2ee95f20b2409976bef77905643;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc86801b4a4b8f6e1bbe682d218cc1ce52bf8ce1742;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1238856977bc12e254709a85532c54e5002f8b7f19f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h67d5b2c01d1530aca887812b50450f8e4a38056c08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9badfa0377655b05ed04d58f3d6b8caa343d9e0635;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd7a520fbbdf7f2222877ec03416d5e77a1aac7960;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1849778e657bab6bb539c6e683c9c384e3ef23308e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3333c7a1792c9bb8051aa4fff84aebcbfc00e35239;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he337101c049129aeed598129862ba48b1665d432d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1967d28867634a416ea39763c9779dcfc7bbd91b4e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e91e8d6b5754540574b92629c672c04b7424bf9ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aecc8798849933492eec897071e4aa64edf12c1717;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150b739a4f437e013b40bf68452e0263352ed705f21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f94c955974fdaa04cc7c2bc2a3d64480f8ea79371;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea96b127273f270a0688d4f48893b4dee6693cecae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ac733780630449345e10a921cc531fac2986fcd26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156bc8e09a1f05a574ce6524ead8fcff9b47ecb3021;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb458b40f096a75418f5bc76642c4dfd0914250dee4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36db6d480a8549e38a5d9f516a771231ce7aaf1792;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he548941fce5f1ae7b9efc1a4865f9f82803d804b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1593ede04d58db8710572d6b0528939793a2a9662ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193cb0a84c66d628457f4b11562d0a42c5e9ba4aa9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1341ed0c0fe12a62cc592266d326e231988f272dbea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h189656bb67a89cf25267fda05ce6c89ab42eb07e1cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86b2e7d1a29873fcdccc3fa4613e73347250e2522f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe49b2aa8dd994ac69e3a490e10af4f7a0bd7fd93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c27f6be449ec83a05b55a266032d03ee6c93d3ca6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159b10f6f7d7fdc96e0dc2e4287d53ea0702851636d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b6b992acb2971bd65d7ae4bc0cc658334c5ce478b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164d1e3b540b5070e5ddb129a00b7969cc655af86c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2bf18c7293d4a42922d68275ff17078df48f257aae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11783730865bf4a37555f2e93c7c203125c051e93eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19329997ac98d146c280cc3d267d4bc21a44214404b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbcfc8548e4201cc349158c651481a114f695372294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec6c63faabedabb49e05bc4e3180d1fff14a6a741e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd11fe435dd1ec958895904a644ea34752b47dd31b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b7e4d5fe261051a7ba0bb94d35cc3acf53f6856d39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14865b32e43ffb22786c4e1af706d802ad8f9528445;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f25a99f307239103c43c7bee3761e2f0374cf342f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf33311aa685a870d1763a95222a6147995be143db9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h665b36c638e0ca87f91428198766aa8a2a09d98f76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee2ad20120fbe403d3b2ad1f072accece9e4bc3966;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h851f265ffeb42964561c1d44982dc0494719984956;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfda0e2f1b6b6fcbe2ce9f97d602f0dde7ef8345dac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d4f94ee057b9eabf75b473cabfe7f29842b3d7d9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2a6145884e4aab4e4c268bd8130d71324a2b9144a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106cfb118fce4c3709a039ec81f9310f24073ad6096;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4087dff5f2c64cf94349c410542a650534c367c62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89d36d7ea484ca585df9dd279ac03a8083a5162b37;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfab6c6ff558f009f41aabacb06904ceb30793a1a8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf38a4ab351eec5c57b77052f57b79b74fdb66d701b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42c777b8b472184ed28d2fcd078963cfc5543f494f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192142cfde0d1a9c7d07467b65e9b0dba1c2cf13579;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a93a06b25308b0f2ad23b41ef215a93861a52791b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14507e287f3bcc074102c7a119929b5fa3f4566c4c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc29201f5f1822ec9189a79dde61e5ecd10c47a8e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7f39fef7bea6d904f56fed6a5ef992e260e4904148;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170d0d84484eb9b7321cd740ee7596fd2636ccbb8cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbcbad350557fc60a217cfa8d69d49d0d94613791ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1240b7aceb946bb0858026db43e57dcad1bc19068f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81b697829a05b11c6d55cf5e4f0d7fe0940c7d8828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ff7b16234164c22087bfc49739f65ead057cdb82d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157d580a610f0788c1b5048c255bf092494051d79d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f2c58e04c472250a7f83608f5c1832704dcffa6d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de81e2b6d2e82351e0e67b7994caa8d9fe3089cdfb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192d2f1e32a6845b6e65c390f4c6170566db5a1944f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137ab43af188a6386c58666bd6909c27205991b0c8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5e29d10a0e200d9efdd5b3c9a74ba2aaa5b8d2ebf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e32c8da159c152289c0ff11ff312f933aa0e52068;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e215a583d34975c8b6edd716e9e1c1016cee81e05f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199e81f2ca6c5f43d022b510f569d90b5594bfd8862;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h992a919c79557d868ae56f4d6afd4220a9d59bf246;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11be9198abf9b2900d3f7dc26e9d9ae77c3aaa46d0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9e72984f73d61df8b6124c6bdf6a674b09c79c53f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb21a0fb2e863d2abada16bf2eb1e7800a10f792632;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1504682ab7e63850596cc081ed17ddfb999f76e70ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e62929aa84b78b97b079dbeb843d5455887e4ed08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d5d5c5a5dfdbca2b1495588ca9ff8418e07912cb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17bcdf60001f31a15a19b95bbacb56e778395c30450;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcecfbe6cf4c33769596c61ea436e15f491ba9d703;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h757d359bef796c078f9ae0fd3150f8e7aadc9e83d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha14d1de4d7835c89244ed7ab3c0278165dc3a26666;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e02332ecc3cb067a9b06bba0baeade50a0165bae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c473783ac16362b2e8f7d30d3235e682656ee5744;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee62bad8f2f9dcdc3e84310d25fd40291b46f3b2e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h501c8db51cac3f32d76790175aca95ca13a37f6954;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f4d9a9190343fab93b9290fdaf3d8e41cec9c08a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52f635d65d7e8331fa019a9380bd7db8abbb820c72;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1b40fd02eab27504992ee8f7ac0a4f463e3a486a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a67d18968bde3ec509c98d1f85e2f59998d490751;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d4bf53aa8da9b31be7dbc1e5b66ad8703b6a43625;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a16badf8ac47a35c913fed9812b58b46d334205515;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d07815ed5259e4254049cd9e8d3027040a4a4c996b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aab4692faaf3c5abf709e9b5484b1482fb6bef09d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5581596a72aa5f8bfc009a293491b6e5b69aed5cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e078caeb460fca052947b42a4e341853949dfb94d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d123910ce71d1a750758d1905c81e0e5d132477bf8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h534051a274b7a6e4db69de216e77026137d9ac0b08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118a52ab641e23d872b6a66523c485ebb5168c13ae9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h332f9d666c32f0c35e08c7439fe08c1db15ef229f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ef30c73cd4625c006ead4b959a961116b5e1ad160;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35efe381048495906e57361279767906154a5d5bcb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63549a5452d9311c4e85d08eefae630bc9c3d80ad6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118c02cb50d957b9f785d6d2e96d9125b7b3fe4403c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130edb5a969388c147e40177dfc40c4ec7fe05ad580;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5aea733382ce07427bb2e34a88803a115c0635311f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33637aacde0bf7df2b8510c2501a3fc568cefc8e9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbdbf2fc2135ec17da6657c7d6feece231dba138f42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ed792891edbe13f4068f26063b08233fd930b34714;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118e1f85d0c75ac6623059a92220baddb2424e747e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdffec7c29fdf82f026283edf2a97714fe44a7e4154;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171f09f27da3c7aebdb38ce81900fecb8d3634b8ded;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30cfa20bbd47d45d2410283e9e26b1d347acfae192;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ef9eb6fcbddfc7cefa5e14bf06e6a162d67036bc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h967e949447b24765c421fc9f034d46d8fd98d5fc62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha845b215cd95d41826364a45efe3a1492224a8db7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h264bf68aad7ec60701e9bbaf05c37c699e88799c15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1569ab34fc0c6614031f3e337578fa3f334fb72dc6e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ebf030ccf69b3ef4a8e5439757c934b10a0c5b5d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f27a070287b14509bcba5e6781a4d348d5752b109c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c5e06148d8b9a4925fc69f1fb3357a4aa98ebc090;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145e5a2d52f94772bc2684b68337a94b43c87235b2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15533eac60e2f7173ef92f5921d6c8a006f28d82ac6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee4a8563d3628fa4575a2ac34d422fd8ced54f42a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce7ba0aabb63bf00685c5acc0a32a95394732f1d4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19387a6fee5ee9ced9020c40f39b53979663cf43723;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13359052d0924d0f5af64ce47e245a7a7b1005f047a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1761f313ce6956e998636f9a07a4c625487bc49b1cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bb7a8c88183db9b8336f8f36aebabf3d1feb2608c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18777faea71939b37d87fb0fc9a8ed294ec0ccd46c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4097898d93c65fd7f5b09eb9d970426d157cc777e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0911344374a9eff270d854b550fdf9d1038194e8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5947728981ea611030beb466224cd61db9054a867c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb72cf4a03b5e40a71081fee0f1e90988909836d896;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fdf4bc6af7948828abc626f959ee0ca443fdb0f531;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5942675804246c34848fc925fddce785046bfe2e99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a81af556705ae48d1e3f1b559113910ff02520f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h940975c361f0e0ad8f24160aafc33f87ac47402595;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d36b59a7fa3f2c36e68e769dc69a50dad6e776f51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1908871c98595fccfe2f1b5a911c493adaa67cfa00e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fde793205db23cc250bafcdd51e8c39023d0fe61fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae48c2966ce5539ae529a60bcfd1b5f21a569b4e4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3e8cf668113a47f9f1e015a29259d9dc0b70feb1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he83283d2c3924b6b9b59a76d38af22cb966c2ebbc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53dbf981c08c60c2bbeea1f9b5833b13ca6d27a4ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffcad2aa574f9c6ef67b3137ba623c732c57a087f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c383da60bab1e362068c50238f22236d30807652aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f545e7be69604d0f47fd7754630d22f8404da4b2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119f19126521355e53daa3624fb13f0dff9efd0cb39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3916e7bef5978385833fd47f3752b656b1cc10462f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbbf882c693a327767062d20e708144abb73e48d5ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f43d339ecd6d5413f6e932c8797bb0775b7e30047;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5763e63e6c35c299a1b2ac13aaa372969fbdeb63e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142a5db4b590921701c7c982114532d26a3367eb3b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1118c06b6ed6465c1af094cfdb89186bdde0e1ae5bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8f4c34b1fe679b313c3c943290bc5971a085b3020;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a9753fa275e5224df18cc62a8748fca1e16137aef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1070e7c87ee6f98fac095aa7858f44312e08c41a4a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8bf655566f405dffa5760cc60b127fee8abff084b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12a42805c2352aed52212ea01f177c493b4f391d973;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h96c683683ffa8f26c772a9a7c529ea6ddd1100e851;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1706e9c69f5510b424cb69bfd0ee4cd9f9704192a91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148c8fbcf19531df8e3b6be7148eabc061b2212a214;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d37034d7db6d70b1ec7d53efe6179dbd66b8d8e33f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59f8b54da13b8a0bb5f85ba871bbd8261400b58957;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha61a39399bc7089d7b76f3f5fb09fce6abebb88737;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h109e8c2e3493a932d0b68a2bcae74de2e33509189ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133b30a92ab76751ee1bf9be2cd7c279f000cc82ac0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c0dc10c9c9ac703a6c335b7f56b8dbd8db518a1c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecde63ff7734db55d868277aee02277d03d2ff5fa1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bb1165f10d9fdffb0f3b465fb2a7ce344c64fa13f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3bb55c9e954bb0e2ed5da8cf4bb49fadbad5044c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha13da9e5a2cf1ad46ccabfdc0cb53cd8b9b7812a6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1866f2824a0b1be4519ad95611d6bbf56d74f8f0ed2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8f597eb63931cc32c6d9b79adac2821c3dd9fe9ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b758a8e7f86a347e6afc3d8a6953e3a5e2a14ba789;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e575138d9d76bbc12c57784e7138335200336160c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41946ac1517f857e90a76a3af2d31296b8e5e3b040;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd2a8c58b1547620f8537aa5a3ae522196ebbcc479;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51269bc7934719f162533bbd5a965c90922a8377ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5adc40bc7f3e7b4d6282fe173bb9954d68b588a35b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1668c0f3bb3703c7570ae2d79855578bf5709f9e762;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fac5c10f3876cdbf45b67d6e420a1db0e6a08999aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e766ac3ddffe9f99ef44a8bf5ddeef1ec495109451;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113a7e7bf8298d1b08cfabcd9b5ff2ab211327bc522;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6fd2c124c84e7b3d7fc31b800708d8ace8cde65e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198957482c15d5574489f39aa08f750509e920158c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118cbe20c9daae080b09511ab78a9b7e9286edfdcd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3ef23c818abd85c64b98f7ff9bb94aa9d0bcde14e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62db36725e6f4f33bee2ffb3ab1340c6c7980bcca4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2889683cdf7973170e7b6e248fbe11ba226033bee7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8893786f723578979ebe3f1d004fc52d5c919b35a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h787ba543735d17eccbf739e4cc376bb044a1ce61e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb85bcd0a38ebf54cbbfa14fee1ab501852632cbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178d1de80e790090db5cd5a5f435e30dac644f0f0e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16495659758fb1ebb45807ba723310056308bd0ca1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f460000465ce1788baaf8ce9158d83b03ce9260ec4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b719d466b69945d7d9d741bad5bda337dedbb62212;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19169b7b1445b841ff30839b0dcd7b6025daf5963ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb28fd8c42ef6d44ed233c4ac136418a4d7505773d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1160bf353b3eeb0558ba80aa2928b011e50ee354f64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e65aa32f3b4f8d67c7b727c2f61f09a516f8977273;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48d9133978c8926ef3461f88be5b7032ed94078f05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5248888e439e5e03d6815038acd7dcb930c592f53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b58e03e7daf2e3ea4b13a4e4e0a7374337a074eaf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c3ec61d2721e2cf102bb1e471140b5c755017dd0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d3493ce94bd30e5879cbdb43d51c7adebd97e1d40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c93556ad2c45566bfe146be1f490f8aa3c2afd620a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf587a26c99dc3b36bdeaf8ab66841c55366dec4479;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148949fc98d63af3b0912aac63732a562fb9663a6b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e6298341be1403399081a2c2ce37dda0511d5c5ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1499b90371ea1be865a9fe1ec6a1e778d640e075cf2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea51245a9f42022c08fdbb3eb3cda7ed49fc0a24eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27281d0d47faadd10685d0bacf5d29a7d9d4cd0544;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78ae673c277b96e8ca0f3c0936753ab10550ee14d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47018a5fbe306a3dc3e109a5e7aeebf6393e890acc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1984867618d86f189c248a326e5bdb2ed26ba380bbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4fee652ea36493e92ebd5ff3e285e5446d8aa30a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7d737a4d62c5be528eb0f17e1a5fa9860ecd2a569;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1847273d1d8baa0b8be6e54c8b2c751a7035f1a9952;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f21649043e6bc4fbc5b1ed82ca394c380d19c6334;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc0e3fef70f50125bb371bff88580864ca6cde1d1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a586a2e460364f398fc40ae70451f309b03508462e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bea56336cfbd1a4e2fa9c59073524a2fef2379662;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f1be2117db76b0460dbc2bd6815f63b6ecec345aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11aefc42c211025ea6aa41dcf22d0839a3cd4e08c1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15929edae4ff3274433898394879a0923c51341f019;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128617526c91a7756d67655638fdad775f2b97b75f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8c78988f7be1dc83b3d3547b7bc2a8b03de4f3dc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1684b17f7fce8e0a9c395a7a0948fdf4074fa0ab57a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1073939a35edbda673a6da76dd06dfee4180d19c589;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e1868639920183d8c91cc2c220bdd4359dc2f101d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e6773f01128ffc7256fb7f85b55d23f05ef3eb09e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fcaed65f05127b687214f0add3f6ee82ac04ebea7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148e46a8c574d8d07872e80156ffe9aad140a98403b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5b755d0807ee723ef1ed8a6022a0ae7258349904b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c0900d657dad6e5790da8e26b0fe49fb337ab6fad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c005cc54c73acfd381741c5e018ac612fee0cc6a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33ed2eb4d0ac6344ff29c89b3d1a34ff6b9a500a95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h43310e00faa605da87f2e8dc6830c56d540e09786b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd7d3e6fb6701a05015a63ebdf28b161fd0f285c1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c201fecaa5363a86b46b9dd0ec9ea734ddc5348376;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3982b6ab36f30f979e109544d1d9a3bf34aa58b4fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc4f1b2d5ce64ce1cca0a17611003806b371c714f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha82bbd4e10ee7a64cd63fde88f72227f92c34b0e65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b7d713427df1cc1a650298bf7329f11ce1c812c9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c140deccfbac418ab8f2105a39a3274d0d9019a3d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d7fcc2700ba9aa0c172e14b5bdb21f780d34e0c74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdad788ac32789cd1384c9740199f4ff3f8107f28a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae22948c36ffca5ba1872eb31ccaa2db2d944919b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef537d15c62df3e9aaaa410af840407e403e096c6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cadfc02780df77039d6c91b2173c640f776d1957bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9ddb04dd37b91d5248df71e530f19421b7e40bd82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc3353e77b8453363240adba21d19ca6d75ae43164;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h905e8a3c6099c58413cc4eff5c2301c12c69c98757;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5937ea204c22ad49adf3c55757210299925a521fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cb837434755946e491aa7cd567dc1c8946b3dc5a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h805e0340ec912f618cce5178efbf4322304a06a4df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19123ab347b48a9f5cd0c5e9ddfcb61b9db42bdde72;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h284ba99080ae494ebe2d5d1300ce880462d5983435;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha127626d8f222bc6ad57fa8a12f5688e496fd14c69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb62ac3af4a246571ea729614b2ab895e7a7289b04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f2d7d3c30b31f79d22f07cdf9bbac1430f3ad415d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7cab26ca55115ff5674e338e0e5d22f691baa647f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9580d0d6aa85b88c8d4ce8381589689e26067bf39f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b64e355c7f6db9ecbf4056439e55506073d0ac791;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb80a57d100d5c14a8c82921014d75abb6ab231f8a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e70112a083096b3418b4f687edc73735ae1f3436de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15057dc0f9e8aa820e48c1d893b1945c0e01ef33eeb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h480fabf48dc98fec716a66e90f217f5a3ce49d4b06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e090809382835ce17cd22c0b2926f3a22ce4d7c1fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8316b0040943d6afb613985d1a110af2a7dfb3a2ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h196f9c3c665b25db80ec9e92bd0b45e63a9a46b909f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9c5bd05d3ffc32a531715f3a5994f452e0c93a11d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1365c723d43f0cce8b35a00263b495b415496fb5557;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53596ba06b7dbb0397308489927807cac47dc336d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195cd56ced6d7757fac910a23efb84093d673e9ea1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d95c4fbf47030a6ca44bbcca159860587365bc088a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3b877da0cce76425e339b7a46c7344cf7c0df578c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb773a45fb8284c70f2c406700fb7858153da1190aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126ca95a628c006830fdb8af7d97fd32dd6faae30f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e384bb5690a173d2b97bb3e2fa678a1e965a07280;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6f7a61e92e47fd45b8abefd6dcaed58d3dde2748d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h905bd07174e9039139ee3dbad32c452569d1982ee7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1190de14174027aa0249458aef0fce87e17d53190a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16daa1e346e335dea567201bacbb09bb39165aaec46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf66b9862b88d1b9d5c25b2380f19cd6efe13c78719;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101e6ce0e9b4460173e115ffb1205b7a447daf1aa91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6677c5ff37c7d2f2b7f82274c6195cb0d1f42a064;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8a51582f6e3f2121ae072926fa59f3fa499f3c5da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4327e579ccc9b9bcb770920292605a793bb1403a40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefeb074dfd88d725dd050b148389917f1da88f2f16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172716f7128e474db5be90c353677c5bbc81521db85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf4b2cc80dee069c1c6870a416bcb1335f54bb9ab4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef561cfb53e653f7c016b3cce5465a270880d98144;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d2811377bd532fda04ad72599113a3521547cfdba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133c419534ba067a42a8c156f8ec8d707b2a7f09b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141e1bd421fd0ad457054cc33dd60ba0e02516ad3d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb98d7f25719f3920a20660296c46180a8b613d2029;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130413da5d6c01158c12890210c6141841c22ac9ee9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcb21606c719d84ccc9133b2b7065f40c91761bd21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54a763425b8c95e9cc209627905214eb6dc7561014;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b33ec423652b3c7e5e03154a402fa5e13060ffd45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd474a3a5e5231de7ba4471b705e97fc9dfc3ab3f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e1a593153b6fd635301c17fc7a0262a0b1259981b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c1e20313475821afba909836434a1312660194466;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24988cd47453418251feeac17c7352a87b9651a5a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e7884689ae879bb8da769d9041ea36857593c4886;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4d9cfc9ab03fcaf15aebe0c65eb0bc37058e6bca6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5b43350edf89a6b4d2e8b6908a530d5d084bedc98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146cd90742d9d697cce6232985fe4de054d37fafae8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102e49263ac3861ceaf2a1b123167940063d9d20954;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbdebc57b5319f3d16193619a3a5dfc403ea1311fb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6847e53b9ce3411ec508b63fc43fb685cbc37de74e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf583a0eb864dcd296b23f01d2f8f08a100cef0318b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bdc88d340993761c071db45f2641a85d310cc7086;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a692d55ec74b026661df8fa56234646943ce688333;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d686ebf183f54774b2266527a38b0d567c3b0da6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17542b965727363abc154eefb9b74e766fb8d71615e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h836968508a23e3c361e57b05b7da2ef67cad86e99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2928f91db14f2c5d83822c7b2de7fd4ae4ce3008e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6d19b0b92da1a1497e51b0987057d7f14dc08aad8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f7064abc1bc9fbabf2819bb448414ac5c8a1dc3b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58fda057525f3302410f1285021d6b7faddb7327ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1f7cfd3b8cddbbe357c7a51de3d21ece78daf38c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140c2eab8cc5b61705118fcc2dc7ea98543fd15e898;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73c298343400260df1ac4fe040e2edbd0f1cff5edf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6b5ad8032010fc98444ca549b88942dcc1ff398cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8234816701cd52794fbab235e3c62f29be73961553;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h98f2232b87f86aea76107ac14f25712386c2c7a86d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d44a217d42861166e80f475ed6d16548d42297f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha9f51c96df1adae98456fd23c57b727bfbb2d4d17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1e748a771ad8404ed9d0f4b8fe7f0d94369bd2890;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5910828236490ea6712470ea7716b744caecb1ffcb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18973287b1c8af4ca56b835aec389525f1f31694aa6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aac6fdc38fba0d3ce189cc5c92c8521958dad8eacb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113344040a392e1571cbf5c7897922c144456ff7032;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106e92c9b005dcc14dd82c97dd80c9dfc3b9f13b45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c5b733bc07683aa01cb4aa3829609fd8e27fa256e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16414c5f6e1990d7bb234295e5b2fe17967b21b4633;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9c836a62a4c97d0376ce637ece985bf98d6a8fee7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3df20fb46394f73e1d32d391a0e595aac2741bdaa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd63e722f63d5447d2e533ec87cb63b6cccce60fd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21182e731a8a82c8c97c2644b9b27d7ea2ac7e2cd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165ba3a6da37b843ea8e9e4584d0bb68fa36a4b4b8e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h340d873348440257fc9b8493d9851413b1bd1d9113;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20f14c6ac8932d179b6b96bb0f5ebb23f7c6159dcc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16708d778eac800b042acb648ada6a840654071f208;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19123bb49183d28dc576e99f56b6caf8557d4b63b12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15784a824c7201f3958649eac7acd3589aeec144af3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha28ec12e2d04164f4e0d91f07c8a5299e5f695fd7c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89db733f3c48c860856a0a1d9469390825f54936af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd86fef26460c19e9b6a4f5eba654282e8db2bfc4a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16120bccc3f5dba79bfb160c3d5e3ff9c385fc6bb02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5b7cb05835d1364df9b0ccb0b5b9f164128a3990c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91588b7dd45971aeb179b095005c9dc95f4f30b551;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc0baf07a112967bbed2054f69f5fc45a9f0ce4be5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0cd7feaece595ae6eac3d7b1009446d5e704e8e35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1611f03a9682e3b7beb2a29332ec03ad63fb023f41c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9f18b9320bb993b64153439539ac7657ee053fccb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c89c4ea1fbdd804c214b9157b231ee55bae3ee9eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9861feab3977952eab74bd8f428dc5a248537ed401;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1803d9c994bd88790a9ab62899082a7cf05345e010c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b20aec11e024c79ede3b650e299a3511929ae8068;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32317455b48be18c0f3e3eb288f1aa11ed9d0946e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128c6d32a4d975869644fd2f83b54ecaf246d16e87a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14bc071b01f8326ad66daf9ae792404aab94ffd3b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a08956b010194ecf61df7af2ee39506d8ee7625d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aeb5dfd33983789c0ac71d4d83ac828d1cbcbe9399;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19234fa7ffab45c4b4decfa791bd4461e89e34b808c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6129116d485061e9dfc44bddc4458d7bfa8608c0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123d43559aad3ec73e4828341ab7bef85a9c54e3994;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140fb7e07e254f10392ced3a36e49775118f483f206;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87abc005e727f488639ffa611556d39ba64afd0ff9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcba58243ea9d42947113b41cbe09dd9aa10cd7f6e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff005b226535b42a5c9b4a15c9291c5ffd222f2ab5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b3335f81a29802e0bcd39edae0ec445359ed0aab3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c3ce81a5e6bd2df51012bb8577ac354d200d5a128;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1120508afae5e7ec12ac22b61c29e4bd544b1853a68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52be3a31a0f53d61be9c813e76bdbcfb7fae355326;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1e5f8ce64ed7999f450b481949af56305b373e08b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1165317412b5878488ed3b1c8ee5c76d60aa6a1d0ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172c0875b803d2a9dc926e2fde3d50e8062a95b704b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cef6a144e2005566fe8dec97b3cb344f7621c4b5af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110c634921c7ef202c58afc2277c9a87829bd7f97ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6473e7a5e6fce7cd6be020440fab961076cbbf00b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c65ea872bc8df232cb5e3bec893060285c60620ba1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa2b7a1d0c8cdf9e11f3e67c274eed18d6c174cebd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111d306ec6e40c30cc6c939119760d8eb73b8ba3bc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144a2b68756b77de8951ed6493f9358bea7621895c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12053641c2204671d49134f6a552a650d3af5da1d00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b1e0af0d99bac3e36850d97cb20dbe4fa89310073;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed6617af52eb53db9bc9c3529e1c046eab8ffdd16b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h151702dbfa437d85b8f708f5a01c36cd4c163293449;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d835af0cca5de1f09d05634fb734e0acd1583a57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h139cface7f110ec4fc6bb6d2c69860ba8bce09f7fde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h357895e0a48ac145ba661eba70436236f0421c381f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h204a3e53b7e1e2d33f1d5c8b20f9890cf43017872e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122e9eafab2caf6498ea006bfc7bf6f201192940186;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce1491989cdf329156ed097ebba19bc50f6050c8f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b851e2d448901bf391297a1272842d64cf2ff8185;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35e6968859e32e13f38b14bbcfc98654320e4cf202;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb94e3a9e4394343b976929587ae6b2b574f9310fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef3e9a18c471877974da72e1c867af99e7c7593689;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162f614120dfe86429acd910d400f6e639658a9ef23;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb12b9e092c00830ece33b51c710b86222f05597c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h311ecac906f72f3c3a0582afa0aadd025a8b583073;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1adf6b93eb9f8ee425eba77328fa4675757bab83d95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h881f614c11c791fd786303055fabad6e60898b4c61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6292206a3fdb68a7894e50fd28e1aeb865a872d03a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbb019f33c449a555e90c6dee0ae4b063f8c74ded3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hddbc2b3c63fb3fb14c2f5a9ac1fcaf18504e1832dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a63cde5f69b564c143e03481a1a7817855e35aa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e4ad58ca201f48a53c6d46e07f12800947afb2874;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10006026f8caa0a3e22cf2f3eda43d70fcdcba271c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e44ba925cb04fb595ef73f07667dc0d4adad1439c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c54e85bf5abf3de12be7153f954ad232422513a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6076a87237c3d76830dc1a9440fe753db6149e0794;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127822a1f0493011238f50bfd69ae305c227502a972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfde307a73cb5bfb13dfc691c7a57a4bca1cb5fac9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e76e4ca5c1832402ffddd657e9777a8babbef123af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e45a6282a05b459f93ff9242d99659db683e8d6a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha169b07c181fbd27f136d743dd1ba91a94d3750567;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53f48c32f2fdc7d9cf0f93d03ee98730a1f09d2f05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac7723a5bd04672f30955e9f22b5b3bc86f93e80af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3f27e5bf92735e6ba4030718998e79968742b5208;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af02cfdb1128064aaaef0199f9cd86a6851d82b18e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd40a263ba40dc025752044c5fc226299c007dfddc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h49f5b2fd92d538ce4423dfecc21453fa843e30c044;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fca4e23f010ae7a3a5b26f4274a7ce103f77ed9fb7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc89ec19ceeb98bd4531a1dfa12c718cf3e4a8fa88a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb94c1287d42efb527fbd7d95fc9ee42426d8f0a620;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19441adffd1eab447b27f02231037df6444254fe2c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178fa569d378ae85a064c7850d6078f99388bf8de0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14109051deae99477ac49cbff2ddb4c65037cc24de6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h929ff679e928dad0f71b8dca33e26a47eda9fe4f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e23593fd37bb4fab9fb1c26bf7674ef9b12e0a1a74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f54116290213b5a246a426d658e6c8e1c8ed03283;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185d8ca568795881e6c91f85c7bb5ef33a01c7efae3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd65f0ce884feb99fb82cc0864d02a2ef8dd4a4dae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2375da1c820f98904913bba9c88aaa08716a622953;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edc65508388c37f2bf595460985b30709026a1299d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8926770fa10e1b2a1f80380f881093e3182fb702dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f4d87d7e861ec10d0116e4cc0c0ee4fe261fe8177;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135fcfb0e23c8082f517651554d3da79e697c178d5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152baf915def88ca4df7d3d51ea1d89b6673c1492c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d5c2d4be6a4e59e931fcaafb1f443da38c2ae76dc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d6f84fa55c397f3eb1001c00cf7da2d2cc1667908;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7fa281c60a9b7abd37ad980385402ded40a073e05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1079cd3b12adf42f6ac093d97582978d3add51a52cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1837437cb610c5d345faeebdb65ce8ee549bd74170b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f13be254700ddbeaefc54409879bfa8f7da42fb52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0ad883c57c3c18ccb7030dfac9d59536fb7b3bd5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e615782ea3e670765318becff658861454919e559b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118a6356df718331365f320460bdf9b002a1f124c78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8beeb595ecdc561feb5950aad6c7aa22503296e5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166ec033b1d2c8e3097f8ad13808256036ab3fdc476;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f892aa5c7bc8eb3f4c36da2ead645bd3dd252d3286;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aee7716107cde4877e9d0a8c021949b1f7f6bfa9a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf439b602f0cf70022c8beadc2f42d10c1a8c60e771;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h136c27ef23dd8901f8cf0ca01c1651a50907e158c95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hadb9089bf1fc6064e6ae4e8c85c3ae15302f42b6a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefefb49fde529b1990a8a2a471ac51790f9c4a81f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h429c1ff5fa244778e9ca9e4963556c7986d5add331;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57332c267ae22be7efcb23c6b089f9ffa677d8bf51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87f95ee64a90438544201b09e79ccefc0625677d4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66660e110b8a03ec4f5fc836c833e1cb360f91d363;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d66daf1944af0150927c2a9c63acaf633777179c5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1137945f7eee4c88705c71e2f8bdec37f7f0514122c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199c08d99380c51576a73a07019cc4ed95afa583cdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17300baae47619086b01e76c924eb43a69d7d8f77e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89ab40e57e0e727e9539bf95ed0ad03d843a9b6571;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44eebc8d115e165619ddbca7bfff468a75c2800d8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19300cb12e8f5783b78ccdd68355d379ed0d84543a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8c2513ed42a50557ba0f6e491a9ae487a39513fd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ab30a697837a50ba5437bd00095c6901ed2510803;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he87a6e72f9a0647c156a9483723df6aab82b15f0a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h625daddffd822f4f7fa254ae797fe5d978df7dc031;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19476aa56d1263c2194dec62b924db2a8867662ae63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b635e9acf2b736c9796d815706bff941a19a639a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc244db3c719dc7aceaa84979d82948dba3ddd80e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ea9225bde3eacd3e29453244ddb96d3e364d5138a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc8af95376137b28c32f95147232c6c10e22bd58ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3aae2c4fa9424b0eafe0584af6f50b1c54012c121;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78b90230196bca79b184c1a528d897eae3071bc917;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h342b9f0ab87722ff1cbf3e574217d36da85a0238d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h670634f8a023eb272ecb4abcda170c8a4e7f2a60ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bc189e98956a89faa6a62b09201a4ad43cb2d39ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17cbe1092bad676a5d7af95bb8c2ebc36ba6ed0fc19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6f10794885606a8bcd553c57d24bf2a0c523bb629;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f123e601f953985e521469e63085a27ea57dfeb9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190c0629e941a60b446cfd4fc3a2ee10a5bf241c82b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc9647d790729b663e2ab46ea82f959399c815a639;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e74bcb255d70e7e63e379a2459596158731ecafe6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4521273f7c6272741ed5f3441d38cd723dbab3464;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hceef90dce7187c40e60ede1e96a0233d075924268a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9bb2ababe4a6e1012e5648bbb8d6ca013c51641631;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174cc0a0081011aed5115b863b1f1b82d45740b9c5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1077ace0e872327ea221b60c1fb1236f0873aeeb10f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c9a053cce272322155e19836b145597f916b42e3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b37450f0b305e7740322f95198b1e1ed64b36f315;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13aae045f69f63d71da4af1fd96dd79af55a4d95db6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdff1eb63e4400225e8f9f178c15d29743d25e09729;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eafe43d938e838c9ee92bb1557965da5304924e83d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11204bb09af3a9be1b2d7224469b1aae43105db40f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd29eb01396a37a1a7edfc06fd9330de21b9be499d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5796d5ff73ef78d7fede719b9d25a53d339de8b698;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8752ea02aabd50008abc44158306ba262db4a9757;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfb7e728751d22bf869363a0514b3b85094c4e05f35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48093dba722e3d84307221351ffd7526c9d1aff036;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9476fc0216f5040b00d82e2c369409c4d96f8a32cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7c2bd045ddebb8213e08e065fac9ca124df7d940d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14dff4c6020224069ffc77e7aa896688c5c98deb602;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfae38cb85dabd776a5f1cd9f68fe4d3cf8e8a45d3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a0736851e1acb8147e5b76d0797403b5256b70b8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b72a70fc7976d5b02e21eb8f9a5efe85cc3921d858;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h522fc51754b557808cb74510e059543c77f5b59da0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a42bad2168a80eeccf5471d373141ab55c4c1924;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3ec970783cecdc34a3186bd07513de174a0512556;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f35c79393625d77f983c497f17dda62f73eb29645f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc956f93084dc8efd0f4cb364257106ee691aff0c12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148b486eae0a06c29c24b06b2349a3f3bb7089135b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f3f6382a4f87bd9fb7aa0c0949a8b4c74cb9835f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf51c31842ae9567045505d1ab8c5c30b33b528a143;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1145ca5c325321ed780c97e4beddcbd3c9b84a9492d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4a990f4870da144fbb67cbca6ad39a685e5dc20eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7f5102a510deded17abcf9e8f71cfba91ea2fea612;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ecbf581ec9193c48c728d0b0f7e1570465219a31b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177425432043deee8f3726982df82e2770c5be6a892;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c207f609241d5ac01f362ecfd9bb8b956a82bb0c62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1708d6b4a9614d0e704f65e5cdfecc1b70b2fbc7549;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9161a2638aa2b5beb06b17914ea43ba3f716a931d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1733b6893a0a875415b4b9b58fd90bb69956e275c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24882ae557fb04a138ac312e90732590e0c89072ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcdf332231579e427033963e209becd4eb101bfd3a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143c0ba85cf127a53ffb3d2d37919063c22c56bd914;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24f5cbb127752884fa66752689dc9836b4d4a23719;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182895a59fba4df30b0f2c8daf51af0f5dcb0483474;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7263abd8beff6b3d48f29ec914b4046eb15660655a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4216d410c3806c9b80f3b49e0d0000414ccb87906b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde3f7b713c3da6e2bd5af04b110fa58f736f83f4bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1659b4998b05c2457e2bcb9a22f99ae96c57bcd6971;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d63680704bd1b5842291d4a2e3857f8d74b6e8954;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b30dc7ace196ddb985a30434828c50fe3cd050de5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3019512ae286c621e8dacf1cbfaf13c723a6abcbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aaa208082dc2f9469ea62325abfca6f7bb3d3f1c7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31c470c8adf0ac92b9b96a25479e72966cba659da2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16b3352489f25878de75a32b7af5e23cee60c6e61af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3f910692648de3136473e1c7a382f0f417fb5a016;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1361202208abf4b01ba1292190db54ebc0d9328dbea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee5e1deca494a97b38bb052fa51041a8afa58c3d0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66e3f2bb41861f133f333ba348589f1d9910a2139;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44c6005d9c0e3a16d48d22c5ad0f69c002e1d36c6e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7853fcca9f4e5de215c0c464daf4ac372d37ac46f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac349a5ead2e4087cefc9904e9faeb550cff268623;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3497e14980e642bd4998532634f1db8a9e3eb367d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f466c76ef83e0993fd1697ea5f9a9e41f7d53117ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138fce92d7d5504730ef605cf6d84530ec692f095da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h438a2aec33902d01637da1248bdb2087aaab2e4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158afcb53c2a0f721240808d0e4c0dc06c6ef2dfe9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15899496106e8a8d2ffebf6f570c0a5f47222e91f98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17afb624f57f8689bc4bb3a02c62b268ba6d2ae105;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca4c1ac7116435da3fab8813771aa35dfad52a69f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f6159fe77eb259fd161894112b48efeb0d09475ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d0c75a11308ac34672ce5b9172b7306d436e210d17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41c8ed8b3cdee68b02cc4500ebd734f46d71f57aad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ea13314ffd5fc9c61eebe39a38bd6b6d91b7c28b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb054740d071b001f6394d9581a8fd962badb82393f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ffaf95a68603540e10cb8f03c19ab34c9d3da7bc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h136d80b37d77910479f300db518540f30bb4208ff51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185db7be4f2a81a350f437513c7437320ca040d04cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26bc5147c3a405353ab0f5de2b898fa8ccbd9ecbd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1060d0b270bc8b76cfab39fbbc378c3d11e0d6e9d7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ed3007af8e4880e5a5eec7c65ad2351d991140f111;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16eafd01643d3dbc2c8f4a86ca53642124ffcd63bf0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1418ac3c79a52e6efaaed3593eab375f8d555736fdf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb308156e6cd6ac16225083e2044ff0bf1b7ebb1cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6048f59d282bc409ff459d0c0aaa8ea62c5abd228;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14022a677f71b999155281b93af1ead399ec091f195;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he86ace774a12a48c879a1ebd2e5e0d52b2b16c711e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea92836d3889a37fa958e947b85f6df8a479a26bdb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a0e9be6cd0e99a7fcba9ff59b836e5262e43f4e42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1827f7b681abffbf559f13b8828c8bfd954f594f815;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heca61f5f06c01175fe1ec2bd00bcb406ff0d9faf1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1946236e4b3b7e613fa3649f77c8dcc1ff9438fa13e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4223ca045309b13c5554822c5b1feca05d2f76fb91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7e9a27c7d14458491c60bde42bf26c2993e711189;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8adc55b0a0e7706ed975a450e8342bcf979e91f83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1416ffbc818923b30be29db0188f781e913ecbdba82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h846b3022d542cfe184b4dcd9587384869cc2b9fb77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4555020597fbeca89cad8ec33aa4f767de7c8c144;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138507d6fc20513dad0a3a3c54f013c85ec97b766e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f63c0f23df83ff770215b0045d1ca767fe40cc2124;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17638e75d9e053c87dccc361249388997fbd3c7b739;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8bcfe10117242b6143250d285cdf7500015be33ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h129dab714436ea0e95a701fc79bcdde9dedb0814c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f37023f372fa3dfb040517f36a721bc857d445475b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32a50482763a0f1087b0835e58b27e3bd40043c7d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0be00f0621b754e7f66e085a83620610f115dd3a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92d2cb650b42b641de63b8ecfcb6152888a0bea43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2ca74bad3264ed0ba11eb3b6ea9994eb7978ebe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e831a5e5f8a59fb9a12cc810e5decae730460cadbd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194041f73b31f33134c8e4ec4ef9bc7f0c377ddd57f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131c5dbb62f58fbcd2172fc1db6cca2ef7b0148f56e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c695d008aafc63bee7bcfb5e910d8166210354b4fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8548bec285e00d8e8e32b531a64ae902b33fe077f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38f1dd44e84b2397dd66ccf950be0a74bdf19ab2f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a48fc2035ce536baa0ac76d46a3c3e3d1059d8760;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64d365adb252a7294972c68364104776ae9c74d68d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1167d6adc21c50e6ee5ebb3e65b83a72894f44f7100;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9fd2eee88a9294da296f17890ee2f1f44a93cf4b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1859236c342c89b2eec8d887f7f729683a43223feae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he56dba082b7d251693de83689b0acd49095c7ea6f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1feda0d67f77ef76060a363a91604b53ce6e634dee3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63f12ab8c556b192dc1e8890b441410702441e184f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7df5f1f19c6548d4d00641a3160206ef450437d7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4becb4d7af774d592319ed1395a74744a26382095;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97ac481c9ff25955c1a7b93c339370f127694ad074;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb3b13f8ca8e152f1ab144eb564ac4e29b0f931f927;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf3aec173064d5fb8655623b5a0cf742746645cb60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb074fbfbd00edf5b77d74e8abb49c986bdca3dd806;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131acfdba47fe2a8dabfda70f4d6038358a6fc6b821;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0e449d77f49e941568dc15f384e4a7042151b21fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dda6b2a91211a5a08d7e6c4c075fada8a317835306;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf149d3a12b0e46bdd512b469a8506cfaaee478d667;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15221294daf2583d17dedc137f3ce24f8fc35fc43c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2808ab48ab92c135bf7cd55334ceeda6d6d8614de1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafc561e3b2da0c8e70cebbe9c99fef0e31d5024a14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187b75f1ffb031ac7ff7ebfb95e86e9b190b7da9a79;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ff180ab99111bfd2f2d1a7fa591f543ad7048177;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100df8de312bd3affb383c45fb79dfb1c62d54e29d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h67d0084aa9e84821f66b4f9b07e68d47c40e7c7d92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47a30b00dfb48bc9ac9d63eecf233e9af280ca0228;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ea909591b843853d6216d3c4b9047e7cc5588bda2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h46a7284cfcf6a0b034d8de8627e19440bdf14ad64e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab3a2b2791a6f00fec12612f58c3e14446f9d93080;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8aad43f5db917c740c63bf40816ab333dfcf0172ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3ad96e0a798cc6fa0b9eb3213025a1309068c8aeb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7ea7179da82adc636020faf0fe0636ea5f8677a2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161d9708bfc720bbc1e8419f61c906a619e8edcf000;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd60d0af92f8e867f37ca2ae12d93a790cf6c60eff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5db89e904600c7a6c32fd186fdcde23a3c13f9798;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18420e41507057fab90c4211ce48ef0e569b9ec3881;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1360d9968d023145607eedc5d860af310862134aaa3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca8e11be343bbe2cc6ff01f3734af8e7be674c88e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e144753bfbffa3f2c315001901b6494509e7fd2962;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1c10d311615626aa8f4b91e50c27f959d9785d696;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dce6a9f63b14b5c9ef913ee0015ef37d397d6c1f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6a2606d3278c7d9e6abcb7f16a8a0418c65cf7d25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cd961c0089b796a849a1c35a2d849e27ddf454c17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89137be3ccfb74253c71e4352dd0f7b789c4007bc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b1a5e0966bfa259c4cf61da7e09bde05e37885466;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c95455869ac5fa3b1adaefeae1a580e06e3b1307;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd06e06513ad9baa6fa1f4353034ac8848a2c2b3feb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8637194fce6bea08bd7082edec562ba7dfe66f4871;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c60677dd308747c8102909dad302b7691923de01ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10546cb9eb140753b46a5e7f48ab91540d6294fcaa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16670407f0b0ad8c02da4680d26fe641d9b509ab9cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7bf360d6ccb8a2030eac1821098b0ac50d715bb8cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17469a2e7d8f1c0adb8506b6d5666a9593f653e92b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h88a511a4b3aca7e25667b66a7d1fad3934715f3b7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e65781331a3ef4e3960f0925255299fa8ee8dfefd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb113cf4dde9ca9fb7d2de8c493e82bef5a984dc78c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8f8994f29b22640c3d0ea31cc3e1b38c75da77521;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h136156478f9d083358635de80b819df600e2fff4640;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafe8bd6cdcd619dac934ae53afe5acab965ae2e696;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3119f6f55eca7abd065da7db139a5a08183f8c8db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3072905dcaf6f80cc2edd388646972f703e0c5cd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d5736bf040fe9f46ae8991ee91b91bcf99d6199f83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5ab17ff56ca6ceffd9e066aeae21eb7bb9a74036b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1907fad27db927de443373b9fa84cc56b35035a64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd2366349fbec324fe5680212d2c19cec701efe181;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6492da7b3bf8176d71290233cb07073f441a2e7d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e54b247396abcb5af23d5a8d0642e7a0e8f0a55fb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e23c0e2411da78595349f09ee047678133b3c8458c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecad2c82c9faa10db60f442fb041e628a7736f47ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h944c20f4a210d289cdcbf14a7310942e60ffeecc98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c179a72c6de4fe2ad71812cf498268b31f426cba6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3fde9129095e2b6ca27ddc9b63671593c8bfc161c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c17745b98c3530ac7b91b4c6951d911c716046f88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h626375fc6994ea65c87baf513f0bc24b97543929cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3feb5995703a2fcbfb0e73fc5c349d49f65534b38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4da335ad5007a51b1e70f7ad0688f9c603c55e9b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45ca7efb9be478aacdd3aef91a0cd8b32adb168777;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158856cd174e5a5e5e353ae9ba9741a9633a09b0424;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f5fcbaa1e8c7b461b2f24d24a44fbd7b0d5fe32e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f84b1343a9f596bf8750be0ebb9f6e6cfd0dc2cda2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h969bdda71754b95aeeb65b16f027babf3d32620614;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d944011afa72d1d56557f1e6c7bec0b2f303b8e56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h997459f7122a82001cd0a40b540856f2d03216d9ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1036624424e6c432c29d1e9f7e8ccfee503db8868c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h275e4132d733100fdbfd655ab9990a8a49ad9422c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6d9fc90872f7e3adf8cf0db79e56dcb773ac6351d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bcf6fab17c2c353b8478fa4a798196bd2a177e9b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1483fe42e3cbaf5b3f8cfb2e1dccec378456c326274;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef6235ab73993c43f47bccaf4c6a9d1d6b7377c934;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e1c5ae7336e770487bd744c15d845a649ac1fc28a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcaa33b15031a927c5c8930b6a62f384b04f0f1379c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefb2604ec45d8af6ee141cdf3185fd7b9f7f75e344;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157cce4d8f955fa0d9b26f0f7e9b8c0920081bd20b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc84e86c1ff18596ad23074feba2f36fdf3a2b7bf89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h880b91664de20bea93f21a267965dc5c925a676ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6c1f01e8ba99387f219de02e8a9c1abddd4dbae27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha24b1ae067912140345c7fdfc8c50c6d5b4e55c5a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ef7d72076bf7d08152caf74f399fc6d8b6b8d7ba5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58d3bf0f3e98fd668287345d8e4b72df55fa646440;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ced956423e36aa9847620ce7120ec5e3b46f41529;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b090bbae6599b597adfda08a123db38810130addd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7216a4a8040178e9e7f615ac3056c0bc83eff11159;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e9701becc9e1789fb595ce5225ee8f8cda4c16d68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc91788d0992d5a0f69e341c71183abf41ca3da7a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b34d67cb7e9d904b82a7d380f8c941005a2ef3065a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc2ee3332bce567d39d6f304ce02baa0d97b07a070a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h432fea68710525ade03c64d62c0afbb2dd85c906ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80a799779b796abf7ccec46eee376a51c319fca4b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4d55b51c8065b4d01631195ef89c2683c6036ebb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fb1dad73266f4716290fb71caf88eb28afdcb98d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b952a16e86e914fc92d0ca34725d76a8e8e9f57e3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h60dd3d59867c4c5eb89168f04f53f492688f940670;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e4d8a799ddfdeabdb37e5f842d09c4e010d18aa9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b0182f361a8bd4a994db2c40a20adcb69bd7b784d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc99200e4c2cd78e2c5e9b08a74d83a485aa65b1156;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3128c0f15a300e960baea26960c6ddbbb7508700b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33ecfacf8e4d276a895bac2e87335811bcfc520a19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1fdfedd2ed44af68f4328966d8bfb785af5c13d43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32a374deaa5f5ef26137ad575cf34c12e84cf348df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf189ea8cd3635e2dd215529c19e99d9767b6d71d15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53df8d99e2d1e00ed0de4704d18fd920304371bdf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92c61a38dbbf65f53bbe5a6a8e56df8cce42b72b5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae41038e6c80bc8ca2de2e68b85815c19126966607;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f2c9042ebee6bbaa5f3ff9c0b88057357180844b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1611af714e455cc582ef7872fcf4822898e137fec4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68f7a71cc47db1585013def3ee5e2cde40651d5098;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70e6e1ee5a7c20779cab50782239813ded59e1726;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57b20da5d36084695adb350926e6c5fe0a9de3180e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176376713eb72b05dbe4531f2c24c0cc3231666387c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h423679a557a5359ce80f47830422952ff48021d214;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h589ad5dfeb7876505faa28783a5c59083b27d41b21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180ea3917512d0e33232572c3475c265d01709e8003;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16799400a10a7026188c0ffa4206af9e48073b72e93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4652609726a3aa428d1a5884a0047c676236101007;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117478bd49faa5889792176ebb7cabc94deae8c984c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b6f81f45a76f6650f480e14784556657e192b37b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5f1a776269e8a7105ecfbc989abacbb26565af9c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f5233aa92fa869c79773bd4bae64af887ba6a8ac5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb94a0645862e08a1b01f6d53ffbb3aa2aa8f70bd8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2eb31862e27306b5042889fbf42c82f1d699acce7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94698b027dcb7e2fae94abc058158e2a35e4334a31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe59c57f9049c52af57cb5605dac21d6fad6c20d69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74bb69a6dde3e50ef790d9ade73ef04e981f251132;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165015a9e5dfe46d1e5f6cc3f73cd6c0681b4d027d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1020d136f603cf3ba430c1109ac9dab939f2329560;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf9521b9d29e5b956257f6f77d9bec0c551fa5ea93a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154bc5bb236d5c051a396029f3b00e22dd48aa160e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be7a126037163aeb142478e8138a34b72b94d2fc6e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha161394604eebbc0c83f402cfa2f18629abc31930b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he48c2c56fc6b91b99c7616f0d7c46a0995608bb89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8652d4044e0370c95d39222662acedd35eaf4ccb26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8413a78aadb0847ef1b7a6e650cbaff61f2468c302;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195fcabea541964df80bcb035b77da76e17299ad272;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f5eb2a19e0fdf32c90dda434134a2c9d2c90d5ecf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44752b4263af69c5e1bc3331dd924f56b806114ef0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ea306618684ef342cb2c93257de5eaafd5b95d03b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h870ed4cf1f3605f52b1f7d3359178bdf824f8d6c95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h84a627d8103ca05389ba47ad19877796093f6430a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2022b1d04ebf199395ac793d32d62104690203cf27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10734ba68aecb051fe37ae37534ff4ec442857c4d38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h623eb9680a780cacaada4bf9490214d5bf1a3ea808;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf23f8c88effc24dcea4cc79fa3704aab7cc799d89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f21277ec6f9757ce7538ba5e25c21eef9f44ff9ef8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb90f2b6a4254499f9d62b660ffa88eda3ebcd2333d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafd064b18ed8d39db860e6b72be1de517d6a9546f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac7458c5c93313945063a853a11bf2b8c039acf058;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1663b60abd90fb36591118f4ae1e4f87b5d169e6f08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15023f41fd45fc541355d53f79a962eb78e0906776e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162ade34bb307517695fc63e4cd9e096c2955724fbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4fe16f6c81c62d7e1d993475bd062e37ec55d0b5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5cc843cff0c9fe38068ef16d2bdbc303559aafbdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19dcc3d84d5d7ed1d9c0e253802ddc11a7652c1e16e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd58d3d63615a21a182b61a7090246349e08f4c382e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155d1c5e1692c4f8e82075be2dc46a3531d8aadff89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h368e467b7d4aaa081c568399d8ef206726022bcdf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168ef3773b8fb90c1e20d65f01ddf3d1469c5f2da32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8603cc667fe21b539c698c1ddf40003a7424a5534;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f90cb6bf847465406d45fb36b8768c05aacbdd54c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd031b379db1a1a4acf478654563c62f297f7586e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8aa77f82ff31dc4983eec24a9d84f124957b3f9a41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172327b771c7fe3e1fd59d52d008fbf62cfa431ac6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a80143a918a93dff8c5d8b96f767c59b6633490c41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h79e707b4dc1548496a7eafa5acb79f477e322dab11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b99450ccd0c95683560cace4a0d79551910065bd76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f53bc98d2c664f9f10779eb9ff1bf4059fc98fbc64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h513bd495b12165deb8b47467b7fd63e56d0dcd78ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15fcd3ae02715c0d4cbd546652ef05624e5266d6a70;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b06da36671a3d19ab032f27ecb8fcc28d21dbe47f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b11523e7cb3d24f4d04b832c2f6b80ccdf677009a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8113e5413dc46e2b784afe58dc9ee68ff03e80a525;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108655da8aed947a74298fc31a3a8f6ef835818ac50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113cbc37c8a103a10e0e9c10e087bfa9d2a1e98d9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h394e3b038262a2e5f1fbf0526050848950a960c249;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80aaec78dc2c22197adbb84fde725f6a7a03c9e100;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd932a29f2094d88922d04321544e9c034b47f4b39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192376d0fc91a76e37066b1ea978341373add16ceee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2ab4839a8688bce502cacfab81424281f4dac8e60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2aef2df787e59cb14ba9b8b44505b233d2a524ce9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0841a1b9f0bd0562076b8f86ece21cc87f07b6c42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11b0226de735b6c70aa5b3445a204febb1b2f5eb0e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a9bc6a119736b918a87ed48f51ca0e14d49b5d25f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e430d06df18f5733a0abff2befe64da191b7571c32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8f5f60bf15ecb65fee4d431aac4209fb8fd276d17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d19f7cec0bbd6d5c1be305d4af2c72326b93f6ef85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef596422b45e5599c6a565a01a287bfff564dd4069;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce32a9bae1bd106f4aef2939138122270537631bec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e0c307b5139474c57a873020362c153295e18b868;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb7681b0bee985f931ec8a9537440e5ebf884fba58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c90ae7b004eeb07eca9f958f7416e139b09302ed4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57302913d433a16a6546859226808ec878d2440a28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a210c637f32bae01bcac5c904fe3f98812401af72;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be6e608a3e6bdedb10212e512067eaafdfd4025ecb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9701ef7f92ffb6875203958c408b737139756af519;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h795953279da95127e8a9149f85c8fa832e38a26d9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1187faee05a9034612b52e54bc0c341795432c7cd80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7dbeb71a660c6d89a7f3269c9d717a7ba50912c6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152b5e8b34e8a733551e24b56f48459252131a281a;
        #1
        $finish();
    end
endmodule
