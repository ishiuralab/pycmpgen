module testbench();
    reg [29:0] src0;
    reg [29:0] src1;
    reg [29:0] src2;
    reg [29:0] src3;
    reg [29:0] src4;
    reg [29:0] src5;
    reg [29:0] src6;
    reg [29:0] src7;
    reg [29:0] src8;
    reg [29:0] src9;
    reg [29:0] src10;
    reg [29:0] src11;
    reg [29:0] src12;
    reg [29:0] src13;
    reg [29:0] src14;
    reg [29:0] src15;
    reg [29:0] src16;
    reg [29:0] src17;
    reg [29:0] src18;
    reg [29:0] src19;
    reg [29:0] src20;
    reg [29:0] src21;
    reg [29:0] src22;
    reg [29:0] src23;
    reg [29:0] src24;
    reg [29:0] src25;
    reg [29:0] src26;
    reg [29:0] src27;
    reg [29:0] src28;
    reg [29:0] src29;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [34:0] srcsum;
    wire [34:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fb5a6b5ed328204c69b0b0cdba39a40e9eab61803b5e7c482d0a508168a7eee9a399f22ccdc36a9add1af2e7aa6d48dea9fe8ec68de526dfa54cd789b8499e9d0ea555ead65b9868d9df3982a5ee35c17ffecd68a0fc17713112a5e56669f805cf95ccd44f255fb72929d1ed477f14b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h696e145153ce08017c5cb2b0646e0f2e98142ea6e89903cbc09ec6a24207cb8575e925f33e77a60a143214f9b65ec0297e22c8414345246d984c71a119a9720618fabc1d57383cfd343642baea0470bdbdeccdfecfd065919d52b9f737edd7fb6574b079cce3a9f0a6f6ce280c7e9d286;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3dbc1c07f97f0e40ad1ec4b23dab4339ac8f9854c175bb628383dcee178fe924d579e144f9c9b0c4f7c05b45ffd415452f1a1c4c4eb64434e7660e9af177ba692b178c2a4cf4449c4ddc89c87e3ab878aa03f5f015178b29a272eccab6ef3e64acf7258fae75705d2e05f26aa79bd536;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf28db8acfb3bed1e9e1e5bf062464daef3170add245aa10f80cd896029f1ee34d62fb08a9bd8c03f3d7c73e998424e52d20742a30ae970efe439f74d2383b619f582bfbd575bf0a5ece043a60e1ed561f62dabf863a0c42b61bbfbe313a754ac3da592219cbde89055c34b8dd19a3c1a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c0e7728565c50a5395b289e4d91bc1c554ddf9654a64cf6e28bf6011ea135eb20e01a94eb277199cf61f4414f613d3959bb8206fecf7bda22d2e374b4b919c1bf1dadfbed4146bb368d9eb2d84ba8e52fff53d8a7a91df7527ee6a1edb145da2b208458cba5f0e6d1c22549c629e6033;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h533a619aaaaf3ed937db09fd17cc92b2295ec0f56232786b13312a3e8306e76912889a8b39840daef273757a3559334c4a83162ecfa2c0871843e3ff7bae325a728070d8d480ca8631b593d9a6d1e4486870fb5258267710162787037c07b21fe19c9b6e5143fdf69e8e2c06cb715f605;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa27e372ef88c774bf96a3e2a1e7838fd34cc1c3ab3bf87c49f4247e230bf570df6f0c622c0ac1a7e3d6507295ce76a66709e293358d39d464542964bf3171f0cecdab79f0e737b9a63ef3cc428618255b22b0b05008526e3696645a453318b8db57f47dd38c471a7665bd7415060c809;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf539ce19f7fd4deb0fa2b9382a543b54a6d9a4622d79be767370b63cb08fce8c808f1e79e023b41c57885bcd28e50ef1e7432cbc156754e0b7b81e2707126ac7b358c2a3b095ebb912527032401d538e164a40da419c784b80c854b7f34a125ba28b689ab07c4658a302bfe00ad2ff19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0f9ebcf596a13d1540f4d77ca5daa5776b35c81e15604e3703fe402b1a6d1d3fa2cdaeb1888c50418cfd342a2f4782b544f3d283320b81a05fb3eeb6f84db3f73ddd944176b3dd93b978a31fbab48e49e2e3bc494bfad56098a6d8b74e9df970c7ae143dedd008914069bdf90b0e62d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he22e023e1e7fd48eba8486785270f42b76be025ea123fddb7da46a5e9b7f310b2a0a3d543c2d99821ab95c97618053b7adb1d44442d2e8ba064e5e735eb93f4aa4bc4eef2fb1cf2aafa00dfee8c8195a3195439072af809df2ff47ef7edd7a3f550dc832bbfd8edb675e3666f04fedea4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha79841d860c07e0be69b0172f1a41a79677fff5803c841c1c01e3f50188cc8345bd32210f9fc868a57453f986fffbc7fe91c14b2d4ee54e29b45f6a72235e174c0e87baa6e9c4d0ee1274c7cd7a955c5e6c480d0712fdc0044316e5b3450d5e21c1314c570b08acd94cdf970adc2afd83;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb196bba102dadb32cc5de09079217626dd93b5d537214df223809701acea86f04304028e0cbbb7a350d19ab8dd787ded677f3e97460ec1ec5520368958920d0ce4dc17ccd9738fe829f8ee918bc9006c293f8a3de92815fb4a5fa85652e5c12b57adab21d922d2f376dc402d509d3efe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ed0efc71ade5d869a8b2acb515cdd6932eab7c0011f36499b40e894593a05701fd030eba70f4829d8ca0c809182dea22ce46b1b6192d99030d1c1fb3d15723c01b147c3c18ecd2c05a50bac291896b2aaba1a51819052a73ad5523da799159f4380e5d5525a3952e9c247cdf95403cc8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca021c0f2787f63a41ea5f9499ec8a57b6a3be686d92e9f45eec6feb41c2fc684f34fa1c1f97226d300b21bd3ab98fe65bd02e61c4cba808d1b568071a24ef96c9b40e0d36917fbc4e16936ec1e68eddccafaa0d36cd4c5700a5373195714c2896e68443d1497cf3644911a8b6021b2cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0f35fd2eb179876e2d1882ab84fb7111796ca47bbd0efd9cede2a912033d37ec4dd57e73887646d28d8ba1d5c2bca433d1ef25820e8ae245d5f13c65ab9ba967cd803da3dc5c65beed6e4c6c15a934908efdbe12003936f3139756a7b9c93d48ee49e0caf3596515a326713a969f39ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h897294071c42389ccae83d0af98fbc77195669a5abc3d6c362db141840e86905724acd9ce3f5b008a8b53180a709f70849189460567f583282ed8b4dc1436d582b05a29a87efda307b2b001259f61b8ccfd68bc7e6d6402d2842bb39c58981c544fb9775ecfc5d59a67439477449af5da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb84d9596cbb14aaed50667f2960d9791fb819efa78fcfcee90390eb3457072dc7b04cde4bd21dfaa2e327ca0f06319367500fe7e47d36a1edd2e9bb1707bec13554155c12a1dda3b84d67470c777f27daad5b7d04c19a9a5b5dd9271f5b9c51c74b00c12395c97ac615b2ba7734e834d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cfb7b2fa3dbb79a93d0377b0c9137e73bea50b8f2c430c308e009caf7408177e2c0c0f685c97e08e038b2237dd53bc7aa4d5c853c6e1459070c1826160d039b333cbc76c36efb2c290b5aeac40c1517e85de7ba19037f470653185ceb661e935797e04d93028a22df3d7fbcb223efd2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha59e717d30110128a4a96f6157d2a738f94d59e7cb87dcf429efd6951b2f2031c7da08dbf4a64e80917e6b982be3d08bf5b2a9752a51fa4a1a8605e3d4ed36be87290418b47da0284d37e1f40445d2a3899f17c44f605fe905c4e6d4b8f58556fda4e221dacf027e1d9e615dd808dc42f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0603ff9a5a99992091a7199916b86e5cb940bb44275afbd9b2372dbe145f5a495d496d8efddafda0e781e77c8ef698c9df1a1d922e54c3cb075a81870a20d80cec6a1399486d7583855484f8d7762072a9531842aed5a38a91c0aeabfa257e5f4d9da5bfee1870e23276c660c7ef741e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha80a40b2863d9449e253eab0ad6b0d3d408b929c948ab16781973fc234db2865285aff1b231c8d4bbc0145ab2a64aae9947ae94b7c0890db80f200ab733ff9478ba12d22118e0984c138f07f7236b6938bebf733f8714a3ada42d0a9b1192bc8f58a30e8e7c39b16471db8f4c8a7d8b74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h845be1f5639f9b1449eb115719fdc2f95fe4f4f3e4ad1d60c5501b6798f721d3c84687246136c7a8e77b9503f1f6a5c2f1f781b84fdabb83e912431e3a8cca7d06885af6871848db9f5b8a6fb42ae8f6a17416998fccb1d1cb51370406b38a84bf1451eb7855e83fbe8741047435cf264;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb0507c836d5d84068d2188c2455a66ebd96be3ec2c3a1baa34a70e7c48473201b32354b694cbc176e092824abd7071b375bc201d4b8b9d81469589f90c681af72528c514e8aa4bf73a570fbd28f8f383f33774bc93f261521949c5befb2c755fdfd981d406bd96751013980fa7360cca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd03afdc61fd7d944d7fb696d15afce3dadd56447c55a87063bbdc4c4fcc405c8b3d2d4f41016681b67c32984206508eb3d84e00ed66649aa48caae3a7a47568bc14ef162cfe31147c15deeac6d4f938f395afa9887d12c2ede3a64ea977ac80fac87f3b8b38b41b60e2658a894fce974b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h922ea4e137063d521662433b41b900818acd92dedf43e590ac29ca54cb15c6c0aeedab0b5be8f24ff4be681a0a4ad5cca22b6e33ace76c7bf7cc141ef7f8b96e0ae5840d04298d1907df44eef2e2af7796d6fe5a87f85d9f5d65f473147a5eb399a07a16ad710e45e87dc5ebd853af170;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde71e09db5b9470f4e92f975a35bb5d115fca06c8745c9304e05e08004169eb1031e3e5f0b2b4ed702d16f233e862537922d3d0b9eee5a2cb841081735cf94f0ce94060bc2ccea956bf4839d1941ce3da356f8360ebfc3b147c5d62a1a48da3308d581e6f448e4be8292cb8209a58239f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d209ab0fb4eca48be92f19d9db20e5e62f324cea9ddc8d4914864c66f7393a298a0d9b54d15725a3e8455c5b9148a93f267b3d042cc4aa871d9eef560d270e37d42535e74bc03d0db769d883156c6ddc0c2416e5ea5b2ccbc32b8e715ba70f16c77d112abdef2c3505e36cde5d6861e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h339a08dcf21f01e26552e4ba825b7d8370a48bba11ab436092be2af980fad6e64bb5042e9e43fed36d9ecd9c4a60818a79d14cace6dadc9e3abc8437ed18dabd83dad6aa4a27401b8648ea00280845fea1386e2bf85cfa0ebb90c5b838df1c5f828c35ee3fd9fcdeeb076e7d6a0dca7cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ed7135fd747661d71dbdda2083398363e10244d14acfc8ae5d5755dfd8f1d1b3ab0d64fc00fe1979bb5d7562552dddeb1c25a80ae874d85463f3e84b59cd9ee5dae2f1cf21a4fde40e370d392001c54c1c32624e34a6458b38fb59fb34e6fb1246a51efaa337ac27de2ec822238dcafa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf57d3206c0ba382abc6f8dd4841c8b37b11513863f03c226ff5aeff9e174490916a25a2da2b0fdc10c61bd1826a946040f542cfc875f6318aa80f49dd6497ea5b3e6325e7eb6e1551e350d5a9d3f9db86422bf08e7933ddacada8e52e293a10cf02582ad994b4e0ec7cf14eca356d255;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d14f7860c7cd6c10200cfe7032ae6b271b2a0b5f75cdc2074add5e53c11e98781dfde2b485cea4cb886cf773f17507051c6162f5de6652e9db361b52ff38f579e312422597f501da3ab3f1786a180ece4822f0606987a912f4550e1a78b2f97ef566d67214573ebf6482fff0678f4501;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc74f25abd5a694d3d7d7d93c301620fd0e4e19dfdf5e383ebba0a062edb9645f63291f6a68b3587beb402acf94cd1495db473522990726ecdf97d0ad126da1166d39a8735d58b760b643a1b3b0bebf72ecca96f780200225bba6a127d776684dc355e0516f383a85131c35c5876f66792;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55dbc6c54a524e1e163f1f3d4bb9f3b32ca849ed9c86d27e2d70b6a5aa9a4481c67119933c2a8c93b50f11ebd9f6a2b41cb0127715b815426644b12ff53ef13118366fc528b44444b6e143b666c0f0a2229961030552f3b3aaa20a934821bc50cc727c20335145caff1d562751f9283a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdabfd93b6026b320b1539f38d658b89a48789df1a91746f1959ce0d010eded3d3bb28bcf80088e1ee5ee1943aae29f87b5d0bef6fff40e84ea495071de3542fc8f3a4d2d2640446b0446aa21b5e9070e8781f1b15cb2e94bc05c3fb54823419b4629882debfd95f3c17a7846286e88bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dbe2f123047fa4c02dc28c34f40995b80bcbf9e0f13086e88517c52bf0e0f6f3314052faa5cea2aa6a3eea06ea5ae9c38ff1fa4c980dc1503db3939a464be9027068f6c5f87ccc53a98ddce00c2ce01b2b3746249b734be7e041088f7c13e7e0890395a9e3bf82b51b7aafc71b4a76e9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he599c5c8fdbc20f2f772e6a3411d73c2a73321769a04d728530e53ea24a6cf588123989f5ce744a17245fadba6ea3b90941ee157f1510ce22a3c6653ded25c57d15efad3e4214f9464dca6ab3803769cdcf54373e5e3105f8af69fdc42d055d721b3ecda4e45ffc9e9f8de42ae5a710cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7098efac9356ef76050e779d3798d73b8be0c4a3921f48ae79317391a7153c8cfc70d365852c00f6b98d1eb64b20ce53325150b37da20465e667361d9d8447d3fbc6717661342eda9a93fba7461fce5fe1680a1a9c100ad943ec7d11dbddbe04e8e12dfba794185fe01ece762482df1d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaf142683010feb516f0dd6f94c734e3c10323486b2eb74de024f480319ac530d629e0578afac6d6c5ad4e134a5cf35c036518bb72cdaeb8a5e32efca501adc5a6f8a83283ee7708b5b0f5b36255c721963de105d1315a06ebe7686468b2b2f43221c4defff351c4f208634219e05689a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe123462919e2ed33155ae312867ee2a7775d55f3ddf18689b7a9b6a14acb188a0cd7ad9d5df30da7b5153074d035388f589168530b743eb302dce5c7106c0acfc85abcd6f5f4dc9349f2cf515c2cc919594a28c92f66f33328d7ed171385026a447bf7e932787d9b2a15850ea15afd8b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e73a3fa288a9ffa4b18996189e28b1f0c40d1348d595c3d5f7688bd5996dff416133b0f5f9118373a490c77aa441d6449e1ff71e5a9a34dccc0fdf0539bdd51dd984c51a22353985fae528f10237fcd13895e278a468912aa50113e342ac0e79f68217ca54572e3be488d0c32a8c869;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfab72d502a4bb17e6093c8b8a32531e4a3307b99542157ce2e509700b294e5837ebceddde4f58ec5d7fedc852540ed8bd4b2d492c2ead994794f1a24fb49a84d30fb381f12e126cac2c16071473b039849c501c0caef5fa794bf166560e1d46166a211525c6dc5fe0f0874a9a20e48e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc681bf96b10b2fd0245571b42e4aea93aecfdb71137006b09215dab711906fc5e7f4d27b94f6fdfefbcec028a42a98a83552a7a59108d830966bb9c75a5584a20a7f9972c41dff15de6e15aec304d3a0bad3082505d8e4fd0eb67f675785637e3af732d85e941183632f3ae53194442f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcac984b97f424f1dee0b147de75f973701099d1f0931833a4b2a6ae8f42a5ada38c0086671e9710069d2db7331f016f4c93fee3b89bb3adc2142c363523e3d9dc3886c2d99030b7c1de6d5b764a45f0bf20585f3993cefdee11d7c3a48972d46277b2a01dfacce919e02a52f678511d52;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc93f19ab929d325c5e857fe616290d2d8fb18a00d5d082ccdd3c951e8764857c2cb20fc09c23f8f91dcc6e827d39a4ea6125e4507e071bfc61fcd80a961eb5adbcda1c9db636cf41c861d9a66c47142af46bdadc1cf80f71bda84ae900fcba9b3385ffed909d3db1266d228f2af49f20f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9807cebb8758f058ea6e8b0c08733ee016f0a7ea316c25f16cfe8cdd5dd6bed4752d8a02f1bbdca2dbaff2bc53e441edccf939bdba08704a0c976b1123be54e2c9bdc429ea951b2db298a4031721e42e0264297ca8c0351b41ca7561faec1d860a0e54fe28c7b8e77ee11b9d619b78212;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8aa8058c19be1d8cdc009316fd08e1c96b4eafce04029a45b67711af7c1acdba31faf52236fc89cb4e36532ce0886f7caa77325724029493c7a524dcbb1673ffafc4354d812e1a74862a1b8e5ec5843b073ef964ee8b77c8cb02b79462ce9b36ac43db081083902eb06dd659fb1e3cf95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h308f3cc8e9647f29d927e5f45e327e14bebe5c173a38c449a31ad5534add8faa9dedeb7236fa2b69688e2f5638d4ee72aee97039a21855aaa207a11ba2b7d6bbec2f20e6f8a28164956ee606c7be35c320af0c8d8da58c4756a3d2559cf7e877a527d92175e90cbae9ded098bb518b894;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2df998c2efdf9b567e5c93e37df6b2f7207e3498ab5e212ef060bd8e3585f6c240601e4480e697602928e2330895ad7b89c0bef77d2490a4d0aed7367c06ca5ca160388f240f9b35c1b17b250b4b3ac184781ee4a2b7b385e6faaa688032c6b1731e787153131a7de78d20c5890cdb901;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81e0434813bba8499a9da5a0126cd3eb4108dd0acdc5c39ed67fa6c570b91fba53fe2139fb0dd0030bbbac6ac73ea87c5ea83d331ce32f157d348c4684501f7ccaa2fa9fabeaba0695e21ed0648648964441c7a2ecdb7ae4a40e1dd288e41172ecf1ec79d5faa1bf479de74c1d6bba3bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99084b7d564633c567e4a451ea50bd479758130d8828b55c557cc16931e0e0f454237b11832a0ea4c58bd777bfad5995847b499bc07775fa38c050d5dffa9b8fa38aa7b2771f4cb16a724e3d8a00846c1ed03cea734ca3c5a9ad6cd09ddb5f358a2b15448caaf4238da02c6ad51ffae98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaf39218f2485c440f3ce24aed444ceed6cc7b59d0c48a349bd3b03a4773939177e12f6592f36d765b621d9e95ed71ad5a49dc6615fbe6306e0a5f42bf0526b253f2e14bb2e93c8c132ac2b1dd02dd82215ff2a0fad51c57de1b90f1e0e91aa37b04ba5d03be925b78333da48399786e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa74351461601cbe375da50c625752b6656e12d313fbd446561898f3ce9e82e16974bad7bfcfb041bcbecac79b92a3971d3ddabf00cab244398c536fb81a03cb6fe4e67946845fdea16c253a42ea4f0ca739cd1e3da9e65a9a7c1d26817635a73be51521e4a69209b3faad0a825fd40a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f50704325aeed177db08aa6296b3e88ec79914584e96d803b131d246be85faaa05e6b2894f26a08b70baa4169a8c8b643b9367462cff0f65055d75f1592695ea64ebe69b34c289f642b783fae264f9f1a753f98ac98516be39f6dc1328a6bb99855939b7b2af7ef36fb03a685973ae5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2a1ad934b868936f1f2e4940ddc1f7630799ddc8db84de8ea270f8e75217482de90615a9c450acfdc75c2713d3a310e83eafdd9c8d07508ac6b59d82dbd51430767146916e8b84dd935b1936df8a535dad480400553c17c5595eec8f3fb0cde91bb4e40f3d199c68815f5d178f9f015;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaeb267dfeacc6eba589f320d7deccf279a3dca2c6ed2aec9d80a92c5856691cbbfe52b62a93ac6fd03e4a66c88956fa05e12bc5ff88583fd6cac7fd823b9040874a35e0dfa562fdf62a1cad598ae8b35131073a1b641f664ad12e807bf3edef2506049e705480eadb1992d4c5c4a7f53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hace4fc22ee87d0f9c037db45c51ac404c46e6b8fd1732edad7e08d3d0f82c3f4a076a583d1876cf8d59849080e90ee82864305461f0055479555f963da376550b42fb117b090f1b8ccff10f4c732a72807ba8f155da8c596ea4a6fb29251f04beb3a7288ec6db293cd43d0cc8bea6197b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e1ff8dc9390e72899e1584fba5c900dd10ab3a6a4dccd7d5a9f79a38fb585130262afaec762005e130441a631a2491284d98e162c62cc25cb74d2856f1b254d5429ea1e712bbbcbde3f3ec943b36a330187a6073f4e7d563d7567b192e30ecd86781baf4011fa1e4828b3f096e86fd18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha633388dd74e5d927a9e96420f6c9098bcb954695451d6e7ed5395c0d1a4bc7fe894b78223a5a9a7bfc6b733a5d5d99293496503551d07b1632468f4b3927e5483df4d1a62b2331db5457e9a9762890da06c2d4cc1bfd8e1e6500df3e013e4ffde394451f76f03d5af5df12b335f3a549;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a1bdd2d9469650ddee463724b67a4cb537b25f298f288a0eb5c824afdab7b5d4feaa4d7e12605fe49ba1fd380d87716059f16b7c565cde850b07db8cdc323c7d5cc06eb012ef5d822b1dc606628bc4e894af73c64c0cc4d6a4207cd2be3eaa5fa4b65affafbb1b820525d9cafcb02515;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9393efc19e5512eb1df542906f27ae3088ee3fed51f0df8d37a59ecc4316ce6c7fbf1a72cb954a403fb5079922d8abde28294bb588ccb6712395f2962648928b0dcf34f02dec91cdc9c5d96d3f216b394d5c7f467375773adef39d0f3bbbec32e429fd74b56fe2d80a3b71d37c46e3010;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdca75e0e66a5362c072399829a58a48023db10676b2b82862350efdc832554cb95c90ce2e7fc94615273b4bd5a1d7bcbebdd37a8f03a82e3529ba55010268af742a48a44128e644581c1d853faa4d3fb17f903739f5227deca7d4c5fba93110ba7302b483cc9ea81abb87432d6f8bcd80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8626be2a9d4e97409a1221613128b1da0f82526bd7f2a357760154f68966f569ccf8f6605527725b4ab843c066a22389b89d3a8bbc3c2601c4e47e75883d9c77f2d46345fc4c51e0eb81c759b6f6611e672567d6603b4d25a7e21631e0886da138ec43474603545bb3526dbf3f9cee314;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb61cb45fb912a326dfad5b0cb1df3a6d0129cbaa94466fe2d2fb2c4fcaf0e5300c78bc8d75c26949f5d98d35c9d7738a4c27c653644c7933c2f2caeffb03f3fc009d81a0f7964f882381d8f9b34ac70a3d01ad9ba16b1a57ecf5065721339abb321f912c02f4fbc2f8880b053f78ffc8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h599f91db628652c35db6e25d2b85add95bb290b16860b5ffc3b684b93c536a2b045bdac9e00edcfd438d1247b788631869aff3c8d633aded2ba430fbc308195366be33c608a4b537f1903d30e1f96dc3254d2315587c7b2d61b540c9fb49f5c817397e356e507075e62b2b777fee36a3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd198c0e89294dd906319d93e75f9732ed2260333017d5b1259a4314ed4e2da3626900dced95361ad0bbbefc73d26c25e5914f28cc79a31ef5b2515aa3445f8c4cc34ec806b61855f85e4c63869ce82a5a964674fe05e498aa3ef343467c9bbd625932a1e9735218e7906eb2c7f476d381;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3d053a1ad348ddbd367d75ec5be2a45150900b4d64724a8b8234f3307f1c5206f7ff597bd1685cae96fb3dd3c98c3adb934e78bb8a1b36522050ba0f3dcb4c0aba42bc5c2c3abf38608f455c941b9987bb007cc99dbb0e1e8b7562d8ee42baf8f3c113f7477965e2e68d7cd20d2a6d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99176639b6da49ddd2b591ed7715d252922d933e3755ce17efa26fa525e9ad89fd7afb8d7995848d3d4a7092a02616c22e3f598abb864bffbcd3408ac12b72cec09ce9d43a79dedbe0e451623b65e733e42ee62644bdfd57ca1fd252af3e28c0d0877e07c032413ea11abe41715e9e221;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb5b10a78cc7fe1798019dbe092ea0945416fa22ad5089854c4d7a7cd40db5ecb9314f4ef298e33b725406d6009aaac2c93de5c2a694f354794f849a21d9f1512f39e003209945d0c3e14e4a1e2951d38c4f196ae19d7e0bfb811bc80c192df363e8f58136afdf6dd29156af1bf1add2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf4cc63f5fa0656dfb2a4386051aa2e5fdc8f258d8cb30e986fa2bf8fc198dda153f6d668ac5c2a43650074eb01495fdd80ec71a5252ba5ca11033c41f0d4820232721a19b28b3b948dcefcec631c2c4fcb78c1448681e1958936df34703d05bb1a255b42b920d84db52e1a91be29a687;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he76213f1a29c8e206337170bc4af64bc7397aa974af7eedbe72a62528924253f073c67417ae4b6782f4dad69517f6214fbdb8b7012372c845e13dcf12e31eeb5ed25ff922d44d13e87bc20dd8a2896f7483a64bb06dd658199669d07dbfa7a23836745a092704b7d354928903190c4b70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f05c07cd8862f227b8e51e0ba7628385c69bc7ab0386df61ff47ef8e6dbf0dc17378d4425f68afde4dd220446035b88ab7561ca66a14d167ad3fe1a35a6ab0ba44ceda8aaa1772cad34809460aea99e6b40ec8ba2abec3914e6cebb6da144f1095ba9c76ad64e3d80fe2618f00c19188;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf35a365b5ee9eb108847d1fac5ab8cb52f4408bd1898d9833dfe4083d29de7aedc32a927f0efb8d3b23807b22e8533d94b85273b9ff3470cba8d484737ff9f600f2dff9274aa0796d1a31ffde4f3d3d6a6e4dd5fd9b91c1510631b98aa8e0c6c6f2c1972afe201dd3ef63f3bf7a7f30be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6967bf499de0855574bc73dee50007d927589070d7414e607773730d35322375898365e82d49f98169f06bed8f8c26565f6bc9050c0dbd8f0a266171fb85f125ff903d0058e197134461af77f927cfe75a06500de167262bcf4af4a4a9ff8ab8dba81e05cda856f896e6ef23841c794;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf9e393ca95c16007c97eeb77c6c26fe0f08609ce4abe6c9cff9493d95a7b8e7670fcf7fa3f007136158175ee702a735b0b89e5083a06b42580cceb3f65579a7a7592b57160e19319444b04442bb9b9213e588b3b288aea661b61e80613a44aacc04df59932c091b7a79c3a6e64a7538d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc763f1fe03c507d2626a65df70ae4445c65939d5a975b272bb08814ed13629c664e1322c52b88acb99fbe49fa12840044be7132adbb8f7eed7a53e8b19b8b2d7fd091dbfcee796329347e2ab5fb09c689b327fd1f327a95c3b2016071bf0745a437cf2898c6aaa5bd528956c617d57c41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2bc777d8c494078f49ebc1d37ba60eff7e2417c68fbff52b07377c91652a456fa5ec6004151008b0a042f3989badcf1b3687d3a26322a77c02aeb81e9746eea3dfb2390bf6a272be48635f8e4dc13d7ac8312d3cd65146001992504a5902535a140ee274477b4138b56ffae0ffe38135;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c137ae5acdd41dbebeb52a929c4586bd47be4e723a31128c0835e74ef09ba1ec0e947f9aa821b2f2f333c7362e955bb2866c4ad32831d22f1c24718e1a277b5cc385ae7aedfeb19c28c8ae34ea39484dadfaa5b6df26f1a8328f9fa7c8c66e7b77765fdc63ff5edaaeee90a766221d2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8893343b972588deb2f43d68e08bac95f960b2318594981fb8ab2b8de14c5b527b04e603db5af720ead6c635a12c5dd25387a59b3e4975e4519dd3ef853fa88c272cefa714ce4226f5fda788f86976c29969be3d753bd5054fc20495d50eab615abd90702d33a3736cd8e4b623b52e77a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha832efca7295138971746a47342263ccb050aa19fc53b8e454f080ea147ef18cb3afc1984250c3f488180d4e039b207cce9ba4ab7976782b206bcbc289097292708fcce3595c87f0248b0e6a7b3ad71266e3216bcb34dd5480878f736919109672bb94d0eac12df65aff8cb80c7ca4ef2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf08fa743e8b82b92000f94a8eac63565b0913aacbffca4707c77367ca084113311a037205745442485424efd0b94bbfcbfcb34e627f61e5ff5e0ff0a6fa12bb83edeab46811651294973fa259e0d249aa5c9af7d4c3a332f14f67db46c310e49ff8dcdc3cb9f1773aff1039ac494ef6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h200c0ec655aeb1edcef6ddb020ee55ace4c2a0d18a5c42537d1c2edb21bec445272e4fa72132611bff5a2938dbb7068a4c52bd9f927da7b527fc65cb31283387c16702ac1bb148732fc18f9bdcad0e6b2b7a0b6dec3ac920b6893cf647f906e5adca75f54fe9eb386abda83286f6db68f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7c8ce2c29fbeaf06771eb0f61d7f6ad2d1143756a585c72ca4b6aed3b92c95ac5e9869c00a139e5cfb62ebab0712a8d833f48ace00478ab3ee79f2530ca3f70d1519990dc1db260bdb0ee484ddae00ebb0bbbfd2c5880a4f5655535d88f6d943f4002d8ef4617bb8fee6aa8190573639;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88580e3bcb39c7f8074a00bfcf6148e32bd65eb525d2b2a2d96f9e03d0562bc621b331df4150f5aebc8d66a851bfce10d4f0a51587e211f72b05793548bb9c082b05d4a3a81a26059c640e20085c2c8b173e113c6cb0bb23c7ea7d59e688664b4e6196e5fd49d04858d480c034affc2b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h977a5ea987580296c1d0522f7fdcb438810b90691c2265aeda63fb7b7241b78fd84676e038a49478ce2f00dc31de211752dd0c2c723e2b8b8922fe306b6339541edf972b23872b78064937cfd19550007363cb0dd27a94d4fb4228fe36008f7ec738999c6e7ebb84c57e335e784e45060;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa01286cde4e2585858fcdf5e965c0dc19d5d190ac148ab856d68b69fe1458642e99158d364cb08cc2569744896960bc475ccd4c04fd4044b4caaaa478abf6390f74e06c15584e49ccfc6f8308ad6a52ad74147a8af165a05fe287a652e07f19542f4541c57d44896237c0253fcbb9774;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdea43ded74135715c04ff3ffff5a8a85ae2e6dc493ddfd2e95988bdbffbf5a346ec50a033b12bd8b44145748c1e010e81ce05fa8c0e18331c4cdb8ca9f282902e95187ee125aab0353a512608dc855e9d8c107c307fab485b377c335e71dae8912c95a1d8d522192c3b1a3cdc010116f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf206a152523642cf8b88e2cbf7f4728d4ca61b994cba362dca1a1b50aadc6dfa90f0f60000f340224a3c585d65281faf8966dcd24ccefd12819fec0c03cd7ef64e3b50ca73488ec2828b28aecc13b797c64285305ed613634e2492f1a14b28607b73c47271d618b381346a4fdd20a7f12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d451e066d4e2b50366a0a38e4c759243a767a4739e24d4c78fc11a746448fb65d5520ed1a627e263f2805f5e883a9bd864783b6c71d8518977ac3a3cfdc4474278c43fbc512112892fd2ae15cc848c43154789db85197c42c73bc850111c4806a2aa7dc24e22bb35c67a597baf533cf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4dbc624dc36583101197d6de1ed708fc44da9dfa67b86a2275fdf30ff49c4a4a17f6647464a8b8e05e29102824847e2a96b122e590ef65d263c14433940ae23ee8f9b210fe930b9cf51cad6c0e5ddd8d410f7788006fe4af919c91af3888c0ad9730deb1129f4e6226cf60d8a1fbf617;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f1adb8b862f2f3eb3233dfb46f3ff474f2390f95d649d10266d6c80a07818715677151a393a90ea497adaed49624f90d03ac0338c19e40b1b629e662aea50a84c3921f1324331ba1ed20915e00df6fd46d7294953c1e3c37862d0df92f9055c0a8865774f0bf934820ef1b1e381ba06a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4031d5f9c3cc6e7bd94080fbbc4aaf7e84e21d71e0b93481c1c513a903144c97d59c8ac55914aaef79ae876bf2d3e92dc584604412561c5f4c1bb668281c1e064f11fb862d19bef1feefb8cbe83a7d176eac8fed00a074e3ab4db85976f43e5902cb25f46569e524270ed82dae4750e6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cf59b80bae38058c00e16f892b14c9a1ffea929db80ec7145bfb55d5d10a0c016293e6b8696cf345dd5f30f1e04787ce12693794ab7fc8260e222103a930039732a47899646a58b2765a85c61d5cfeb628d02b5eeac154babdab581dd5243498b828d34235e42c34f3a34654c6df7e9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h401e51c88e3f0b7af442624ab134e4b351307ee8c542c4c025ec99cc012934826b31982dceee5f9227f2692636ba4577ac8abef43fa28d905a0e005098afb418b6b182c27f00a4b4541f343b6643497ed15bf756b5d1f59bab4649b0c51318680ec9e01a858300ce8db8cc0b1533806c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habe7bf401fc534282898df4e1ed5b6f80f35cd7edfeaedc94a1b3dc873c5ccd4d8849c89ac0f9d42a6d58978d97e1d19607b85cc2c451633053a6c45f60f4da55474035baa68df24a7a08d3856695306e0a22dab7e4a0baaf83d8d50f564e1e08d83f32ef572a2ba1c7d6523ef86bbea2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d608af6d2f2cb2751d198987b99afc979aaa458f9d7411d476bce3f3e4b437bf072b2738ab6fe964659937d981e899bbb70b08b103fd0bb7ee1e23588da44e692426db64c4240aa0a4611e22308f2f0c851e1043174b9513d6a246d9b120bbd8ccacc7d677afc4772dd9f8ff8b9d4a34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab3753f9a4deab6aee94c5fcd45b27d64a9e0007caa388cfa3b54eb1b436209a63d5ad4ec0c665771c20577389e7faf9b8afe084a6c818d9254ae89e2bda5182969a2aa5add75848634cc56fe6aa22625abef42c3ab20fb6653067be30ae9f2ce70f0d31bb34bcda90586595d36867700;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e1bc6250e1e6d461a81cce67d3392c07e085689c45bde613e58755179f94cd1d550fa508f3876562699b439163a2f2f1dea1621653d1b8d387ac9dbf755c60a53e85ce031fc92a0d27c420bb62ad8700a8680dbe4be4a78efbad6cc01a8f3b9ffdb0d02490107167bf733b6a189af1a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96c857b02ad2fd09b4def2acbd2e188b1b86a1f249e52712570e4290f24590dc4c8da01935244f415343d4cf70a0b50484dc0a062aadab9fad6dd55014de367549a131e09ba110d539f2dfad8ce71e0a293973591f365d4dd5a4bc639ee0c7f5611dcd2eee8d8c5cd4211ede5bca22009;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbf1ee2ca1e87629c662d143f514835f44c7e9ca27bba9e9e93db7dafd510fa4ea409c7ed87059bd1568e38af54b1b83a5b9204f68be06ff5ec0643fad1587c7c617e2f62f75fe096abd810f2d6296a27b2c19170eefb482db7029e6e34ea7cd41e562f8abf855122074e282175e8e6f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf4f2ec2c4f61809e58a95be926f11d9bf5e8d5f056cdc839d94b95ad158071bbf6e964db7f992ad13b8c8730472f46236ef89beb00f74730816a7ef9c8df48be2cb39e472199405141e911a8cd6a398ad3909b44f412fac2f0c1ab87ab75280ec46f0aa0b90c973cb9089f1889bbeb5b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7b025deb25c08beb9b55911eb656d7226ac43ad1d4e48c223fa42b167ac3341e029e952d6aa7e50dd543f421272624103aaaa08c69f446398771587e49badb61050ab84edd4337a3d5c811972beeac4356e8ea20dd74ef6a603de127b163bff86fe16150e47650f8d39909484c066cd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6812ddcc13382eec0a5d42240f0952bd5c11c0e6450e004bed7eb09b887689d9f12c28374bc3cfd29a439be8ed939c86c29ba88edac889b2020d59c5a63f1ed46dc19513327d537093d477a1ee30a6bd687651918bd4aa56d8d90f39616232da4ab89e3b86d19797951ff890d09d55d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29218d3dbbd5b35e04d25272c2c1c42ef4ddf1a433517ed56718920dd9b9f263af2028d971e6572a559f1f1320f83d3770473a2dbdf2eacc4f29fb8dff602fde2f223642274cab10a3ea472b2ef1546a638139c28a4e29a27ad838fe24966140d8e032850cfef1183472a1d5d43e47c59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8402da90c6cf3bd23f6eb1710a900cdbf7a9895e259f123851003f1ad6efac664b37acb24a36ca74b7412b40e30a1740fa4bbe1e5b8fafdb67ecf89af454353829ee6ccc41e9924690ae161e8a29f1b2b6d299707a45349d81b54b936a1761e7d09f47a141a4f01fd5ecfe1db7078146;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33df87c03e159105fb9b10c776d26c12643a9cace89e3b7cc75bcda1f5467b269cb0adb9f2b20f4f1c792d0a15ee441519dc5f3702d6fbeb3acd61f64b4c9dab511bc98baa0d5852e9481b36668c73581e18f71864282d85dace22b1cfa29b591ddb646ebf8f38aa92d7c94bd48921c62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb149518f7bef85c503e992acb6553a99221610c6ae7859d37981a086ca1c067c2e2b7e587d1693102fdbc890b5a836e00da8900257eaee04205a15358c6210e2161744bf7dc53d954522cb960d80a36e90241b24bd81a88186ba0b0adffa0eb3a95cb079ef517c2bc6fca12fa070d2fc1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc567d0c5f275f0985363af6a8059388634e586e0607a4e4165fb9ad0beeb23c34b669981cddb821ee9b8873ccbb4a5c7b5be47952b5b7aed7bb7c028437d9e38633cabc82b5251fe2915838bc5071134adde82571c01050772c0290d07f255e75b9287d84394cfce6869bdf3445ae1db5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40ef0766d71372c7ccd29877349340fa1a689ffd6dd845d425e9bab23bd62012e7775474f3e78410c9d123e1c6dca50d6385bdb9e9329e70509588eabc20b2a94f1dab01434c29d2ebc89646ce3163dbc872ca01e23131db9a08b25194937681c04709a8a3c46dc5e986d43df25115013;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbbedf6bbe1830dbf5cbb99bfd0bd48ee941b65a4ce621b4c76ddff5cd8f4ba7d0725cbfd7e3c211a9faf1964e8ea84b82d47f27c52bf12f7c0d8c6ae90cc29f047f0dcc3cf4e525298c1a3265383b89fa1be7e06f674dc880083828a3143764994edab6013e3425c8c5d64076db0cc65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3eb6fe9fb53ec824869b8612706a90ee79648f6fa85be43b250cac76dcf78f70f2070f3fdc7755aa5177e2f0270044f666b3fa6cb6828cf5c07a997af2d4895031ecb234c8323d58655aed72fb0308dc9eba64163ff64b19a013d6e7cb96926680f4521d0d0d9e9808737f84e84919b6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h908cbf93de0d788398c6b400bd0204dd8df91062284dd607705551b3fa505fe1af690f69898dd99e623ccbd2c3f1daf8ef8dcf1952e6231e6940e38373d5b45ec5b76ad08e758fcfb92e34d85d549ad35d7463f74f713cd94e3c635357e163eb9783d419cf0589a786548f0d8745e458f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e02707109d0703d0fc71ee00b7b484d61f14f5bae0fe300ac40dc6175b5bfd6c8dda5cd1af064ed4376286ae70ff71aa3f1cb0026ef2a42e7ba8af1d51ed67e0a2a49bb26b4157953bc538f36ccefbfd047850a178c6d2a759637fe4b5e8cc9919cbfd5db25079918e7efd8c5db21189;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76a2a62e08641ebdb34d6dbee84bfc97f3f840958d1645d988f2ec6a207067a8f420d5d2f279e0de52e9b1585f31c09b7d0def8c8e4229f5577720664a8e39e4e8f1bf5d1f2ffa806ecb3789dd6795274d6ac6b0f7b4c52270414a38e394ebb36da65119aaefc255a776aa823f1b1f43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb83b29310771af4adcf687ca6c7549eb5424f8cbd545ac8174d8dd3b4afed4803d9edd14fdde208224b3f528cfd1ca15796ab98ea46ac5d90e326c68542c6e8012702e1d2e8f50c66f9f489d240b219f44467fc6e686f3bbcc6fe1414272cd3a8ab93df891d28b149ed2a2d5abec2a19a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb71afdab0ea84351a3e0e914129deb7dd2641133cb9daf21753688d56af75c3ecf1ee709462056483763e1fb0ba987e1b3eb3190a9fa53eea3332d417e0cc0765383979c5496b97d1377c7243587c7a40404539317696813aafd4b0ac81a6e766305bba93ca30c41dd955c203dfb1318;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefca6c314b120894fbac473e7a452c9420d2492e7fc252138b82bdbc37737af1360334345d5bab6aff6dde48bb93194d254114f86c26231b5f255ee825af220cc02236f37af56435f9240d96e002f08fad84f4bd49c988c76588f1a3b250f91920cd2825d980f877bed737bae487a7a81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1784322e3aa4989f1de56e2fec008402079ebca4e1d657a7d564a94bf27eef880ca7b59c30a8626d24b286861449b79a189ca433a1c0284286a018e0d8c4b8f05fa77f6ed922e49b5a77d295ec9580d71404ba2c7af2f047a63a0446bb087a7e3055b3c448ed28e597d6c984a597afadc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84df71026e16c237008c8b88eabdb7ef58aab1d216f5cf3fad942bd40404f6c0ae1aabc34f12ee22b8a2211f22717d0948d907be6e595f4b5b3f280aca918cb5acf18859cd41ea54ca53277de9b0f2223ace2a7a52913b09dba2f8931fbe1132dd6d9c4946495186484e6ca82fd83a308;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bb4c08d9fd15317c3caa2db7b6c1f1c995c6da784d43f7d88fdb9e15a6b9fb3e94b1a118c4272b07f7718b9b1fa184d43658fbccd3602d599ab9e6779230e83e0f7e3425722317eeea28e67404fed927de3b4b2a1f4cf858dca472bab83010a28e048da72d2406ba8bd1ff3bb5d6e30f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a270a38affbf299472ffdaa7bd5db07e372dd8f04f6498a844b0c1c015d3c7c4aa9952fecbb71302351d1a81efed7db9491a8be8a2ec1672b641137107f989656e87a3e19ca75cbefc3c8529388b5448d990caa90749bdc31f609d28f0793e0c2bc2d890f0723d64d4c21672938a099c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc75b1e5215b82d01d27780b3232f7142aaddbf64b4444caf9e8de1db19b3e334b5f3598276de1eb96a6154f8844d35421806cd2566da6e77e4304a8a5dcadad17ebe6bc6b579488c087fe4dec5699dce75fd6b7f936e57d263479c11d97fb3e28b027a1b653f418cb45be1767e1d386b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfda1b0e731bf8579942edc5de2753cc78b2df314fce44c67746568922bf579e1c6a14b945c1a3366098df96ce3f8f4e982a9cd912ae19b7f772a142a95bc3cf463ff95a79fab917804b6daf5d95196435a0381079bf306f8b95b0327f256ddc9c72ff0d1bf78239d034a5ac214835bfef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97577445cc35ac571a7ad37978150d81ca0aabe59dbea5117b0c3925f6c99af391848d6fc01f5020cd5d290e270faea1fd9ff7a6f24c997341f8cec8a6568e6138bf4ad8e9ce904a8de5666fc399ff29441d1f92f549eb768225a49d45bc037d9ee966815930782033c6dc5bdee17a40e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b2e3eec27d42aaf1dde54665cf559e26b33bb08c37eddebb8b75767d4cacbda51c270c43f01e877956dbadc6a67146967348f3551da3f64d5c0cf4d70da80334601fd28de4887563ee98f72689be615f50cc7d9e90436409e0cbb27b54c973e9e1b1c975ef9ee004a7512657bc20a0cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94519730fca889cac6472dc8b3f6154785158a0d542e7f87a46eab7a3b3c6c7537c1730517bb48e98f065f672dc5ac1b77df77546fb449e8b8225d78a4fa6801023c5720e63e398a08ee49e1db50369f4da640161de17744082b32df369ed2ef38d2cff88f754ca809f7aecc3bc5f63d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc868736e1696dbe292cf0ded150d7a0f819c5f22974dbb1919b5f1b44ae301286d986b022b1aade964373cc10b6cfc5178cf68697dc06c4508693a25a9bffa1f007a8a4003643fb5879f9ba030462f0c8ac2b72f0a9200f57615a54f9df6d6501e07aa88c9d3a5741e54949125b82d13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9dc807c27d8f74e186e857bf82e1fe9434e07049fd58aaf27738cb562e111b6038426613df3e4e7eb34e8828371023b3721df04d51f5748105c95341f89351583d1df6f773d7d22bb4ce215bb62eb6e4255c7c927e1a7aad5ed8d9ff926bd5ab6be21137b495a46e919cd2c2890f035d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9e841b992e0c7680cce43bcc1d3602c16e07e277a8ff373af86ddeb38f1d07f8ba0c9d20a837b72b998f069c7c3aa123b33e2542e2bc38f0d1f058364e950b882421baa0b1d66c1bd24c00e9b43b6d5e3cc8e8252a8a2f8c1e9e96c08990a18b941f30b38960f1dff8969e8de08a2645;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a32667aa766108e3e79f3be1d92ef9558f0da09fa6d4f8116ef83a70260887b53969bafb6d2d27f4ef7fc6a5c0e887527ad09cfd94e6d015bac60b0f02fbddf6fe29569051743d8ddbefb8954bf64213f93e5af274f1ad2ec3fa4bfa8e36abbeef5c91fbac82232aaa1f23ac29514403;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1326a8b14e16d2dee9fbafda3d9a2186ad54040e40ac5c5495b1db07fd3b8c66b34d232b5f3ad351b3b8507dbd29e4bfd8743d8c103945974df245a585cf4f12ba5a276e0a006f0de3d7df9f6ba13dccd828f5500f453650209ec7167f4410c5bb3bb86c7ae2215d7b93a047e68501a6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43e595cf6e30cfbcde8455b7303bf574c53d6af0469c74bd1fb513e4103498c6b097627fc2f8080f21b9452651fe70729b9dfcd49dd0fb202afd05464bb2917bcd9d16e0397706b26a426457273c6d20be84e9dc11224849f76787776012965c7edddc65fbcfcff631c5f716936ff3ed0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h425a14b96665e3fadc85c1c36dfe2816c742967e81a995072e302644dce88c0b2bfa50d060c6cc7d9f0b906c192e6cd81988b79ade1f0b4b2fdb7cc68c2012a8c2bda9d4a6bea757fb6f838e1f5ffc72ce2ab3377d41f167cc601c2764c3d686081f96fded23ec836b18b0af7041fb120;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67f83b6680e818b68c1108a48c96ca8b0af88bb43676219fa8e9d5d18f1191068efd41b4adc5a0acbe04ac2e232afd262fa1429b264f9b3fcd66ee6b11162644f8427e7c33c1abb7e5164683e53cb4a9061b6829f0d05ae5cbf3870031271d1cea0dc89620d0857bb19967b383aa54201;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdbab51cb75f3684cb6fb19ceee514a5b1540b6b84aed848e77744cce9f18f1cfadfc1a88e7e14dbfe6540ee3110fc58e6db5f66f860a9e36a25ca124aa7d84ebd2ee58b4538c1f74a3cc0c885b86fadb1b71d9a1d366c96f68ca1b965ad5195e564174924d919ea4daa24cc97d3ea1ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48445dcd4bb1b1cc4af76938845f95d31443d99555a5c7dd488744bd86fb3274a95452dc48245275badd0507fea4a15caf940309bd161c717704cbb66c86d4f3f1821749b8052f059798ce63c0c8890bf674170f45755f0fec7c141c073adb38780b858c020a389b0a4dc87c18fc15f0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha89da46fe667474c978bf30ca8abffb162af97b798df72a5713ed21386b69cb157ed5869304784567e430b361a1a4a8f6fa2f60c0e9e263ea158e7609ddf8593d27c5bb625c18b916bf62e3b82d8051f547e484d18e9ace02712a9b32c93198c77b72eab3c8b5ba8b625e82c09ba2b84e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41d8556e250025938ea76e0d486e8a7ee9db2d73783a800c7a7d6a1b9737077c5731bccbbb1f7739d0b8f0294559a85b0139b20eb5afb1dda67da23a26543cbe2043def59fe8d4e2b6775f9a6b29607536e3cd7a5dbe0034011bd4ef36906ce644e92c575a8525fdfd92304762c217ac9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2f03bf03b3158c380fa655b0b0becdd6f6abd7c3ffa5ae2d6f12db980e0ad2dd6f84427ea4e40b4ec821d64300f74876b17601cbcb79012cd2eb6d700d281240fe2ab52516b9cfb006b20e7848c54c0da6f98d7063599c45428b3d48afda1c31e8bd26054adab7d7a7a4b4430dab1a9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57b83c1cffb331c96d0a7d51b2882da39912505e9d8e3f64fa805f13a1cd49ec728c6aa301b1b1eaf35a54e08ae5392b8dee2881daba7492c46485508a054d23d971f8c96a7bf4608f4b6cd8731cf00b5e6c4ab392faa85134117584b70a22c0bc54232708024143b00f7fe3630015cd2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h494703525facb1e5ccda84eca60d8d5a209f1c18af52ab3d64a36f898f6fec3d7474d6d033691d6551c37d98c64e950d7e0ca1e79a9e4c7bcc8d21395cfe71264ee7580d64dabc584300832d14cdcd46629fe2ce71f0a4e312b01f1946720e8e63c59dc0f6a51d045cb2f88c4fbacbe9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac3c85ec1bdb0b3a1c16bccdc2035bcd0b59a12e68650cb453a707e2542bfdb8a4f440f8f95b2b28328011adc89e7d19d190383ede51684294421d56a4cac68537a1a4a002e8f73dfc5401f4c34788e6c89ed7c12ab849dd8a93b40363054f10c19b2cc2033e1b8d98a1f55fab1eaf947;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8fbfd30729a0c8cb36ece7188c93a7dad34d53b13d534eee5ac014ccc64c88bc826bb506d67a9134c0f655a02926c155ba1232155dde62f50a8283804333284a19f06630b9b4d6355143fa0ab00a1876fc38bac91b12249b256b82464b8872ab22905d3481d21741afb074b75798a375;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd53584577d74ec9fd97dc9e8303e56f8c35c6375986b9fdbb8e128fdf2ead894058590af209a464924a1cd736331d3b0643062107b77b6054ef22dea2255dff7f18ca742bffb73fc59749f63ed1ba2d5626a66aa6f1f88968d12a2721e11ed24039c066768ba54375fe455f96b4a4249e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h732e2727cdb378b0d41dcece676f9730fbf0411619e7afa681912369811aa65e28648e75188ced179dc01b61c64d85723b5482722808f6f26e2840109bf30e38b626e968076bcfc96e1b1490baef58cb36843e8d217f3b1132a4681c2acd80d471a88edf5ec413e89ae9ce6c1cdc9483c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e759652733ea0422f7af32b742804bc607c03a0507edbf2c42a4f11025317884b6d9e0bd269fc2ad96b5800cff71ff9df7b4f77beaf6732918f2acf7e192438e4b50258ca16947012257afd911a0135d1b4fe2a678050972f5616d7e4af11de56687176faf2853d2f4fd368f10a0d3c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc1bb09fca4dd5a99a45b74b65090acab83e53bfad01d9680f89e8b74985c152edc92858daaa2f7143d23710a340bc2875bb2697d027a4c3f6d2de8d219693baeeb1b50717ce0bff45655fba374f2c858396e9428c3bb7185069856e0f8ac945d5df385e647c19ce2db1bdcd54ba95343;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4aecab3789d26b0e50451c36c9ae01d65b55d7434c83152e0e2ee4e95be7621773c85bb1791f420ea89cedaf6f4b2a02b8158051bc4f792c91f23646586b0671879629abff31838a0f396ca6ce9f44981926598bd1f5f1f1f34030394788c2afc9999aefc710d85a6d06b4ee01978bd40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h489d01e46251af5f78e51d1dce3ace03ffbeabee4365f774dd6eb1ddef001ff584cca6a97b0453e215716d4b113ace8b252f0715d7e253439594bc85e1ec65bbc2a573be12b9e2ab011be0623596d1bac37565c3d6a4ef7dc37bd4596545b5564ad10cc4b3de6f1743884976501f10329;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4255ae7560a556be3516dfe6787889b9ccfe59920d5549ab63fe09a73df4c78345251676427b03e7db8c6d604a53a697d6eec82218064bd56cd44171bf0f62635d7168c877ba5f55cf30f93b39503d3b17c09205c1185238cc48d8cc7ce0b8438f6636556bc29637b282937149a22441;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea8d43f4809b4598d5e3c6101ee1545269838f0da55377ccd060a1edfd9d435a286ba200b5fc48f918e1e03b19b538900507c895a239188b75a149ec96572e401a2327ef3738a20ac0e6373536b41ed5e09a0880826364c269e9f20bbd94916fda4a179e3cb9496a5d60bbbb7b6ef0a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf34cb245478f964f49b654b908ea9e38f365c0ed9cb023439bfe63d7ecb0d3e864a12b8a1d83eb9ef5c3dd39b2353fa199fe70ff63408d1bebbfd9a7709ac5ddee91d623455ac942bb2b40af36b320f10f398de01a17d179f313f298c390246e990265958ef556657d2ce4a1d575b4796;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b4e0ca024bfc0a1f2f843490e520b99bfa144cbfd6bf1a789269b1d28c83d355f813ca3b4eb81aead8d0a4f765e2ef40cd89ecdd8390d8cca099ef09922e451f7d77c16cf3a7eb14e649b079c946604c1a19db39a9d5eb4b9a8113077e449c9cd628d0b17ce46f71b50f3c82d8d69f26;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3306e3fc821518b735f16c2771e55e27e6a8f84f1822c89c7e2ee077d96ae89d01c5a6638326c74275abaaba060cf5cfc80dabf94658f8b788ea6886ad32c5741e3eb18dd16f8d0c241755ba7aa1d2dc290dcdf0af7700d0a5af26c6a80e15b4f8b96bfb2a5e3f7a5bc072b0e89883ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a9bb638e8c70f0c5f3c9cebd6bb8a993e0070d7c326cd7bde96c1ce3423e720fb7da8f97afd182582a8f8cd66bf787eeca010a1b0563b254dd1febf21e80ee9ad3ec8265f16cba51618ad96d6f45756fec93e12afa8e6741b7fc3b114f496de3693e8db20d42ab5217fe569b454ee37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe433d155b94a2d0c1b2d0f5917f1dd53a61cda4498b727ec3122b0188d0e110e1a35fc7dbab2c1643992cc7e86e736f8fce81e8638f71296b283417ab2420c6b8a363190614ec00b251c5015805ea7825397bfdaf039dea37c80d57025d8d391536436882a434dbf5a4507cfe7144ca9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62a68d3541d8823a3bc854357868d5a58e20c3603f5d996b5170ceae389732a2afc5bdf028883ec6a04b82f774234af8a9f2eadb8f71683d81f88d6b5ae88643bae030f9b13158ea60ec4625e85dd53c35e752926ff1a72e4a555e5ded7d6385e4d7fdcf59ad19befec7e63d99f5f86bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb073b515bceedaa0a28a8c8d4fb3aaadb89a244ca62e99e5a4fbe1f78c5a9342c7e8a157769b2ad8c0ba37c3c4b3fc4744d23f8a6e48fdae04020485d238e7030dd17a758e3e1831e19fa16660032fe6a521fddab752ec4f9bf5932794d36462cbea3d8ee774d4c59f8488f90d1f399f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2456886b105dc8e808ecfeb6978de00972d7668c95d0ccdbd2b7b59c7579fb61cfeb3defeb5b508633618e357a49c8f60902e390e841a804ed84df2e97cc88e1bf9c2003b2016c739cf534606fdf6d10a05f240c232a4ca3e393b8bd2d41541a9fd04988a90baee8a9186793a82e2fe03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ec3c8927bae8b0e917fc6d71cf3295cbeb6e2556a667e47794176079645d0eb11371c12d8d58a0c9bcb4f43c710898b003fe9648e0b9d66f9e867d80ed503f113cf7e23ccb07df779c182538157fe84591303d44436259af4c58bb002c1c859de3fe51a5c9c7a12536a136d744e9e043;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45bacceaddb8f5e944efb58ad479dab3b0cb7a2944ee22b40d8c80989ec3e7af2bb2bfc065912c5ddffd96efa6ad5325be955cd889c64b865600293e88600ad2a9367c0c15bcfe657249b18fb42679e84a17d0800598ffbec889e28edf8172a4fb51cb34764e7b6dd177d5ed72bf51286;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h827a053f4151a42c6a2ea5a4a21c5b903c16926229185c9e4b586c9ce529dd85ae8706340d92c837d6b074cd8a43f3e824a5c73312f95a68b027293d3b06deacb3f8a93e57284cb71b1550d4bf71bd33e084ce6a96ad326b4874c0b488cc91778ef59056998b5b3b5fe4dcf42fa7bf995;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7d22fb524bd5c0400fc0bc92006c2cbaf4332e325fde2e993923b07fa2bebaf327abc58bdea51ca62c5fafa979a3a47f3b53e4fbd2b64434a81e77daf26a77ad471a7aa31cf261fd414b70a06825fd87f6ee374118239dfddc539a26662105ae770dfe8aa8bfc80f3e607a2d1f5b875a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61c59ac212b9d40476db89996bbf0a7a93c893d7d12658daaed7ff5441c5fc60305e9f9fdae94c2d426a7138cf8966b85c9a82482bd521d1056a31e1db04138772c9b073f83721b2a44d832ec7d9cce18d2e87af7603a5e52f4801fd63e2b9290b3e4babc806bfa1ce110f9bfe4a68add;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cfd407b831daccf226caa2daea39eadd8f43b3953070366197f35d81e630bdaee7689552d1a0e50c4ad1d542744b8f7641aa4799cbf981c6f4844c7b025aedef36c89b9ef0ab172dd27849d223b7a8d68d8eacd326766d2efcc19da9b4dd601f1341707ed0e0335512d21539d81e0a9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea2fbe466a8abe56c9982f7340fec779022ba4afae9946972c086dcff1c8b126ebd0f5b8bab6bc86bf6b9ea488c08275f49989d6b34924100e44a7d741b34640f150aa56e9f6dc85016fc873fc100395755a30ea03123aae105f9ea8208e6c6e25ebe2326526ba801b78301bf70dfdec7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h100b8847c7f9351a8503d5e0c595aa7d67444aab8b5461c718a9ac855bda31908f9da5a6a431f9326843c57336ca190f5b5de5d9a51e5713497ec5aa276128c9e62def8754cb8e3e1ad3313e77c6abc49ec8ca56329eb02142297c13a175737dba7fe9b23e3d7a20223b5cd4fcf919bf0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd53e6cc3433d30c57354413f243e57d5dde95d4071f0f2af44931e7bb606cf3cb6dfd18c21e3377399fd49e11821f9b8f39629bdfa5ecdc8715bde738ddc5b6d6e1ee06b4b56a60d24d3b6a42e64e0632750a42814c146958cb6413221982625e8507bbe0850d7ae713a3556b89dba4a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31e3633af1f533da1de0ecdd83341a01b0282b3014c1da498f80b2419f146b679144f6cc34d2fa99da98bebd3058819bc532b39762fe54b9b364c7dc56e9b1b4c2a3b3abcf9526408b1be5b853a0bd41610a569e7b25b34198c5d7d54a1ece285a048e973d053956a998dfc43d9f7ad2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69f8deb2b4af92bb2a816b84c592c28c5c97816aff4ac65a63c47fc49a8d0242c818b2b1676c5dd5b96d99ea230f8578acea1b34c9291bbb4456341e4e819a10ba9b398474c95de505fcac41f375b731e53b45d2acc3916414d4dee2eb778f636e2f0bedb6604993c50fef9c2b840c869;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf1bdbc22e5f7d6e0fa251f12d5001c03c317241aad5588fef65d1239ede0bd72031cdf84d4ce5f532ff7c58348442b6e2b7301dc630868c6142e1a7776ebe1b60292e0538a5b818d83f3ac81c296b5bd14741185ed3faa33011baa659d25c1d276a8a7f09e65308955b828aba2ac2b24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3758def30e66e5eed016a444e3d4b86a9505b91135edc0cf24ba6484e5f57e58789b21d2f56a2dcc778f75343576350378442308d3e5097284336bbc0a5e286d6d0009571714cf07ae75c0def9c16d9f2dbb90478d53254c867ac8342a191656290a42b4e49dcb0b6fe89dc1840ec07e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haffe6feaa9c9b81c7d6c0fb398d211bfb12fbae8a4ec3d4851ba177676307d64992908f0f6b419d258f9b2f4bf3351865aae79e21c09b1743d4e63c5e698969cfa2432326415b8b5844edff84e96235c76b70b7e6859232ab959c452939dabdd4c64827f066d5cdb8ca39fe3a9d9a5289;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0d46852c803e9513765ff668d04513ca410bc0940bedac839731ec65dd5b37601e7eabd98e160573d37a84ae90e42e0cf1a2262ab0e3752b831c066abc8f5c682085c149b08123d2157e8cc8dbc5474a58e4c1f66c59380dffd804b02253d97d1af956d3fb2939bf17566ecc930cdcfb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h189e168e5ccf66d5ecc6f9febfeb6af045f82b75176c32cd0ce51868f139a7edba45a6d9237c40648c804458a3529ed70938d14a737f495c4f37b5997fda77f382b470755abaa194bcf4c05f06ce2a34639b8ef1a35636a594063bbbfbbff9d498cc0f85ecc4032784e5f027d510aa09b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ffc3007e83dc3a6b55b22d031b2edb6b1d51ce63090073dfe8886436c7625c2171fa780ac9d4a310f634bdfe8fa7c4566253de8af730157f51c3991f99f2bd2801533f0d8497885b399710b3b938ad3d0c782becfe6eda30b4fe0065433fa30fe3203832e80fbef05ef9e1b2f2911f07;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc344cc09ece0a4a968a222dae7d6ee51af0f265c999ab2262590925bcac31e8ad158c772ef6bc88f2edc5c8e87a96b8a02f44f4ce0176131bfc9cf114f36904d8c21b1355e88f36b8f5d6f3e657707c16b435dfcad6e8f609561897b367cf91c2c3bc6efd6de8a31793b119c91bacd451;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5e1b538239f8aa3f4256444dbe9a0665a98f3d234e48e3536f92c8869efe6559bbdc3c0af4643722849bc761c9a7228e2cb1e9189289b7deb7c9b79d777039b4c4eacce78ab0ba8b5cde4e384e0087ad65c5d2cf19f7e011563dcca4a42854afa4f9c09223abe472f85b94470c4171bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa7b4b62e2c67a99df9e9ff16521f7f5a5423bb493b44f47e31d0b8058debc000a170d8fd8e53a401120c717872b3e993b024cbbe41b8f4a8c129c0d433db8111d42c8c80a7bc7ecf31a70d4b2c43cd81e1b1cb5291067e4f6a784ed7e802b330ff19adbe37b36e5ab01212a45f945d38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2636dab197c304ed33217d680054f9f9c7eb55875939e8b89e9e813f47f9b3ad3729358e7aed04f0aa68c5091ec945b0dd461662f9befae36532071723be1562d9e929ef3c66eca848cc3acf095151acc6685d8b46ef6dc9d7692b32daf031630d7e1ce2983cb4ff231e52481bad0378f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha554028a2a0ea3ca079b23206ad21ce935f00b8415e313e8ebd1baa0292de87f649ee673a11788a4766a84d23a43a19719536ac76a69fd3112c03e9adac8a46e9819234373b39241d22049cb188cd20c0789d7eaf722d26a7f09bad9a63e8547416030f41930117d56ac06e3a9a81438d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbf25825901f68545d11a197a615d26737f6f626fb683c3172a3693fab52ccbc88030f347b0fef7b197afcdbe04f7588b72e88fb49dec3e308df20af08cbc88d03a585ac30e88da23a4ebc37f1210e091fbf37f47c6443c8d474596b887707f1697bd1381476ea0315232ac2db631eef3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc94f91a1682902b1897937d431b745e64bc4f5120407eafb6e0fa7220d1f8937f1572c2f3f7ae135f3b997491c5fe9abd4dc2ce7018dbbd20a6dd62a9baa402183842c9bb8e408d8c1669859c291f1ca3c270b262fa79e8f7db76c411b4d3db65a986deb43987bf6dc59bf29aa7b7ac6c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h444070d9bb0595e6eaa167cd0297e21d38a100fd9de526fb13052d5147bfc3b549f192e4788ed630af63c8738ec3e0a61f1e0ca46adbadb2f3e8eb7dca6530823186739e167b584abf06a77d48f779076d889e322aac50a59a376191e6aa5e53ca4183728e5ffe922369ca8c5152f88ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf3ed34043a654ce6c6e24eaec935f46089561fd8d25a230c67d09eea5529eb4cb595b337735d350b6bca9f8fa4a9847b15b03dc5f77601d8f63f2bc5b62755d291aae97f4ea018bb53bd85cdffedfb460e1a3c01cd309aa2827ad47b375d24cc725291308310a6b97d68d29105040746;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ab0ad7c0f4a5696b6e91932fc37c41eb2b44676b00f904c389b239823ae646f79495e1223dd6d44649fc400e11d91ddd2a825c3274a66b9344e5b55679a9438c857af3568da07feb79e7f84037e72157ee17f1cfb4038ae89af66706185b93753eaf81b1db2c5e87a8094936b56275d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4602661a2d0eab14a8841c11fc6e709fa7667a3512c2c186e5c117dd6fa8d0413f31a1bf2892a9fbae338cc8638f847e0c302dcfec6526fe0cc5f28828062cea6493aff696ec6024dcad560330ee32a8e6eb180ba872b6ac3e3a21f3ef1db6069f0ca2ac482a2251180bc893ca22f3ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae290755dd77295145558a8e1bc1fc8441921135db8fd02379dfe401048a1c02f953506bed3203d12c6b789f3c8ad1efb46bb398ead247fd7ca20c39e7f780d713e1e8a886b3fced303b17eec5421898a0f58ddad3822b430968689e3cd3755c1d2a175b444e9db16eaced83116a4721e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h602597bb59794f4a52c1d56b5796c1c9facca21dfc43fda7423048363357303e0185c90de7fa4f5728f8972a7e501370544b3260ed41e23c3879335496832d8b70a59ed46c527331ab4456656c602f4b6a9a699ea8dea3356ad423a94e37f7eff06030be297699defe34084a204c8ea02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84f3f3b158bc260ce1d0667d44b9723a0bafe9c0ba43ddec04a55165400cd76619e28d4f3cb7bbd9c9e1f8ad267c5f59fddb50216813c515cfbbcbaf39afbbea74e73fa7505d03b19068942ff6f4e58dc395027254baea69b9636017acfd87096a8d4555887658dae4c20f6f6abb1554c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c6944cdcc60ab2b5ae810e91fc4faa95ba3c016ca7832a249148f55cd4d087fd768c9eb69e96aaf338b2b4b05896fab490299d2c1773f33c7228b8736e095a97e8b1aee49e6b6dcefab227eed5a1f3905e9531ce193da8e8695fa82bc081d7ff10353c2f3efe4c6f2e16de710f1b207a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8929324c882412dabd38103b2b86912e5ae92b5190dde1a03f88dba2efb4e2cbe087bfe5771a0640fada1eea2c839936617d825fafb8f0815e2cd60773bff882e907e4284341e4aff4a9a247e2bed58c66787ccce7efbd0e153eb2569b3b298f5e762c6b4e1250b31f358dcd2a8111540;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1242b7ade52b4ccfc5f50db5159733ffa2be38195e86254467b19e37e4217d6117427a0a65b237147aee8b4a76a53e3103680e1cbc8466d4fc1d7c1a43cc9ff613964e2a4f13b93204e92197b5f0c7254a72b0fa27b200c02ea4e19a749e65b7e43085ca81f0679b663c17661bbaf4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9683b16d0a5c48fc6946de9aff4f179496e9788014d05b0abebc48764ccaf9714ea1b65d1cda2fe5fe2c867261a8c028f01297e3cbe69d5fc9f42f968ebbd4a621d61ba7b3b3b7ee7ea5fa6ef7a95c1d0c3780944767dd0521b7a432f12fca5c82f207a649ea24d025f3b23dcc745895;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cad5dcb7e6759e8bc77afe395eb022cbe17c1e8264fd1c246578b4aa300a6858d1152bf18f0be2cca76d05252e20afd361942c28c280afe552b6ec7528a6124cd72660a43621a9e7fa0e28550d9db9a1131101f5cdf9e5b00d5703b20eb7fb55fdcf22b5652a08ae3a44997ad95b863b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92726230e6a5de337750a07a24299488869dd32896aaee3707552096c614d2e22147fa602a0e1bc964fdec8dc48928a36a34c78f460499d7e752d196d156cec079fba734874692f7e5ec54c01eacb94a93ee9f270b8a92c2706b507a95a492df77f27fc14fd7ef5ff6d37c06383344714;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3da59e34c098038777dc2d451eca0020bdf1589ebed4629c06f1ad9e67b77608bf84c9492b6af5c63b04148e58cb63d324650056fd5572d08b1da5472a1e1630e4e6053f2f4607a6967e34286039beb2314e01ab5300f933e90d053435335909b4095c0ef7493cf81fb5c0f4b5d742c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38eed7fbd047166649690d779d12ee996cd54eac36adcbd01cc77ad29e09e24d0f0bfb9eb8fd8296d79b76ac8feebf1ef9fc8fdd6203d8e90b69f232a7e78b6069279d1679d402271294c35116a4654137e8ad70159e0adda0cd46d7ee251f3f836f0305eab6866370c4dde3016a9dc35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86b96afb45221d0a620163b233a347c611386a04c97d88a038746b45de44bf8870727fb7dcc36f05d5fd7f39b54fc5447d873702bf1877fd274709094499a1c46bd17a5009c540031fc99536fb73bd9aebb9033fb8f63310a1fdc83b0074e76569bab9e8c434e8fa1dcf60699d3b495a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b7ceb575a70771a40817a14fa59e376701232c901726da33b306596cb45894b60b71b6c41922865f5f9b28dc06dae195138d0376adb33a1d91ecde70dabb29df7da1c597dcc24a9a5e5b84c75815deddc805559515da82fd561a190900076fa7aad73a85648f3e0faf3d85e5faf7ecff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcedb39d68beee1ef546f4ca79d56fe4247ac6b4869f19a22bfedd4cfee73d8794f9a1a0da121069de0d9534bc4015f247b9affa3ee7cb6980e8e9677eb58793685d0cf7ba10f22792f0a849b26afe3194f145e12e537df9726d69857b69679c0f3fbe1d0d73619a6501fc5d19554d65f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a52a5c83c58c7fefe6110663dc95640f142519866c560e16792d7bf49ad95122e34436039303f827add640ea14676c87aebde0017218e1c558e1fbb875b64b5498173156c9a313b08a55fe0f68de1d5c731c8ba2694273825a04d16be368745d2d8627437a94cc5111c99bc94e82092f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h980c17a49dd400bf78b176df449912b5fb09e6ccf5f3626e3720a440aa36927d9d7088a703463b9df5c0cdc3907f06175e7d4338dc15754bc01a8a618deccb12e54a62242fbaab9fa699c5dba5d84508cffaeaf4b49534452e6b70f036da05a5db487bd9d03b9c2aab0c6d0ed70b74c1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b16a9ea6fc52db5a2f04ed1839391b2d144b731fd346327080bb6293c5c7fc378f760c0b4fdf9834a9336cfdbb001d59c418e7f6b3a6a8590be43ba8c9bc7239bc28eb0a6b2044c45834f24f38a31af39f16599526d5ebff3749314139548f5487ddb6222cd229d322bf053018ad7ad0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f70131fd3f66f6dd5147923ee3e8c317e19489b4fa5023014cc77af7cbed01181bf53c3ace385bd6fe9c59b8ccbbe49d26ac27c27124d748dd9ae95c1753077728dfd8458266c3181988dd7f9dbcec86f2fdd21cbe26210f1274a14c7246c5c7461cf35183bef583887479e01eb1a68b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a41e5310c079596ee8d6d8e7ce26714ea6e29220d77ad2857b795846d2cc6b284e7229641e4976b36dd3196e90e8ecdbf1a7a725ea15b3e3ceabcca0b85bff3635f178834768327c65f7ec6c3976235ab2a50834ef300a8e417f0f38658dbdcd6d94ca658742d8c72ed47f830e76adc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e01a637e8bba959ac76131c9d7fbe0b1c8d9233e7edeabdb39dfec43b86f476f231a263eb54cc94e1aa554250b56b441fa101a3fa744ac337381a92d90d4b36eceb341ac6527fac97e26ebe746e2545f25aab4582b9a1db38a92dbd06ebe4b232d82fc6c218ca62f3ded70f125a63429;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ce15a7da38c90d8c60cc5c4dab526541a538ec8da9773d3120fb0e17ed9815a42af5f30701831f6148dd462ff0f5f86e2daebae344bec94d33b440a487b34e5b99b2c688f6ee6e0c0e2864986526fdcd2e32e7d0b13a84179f0ceb608a0210ec16f6311292e09a8f88a32da951eb8c6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdfe7b5b6eef7272fac632cdbb6c6e93fe899eef2e85fe4a2ff6e7f07ea725ceb9e570ed4be8f22c47ecdb11e854077a0d13654b6c869749bffd18c79f2e4320196d7a39694363fbddeb59be57302018b91acbd5534cd01d06991c21ef2dd69b7e6bec8c8e024ea4d1a6c3fe40782841f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34fae11077580d2ac528ca60792c2f879ddb3d16905dac1bc3703d17882b5259dbcb6eb8c285fdc7e4c653c4d67009066033dcb26b477ceb724cf00e6eea1419ce02cb1477b68559a7b581a6f98e39c2215fdbf7c47a69b0dc07e2c9ee8e7678aae6411acee0c71db1980df6a3a47313a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h599e188ca19088a9db3c5f39c88ec4e90b8a0f98843bd7bb77efaf4607b1beca7684bcf51951eb0b8a93a82a161372c3a072d4a0b8e3ee498ad2488d4d3de0405b04dbf48238d9219c3b28a03fa85b36ea4c1164f8159ac5e696c185a4c8aa4fae53a7a8b80d21cf1f2ca2b63ad525ec2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fe4454e8458fe0caf165503b241a7f43e468fb41801602c0f6276124e879a72c09fd8d70dbf37b7b55a4b4a1b8f03f3cf78e5132b6aaf5756332e59c64b2d755bd217f418c8607bdbdbdc04893d059cebbad98c2831dd2104490bf785bd3522f76c4945dbd077d30fc63da877ef67534;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d6814a20e14765e533fd56838db29d30db5744c39f06ebeb72eb1c7042ae1de2c976c9137b865790bf8d7a942858120e33192cafbb5bfcdc4fe3cd625e8ea72c9b0d36df0a1a94f437b49a49ff4e7a04010055b746ff970955ba102bbe87035a6c0ed7599bd64eb0219b6f31d7686bca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6cd46eb9bbf0f7e3e99c5551e33e00ec98c4eea6c71bbf3f0a932f74f0a477bbb1d8daa382db99dc9f728fec2203fa9dd0e8f5264bb17258e7a5d9c13b5c112924c0087491b569a41478034e5fd56420d2fd77f82743c665db35197fdbfd3fef01366ecf1e005ab56fdd9dbe25e3c506;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fcddacf913e1ea9b910730af64254b6c0983dbc31f9f4c8b628a210c416f2543eaf0b19a6e9cd85bd2f98481d8e81f3a8fb3dad64b1619b5b72c6f4cbc94444404cb9f07f6383dbffee12c4f0abfc6472df3205fdd83b268a311518c2d823c80fe8c9b53b21a6ad163f177556a9a1f1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7dbf2b22408c77f930478b8e23ea993c93d105cadc54070a788a6c9c9e40cc119c2ed129d53ac22e15c125cbd0ed021fa534cd6a1ff4a54a5f080f24893633732076983b181b0e9b7496dc4242a827cbdf10f19b886f5496e1a7bd84d68bca5332d89d2b4b9726592746e439ddcd6cda;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8370fa95c6214f044dfe40d063716b48a7bcf89847b3aec70ab3f66c8d50ec9576e1fd53d475dd934123dfd83f42c26fff7c6dbd8f8a9577bb2ef2335088cc795fdbf9881e2103379baf1d15ba09e4f31702e0c2bbac9d2a50696921a6266409c9af5cea6ab8033d123b9a7b55007386c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b936f7e642cc9481a5acd81fa53a4915ea8f640d8a4c5e95d81346cde967fe7758c6f1ca3fc6914db879843fac09f6162f01fba7fd9498f4bcb168a5da4f8eb62096f966b768f67bfeb8d9ac1a54f3e8e309994e284139dc26f2b85a040fd20b683bf8ca6d155ce5b90088cfb8ca035f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7f22d8f0fbbda6d9dfda346badc0def0e6adb2e4dded3b73518d232ded3e5c150c8c4fb83357c0cc353bc06ec2441a6811db6f7b3a1fb7bf76d2d01973a0ea2db28cce23b5cef0a36279145e2a28ba34eafd8137f81aa622b99ed7a5c18dda1d2608056286387a4e401d2cb48e2e89d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b3194fed7c5d1be8e8f2125c601afc9738a9ee6f25c28f8f08f5a9d71395b5e43a0034492d1a012a88e11197c2d738ebc968302c63104793c3e7a444dea74a5537b04224a232e3231ea1249f80b8be5f9bea3256cfb0b68bc82bd8190a60ae86520b3520aabd184764b94eff4a3872b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3543476b01b9e20bb5e7801c5758b758642e98cc79ea8bd9d812080c2b580015c6b837fd5dab8cb9f352407d0d5f0d4ad8343c15d52e07973770525971e94edf4acd8ecf61d99ef8362494ee5f8c4f08fa51666a121630df098013687676cca04a614de05db1ba8aa78aae53d853083d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c6459e9aafc692442193453a206f042e007ae998a1ee15afb8c61dd99517d4806064e6da306e4a2171fb5f396b48c0d5bae3e631631f6a452ccc3f2d123a73a0b29cf3847d0f884230def9e996536505dd9d125b2e87dc6a4b0b911390573be2a16a79156343351c1bb3cd5ee50cd27a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20d9a838e37fa20e72b960fe843ac8130c91be7d2edc5e617eb0560c73a8ca82cb2bf3e17e897949f20db97bc05a22eefcfc154aea9198d4786ada6470b73581aa11b8ad2eb4fccdcb636c9db7c6f52b13eff55808784c5ccc294e5ff7b96c94e2dc8017c51646bc3f4c51985ca95affe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ce9f2bc9ea2b45b3624f994d02be5b0f93e77119e37a35383a61b8f92e89a4ed4d92569ba1e52254ccd057b30317c0d448c3e848842159c08e83064ba7c7031f8194f119bde850ba3651cea350c38efea5edd454d8e3711618c1dfb724dcaa7ce1ad7569d2375d6d830f83e2fe36dc77;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2cbbd56dc04a598697be2f33685198243512ba955894a30012ccba989901c97637386f29ae27c322770bf9756a156dfad645308d2a4d730cc7fb19e80a02e1306c18b7195b8d3e51a71bae6b741d06331df7c55dc7a1064e207cc1f63ebc990e9c628099143c2679b5c3c7e65422392a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa4dce58cbc29c3ef932dcee5065a3bfb0632d1a4574b35ff47bbfc218952040ddecfaf52f195374dcf1aff4a714f6da30120eab60a5350972083a0cf354ed80ae96bcd1893a2755b2e09f92e29ec5bef7c7a4e939a5551b0d75cabd661016210f981a826b902639627490476fe0a5238;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9eee125fe5cb36d8a7627d7f82dbea2d7f29aa5cadda927d31cdf10949a8bdfd56407f1254e30024a5b4e3ca13021d1c535a413d28b1e32bd1d0cf2f82e8724f749394a90f37343e40ba33b603c350a91186449b9ee35e407f8352d792bc190290adab9954542728c34cb9b785453b98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1df5d12a6cf6574a2c0b3d29a6789a3cdfa2ed4acc78d1d4d5fed990e829b67e770ac6bd60bf40665e50782a1471b30a4ea5aa88d159e1a77eefc3b5b3e6da6d708dd68b2197aaf9aad216123bfb2534a29d062b0ddc3c7e7d271dcdefca7053074b3c3305bf147e35ae4006d623276a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51a07637ad39f0d7e219c87f0b66c54fe1155de7a9cc1017db97ef96506dad8a294079afed380e35c27d1dbcd2844d35e6bc1b27511554fb5e1338b076a9ec95c9c94172fe8836408d96a696d87e19c94693b2ae26862aec3c91b0582dee4cd54d1017e0b13edb80b1c46fcde2de1d9b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h394c6d0db450623a5024b12d8fb92357698c2427aa1ec8eafab6e3d25c1781dd07edb1a9958fc0b3038272a6d0160f3c25cece70b7940966e62665b79e630f5b3ad58f38b98c35586a3c66812bfb06e153df9f53db3f76c2a7a6c869664b2534359b324f40f5e09ed05549d3dab18533b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce5a6130f7b550a03ef8ed9e3c43d2ceb4d6c845d0ab12b00cc9b4575460ea04c6353ddd5a4fcdcd6498ec524392465b9318fa260fd9d94dc1998090f20a788bca1fa6cabb9e392a7a3bfda2ccb42fb85b219e55fc6b63286dc27f51f3c7ca1a81007a3ed91c9d260ee0521fd6ca546fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e8207b3f5f6d00795105dd34d1a814cdbffd154ecf8ceda707a7b470ee8cff2637a60ccf18bbf6543441aa64cf639a7c11134a209c1bfdd63ea40e86fd1f71bee4f8f0dfb696f44b52616d9970c73fc5100c716a12c9ae01cbfe6625c62ba5591eef5e9f5cffaa3a3efc8b90beb3ff5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5a4c1df4a26c73ce1fcbdf9f6a0730f71bc3bb30721a5ad15a9c69c0995ff9a4fcd8b55baf36ae7d7683e983ff9c5c5903ce941ee2f8ace615e65a6b3255dff1d1ea247234e9c187250ae2be486b91afdbe12aa642d4bf57ae7b1f440652cbbff228c0fbccdbe97b642af41c10cb8327;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467ad411c20a803051dad73f67ae66149c96672ca4dfb128eb619c0a1218adb94fb8f6243c300a17ae326d6c088b7e051367194820acda03a9acefca5a930ac4ef2da1cde35ad377a08128a54867496296c1e9e293e13874d88180c26ae85d45f76394825fe5b1a1f13aa3c96aec04fe9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2e8343cb95bf8d37d749e2fa98645ac955e44adda8f005445830b50802fbf352988b7c3438fa2bdf0916317384291aeac280255ea71e94e091fd7aa37de0d9863414b68367f044a27c521a4451272ba494adae8b2d7782199162b782051cca0d3e6819596b36ef51831a667f2406f66b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70fafa65224efb721a9810a5027e3298e0bcd57e075ecc6c8340b62de9da72ecca5fbec7824f89a58fe40e6c82803fb881ec54b337d2ce8775da7575f9f7c3dc117626ba3d9d875d921520cb726b847226d2c6a491736e791d03bd1392259b41c7c314f2e4f2dcac94302770c9290c57c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27639bbf6e0c55c7c71f368a8da2f61e6e83aa8b284bc845ade61c063faf3023bcda5f0ffc65c09908e70400f34dd05da902686e4be6ac50854057a93d3be790226bd7471524970f66d9c20e7db1071947fff56813a699de8f656b403402dedf649dec08b3d19a633ee0913b81edfce55;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7914b6c056e9852f07b5e18a5f3075b50d2683a158eaa71f2709e7a74efa8237617b819f4a5e9cc255ff3ad58a1a4f033b41c430ecb362547956d084037bd3cac098cccb860fa412ca921f62662d3b1842803aa944d56deacd3a0cbb876eef3bcf29db9444b3f125d148b912b4cbf21a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e73ce0822a2947fa3ae2728ae966a3a5e9ec159a46999cf7b44a0dc00738660d7ab552981487e838bc9039f903242604e3ae092d43ecdc14778c811a837cc6c2d0799f92f6cab7e42444610a1fef1298b12f0fab2a136051b470a5a304fb5e9cc36a8af037a5eff1586e7a7dbec7161f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc4bb1093e04d5d47afb722e2083de5220b5681062d6c1adfdf27e530c2f9ccf423cec18f6d3c8d5ce2902884e4cf564f9ad5d86bab609008daa8472765393bf8a962115320b9ffdd7b8310f946bdadac32d7969df6db6de190a51e39113b9133ff7a7253f899c5413bebab98fe25aba2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4a8c2395fd4e11aa12c008da99731c72060d2ba0cd4f55fa4a04edd528ba1290bcbcc0f5da012f2c42c72a315674c82c2553214419fbdf88610d205b34e21347961a394b8dba385ddbbd50b290491bb0c6f38f5101bd2c84f26a9ccd1fee8188a3e258f789266f3f9c2d9aebd308a86c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41437da3e9c927c289cced40f8f613482244eecd862880ae7322455ba400ce52157264ffd0a9e9c6ed41bc2a61c0f7416108d267ece73e0058b1ddddc58cb58e45be6064a39f29f1da627448d426d6cdd9ff8787cee4c7dbad85e280daaf493fbe6faf53cdfb3fde1ae00e970c37c9855;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d8e4ebadd1d7718ce9cd5927b4020cf08c8fbb9811cc2388eb8b27b7369160856452b42becb79372432ca1def6549624784e75f6371d151e9f56740f11c6613f4f5d57134491d1f378930e5015e4ba6646c3054fee23a15480a9af98f8162bd3b89769ec19c2f1c8c9a30b6bf9c28df8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38aeb3f71e9632d2d5bd3c9e309a07eb2c9589a41ef80a841f1d6136f6499d7dc1629cde1f698277a89d2e94291092e461dcca276a1fb79beac57f0dc7495ed8e5f9669a8bdf7cfaf57b405506ea5462fe1d61589cb8302be1d0be2590e8140d676171ed57e85dd5990ef86943bf5e15e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55a946b08dc7ee710781b1eefb17f8f2bbabe5bc668c335d5c66748d9c1ec264c6e7573f2038f8a406a9b68c82e6de3c29e7d650d2c558634121d83dec83c4fcac6d2f321ca9e45164037d05e1ef95f9a2d4520036e47e37223ae2be8cdbed15033a52c482d55e08b41486cb8da73d44f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb38211ecce205bc5f577b494f809b83c00b93b369eb3880b77079c8b6999571931597b472d0512aa89bee40f5429b476fe27341ed25391d68ee15ac280c28d1a904752aaacdf67f1788483bd4bf17aa2b5ee3b8fc53413985873c135c90d381d324a680f7d2f3e03bd0bf34735e4b2bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b90e5af4618fdd04493ec63c52378d5841f3f787c265964be99380ccb4e1c13ef360f70e7bb4e66c423738224771de48110b3cc4fde34b722981cb0ead7a3c5b64538941ed4a68bf7e7af00ce5a53c5098ba66a9313b9ad16d1202aefd452d0ff3cbfdb9dda8089710acf91de4c58b5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h771919ecb95733257498351a1ad5a85313c5fab11c4a9246d936316e92caff2d4ee1cb7450a72796a962d9103de828b03d462b95123b4f7a66d68644a9ef3996af1636b2eef60cfbbd8f651f2c0c3a1c7f41c1c3d33fd0224ad53cd3dda54f2b131ad072ac1ec1bb422e6e0ccd5789c29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3310a9de5ce3a16bd35946a248bf562d1c34a996f782b8c3f6ec814251513f27c78b94811e404220827b25b811d481ebef20e72ec54b1401aff58779eddf2d14bc60a680446a668936a29de618935bebc994907ca4d54518a465b3abde02e96b97dfd296b2bcf44302e42af2dc5650b06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9801b421ad0946194d6cfbfafaf834dae40ff5b9126e92b670d0eb29e90b9f9c43673853486e3b2ca9e884af2cb13411155fcd6d681d414aa4bf0e6900d59d8e2593851a23eeebb7086a0177dc0c4d090f5d72c721a36218a000222c6e13c9e362eb596e171e9d2277abd35db67002a85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf750eabc1fe9920d599439abf73564eb01b646d8d5b9b2abea56adb0d651625c64335dbe341e153a9013ee3e199bf76694d0b5367a884d4bc542d61aaffd1ceff8504f99b3208514a731fbb0f0bca86dcf5a78afdb4913e761bd37dfd4b27f81ed763380d02114e9460c2c7293ffe19e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f134529aa00f038c2ce1489425b34259a866eebf1c6bdc0ea58e760c3e10d0a369d6882d66e2f3609c4d124916e97b54d172506be31b529cee98c671c1398de351d71601e072b51c95be47fe5bff14ee9e8179e40e46a90b7366cf44c54434344c5f5ab3fdb8012e0e5ee06a0a1f2af2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57bcd195c9f3f60969292f18b79aa480e047f507be5aa97a6ec9f7ef244746dca5fb8dbef3650fe643eaa3adb5cfead33080e7576bdf738972ae7cbeb2b022d8b0880ae51ae9c0c0d97645cb5db66441238c854aa2ede690b651a769b3b5d32bc069d21c1440c796996e7c4caeb6f0c5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3a85078b9a243f446d2ee4a1f306dc9ab6262a997611895262bdc49ec52aa4f97c154f282cc844671bd7a78c5d734028e966738c5795ae001a37d1314d14fe34f0eefe4738c418ac9ece77a7811bb9e2fe8d62566f4cd737d38fd5be6ba91ec73fc049292c5d39541aa03d7b25eb63c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56d0e9ff9521b3ebec82adb054fdf7c4bda09edc7934ead50a98c65568df5868ac04902b54d520a8c7821f2b0657bcfdf072e14b6ad9027296e5fc344aa4883ebbada69a781492b156a3ecd5c4beb738ed8bf64c63121db18699c174c3bb49ce0d6185ca638e7c6c7c1e70e8327bffd62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97b3e38e76152f1777f737073b737e5d1eaecfefa48af1eb4ae8f7b729070896a27f46c77c65736345e38ebaf57a0d08ea7daaa04b37e73790194174c24dd3f3639ddbf88439f9aa7f766564be84c2b19b1eed888fe1ec68142993b45698bb88b0e27a26b874fbee04ad9785e8fc052e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h744c7a448a23bf8fa7a4c2d045ec8163a712c9372552ab815ff5fd4d172c31b03667d3cd57beaa96f726eebee44d7a8dd6a90ca9051db23cfa34aa5bc578a52417a89a8effbc9165179a3a1971a9496166fca0b94dfaca246a6329b5a68399371f8579b24d4f4ddc776132d975975a799;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1680ee74b84bdbfe9d474c39f2cdb90b4e311373f632da91f2bc8a8742c9832d13aa0e01facc8cf3c6f7c487bcde8d2dce9dac94b593afdc4392db85e798c0a7c97b722176649d692be367689c606724928353c8dfb751c5d0b2270e93047029891c7885dae4448f3ea514eea5462096a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffa8a78efd684918384dc8376334cc744f16b471e0509a3129d7d9ce48c70257983c89e10eaf04233f728264355ad244101347bcc3dbccc180c22baf581c08169b90697340060d325e433669e60fbcc403f591a7c6f37b1d125a681b1f9c5ad4b874f94b16fc76dac9801ee9597fbdd9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66f0b00e5d8ff9d8b72ec0c8dd59eee1ce82ed271b46233d62b9c3b12fa9881dbd2e7d77f4ff9d12e7f9fbc72b494ee6330f5ddacf5fab53f397833d6d3bc1f3ca816fcd10814cc7d4bf85be9c2107602d1edfe2360159e007180cfc43c8c78bf0254bd96abb08df25e262e838029477b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea06d0c67d6efbd1311c38ee0a9103766dd43663a101fbf64c303346dc67c6ee11226f2a3cb7220913a71fb25181a06ddaa544286df22021651916a476e41ee9ae5a87b89da866bf22b4b7f53baafdf557b5eb27b09249cf0ab2ec5c6a200e61e460580f9b6a700b0c53b59cbe0230fb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3373684d0066cd77069af464551aca24c3a265fa01d22afcd096e2dec9891dde4fa9f5d28a1786aa8cc164594fea2233d0e0459703a2aa48f13ab946f25310aea77a5035a08cbd3d3c610d3924f7753dcdad61576b54f038f0d67331f10280ca02a898bde5811eb4607c3d8314dd577e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1939c68f860f10c176588ed533a237724a5df21b719a274416c600808c35b4ef8dd152ab5369a8bd8a7a09409a8131dfa240478dbb3dc984e6ba64263b5fc4b085260c77fd417b4dcd6f1f76ebe92fbb2644dfb30a9b9fd5a8bc2f2c89c962f3ede9c57afc1d019adb81074ea1aff1ed6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4228daf9c69056e3afa3542c168ec8ce6e73e831e11c99187f14532d53daca1cd2c63158a5d2e879f6a8ca9b1f659c9c62b490c1651335da4207f75fce314f82b7766ea0be97469d97ad865ec4cf0e42675e4bd33d2da77afaccaf412c1cb4aaf13c33d0a6ba54251f184fe4ff74c32c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24e7bb4bbcecaba58a68419776e8a44d04ed8a16d84abb0d1f21abc358dd40da8be4bf23cd9dda7dc60b775c7438e7c022c9c688611d3521d64c07655ca9c43428ccd05c894da872007d78d27773a2eb75529267ae2b27a7cd7f9414896f0b2828b24b6092c01e17232b210ee9b21199;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc80caf64588e45e73073ad49f3bd78970cb97f9aab6db09f20f563c7df3fac7daffc37c7d761bf69a1fcce599c32218587d57f9661199da42919eeb04949c0289c4a2976d00a0202ffa70edd082de147f3de8f6c85bbb4b8ebe76d936b78ffd014d7c3ab0392a281eac68975857d204f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7947d9c98fad398c7e7594c0f6d7342024ecda802f8db2ad181cef54aee542449947cbad2c267fefff743afb2ebf1966bf067716fad42ba6788b2ddcb2a556ae53cd91a7477f3c9c8e76633236603a30eca780507c44a347794e1345658bbf76de2e9ba5480530b73536b3d7272c125a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fd437ae02a7389f0fb1891616ace18f00ff19147a7597205d9d09e0a77ff7ded04492028535dddba57ce09b57c86e859133326132ae35a639e1550d7eaf67e4d2322fdd68a18ec94766d9ca9a7851fd1ca9e5ac3de6a963f071754122c08f83d939847d93311b7eaf55a2df14cb6d3d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d38204c7e06549ecfb6867625f183324b9af1ad32fb96fd9daf22fe9949fa3c129d52a7197fa85668f897d6ecaab4e334051c9a6d74efb48b8e0059676f946d4e1d9dc72c5ec42a1bbb00e5b534a936630e3951ab6e3baf09e6f1a45cf6a4c18015055f5b56850936e5b18b0177ffde7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6bcabec2334ea90a325ac2297dcd59af3784bfac13f9135e9502872d9b52cfe21115ed150eb7f69f220967f81c5f02fd1e7ccd12fd60ee1696ff8109ebb69a02544a6c1e5dd38020799a12917d6db480f4c9c5f14ade6a2f7d9bd419408bf2b9e8f05e50e53008874a81553bf64f20ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc17319abeb654b081ae54c7a1c22821ef644bc385e416793ba47762e88966cac9d8459d3631ec5d9d03fb23b8d693f25b0643386481df46529729127078e9638ef789700cff252c0bc56680d5d84f6cec3f50ff7f4d8df2726221bc40728410faea3bf0961c60195dab1914677a2e56f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5d91a0ac08cd8dd1cf660284eba3fecd4df0d60c7e50fafab379d4ec78de902d7f92661d90fda7d0615df6612f726ce19b6d7b6591482d1f751113070056fede74b2f1064a7c1189f7f450e68ffa1e744eb9110a0c70f68b1ec3be81e0eed74691e2b51eac38d0a5a6f98cbb200e11cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42e1bf684d6fcd16d7cf16bc1995a958e1adf8b514df1370cc55200e517d5bc6dd6202fbe2be294602d90817af4e7e43ca3217d5e68da642cde879049daa503a488251efe2b9cf46bb23d6e99ef11ba0e454314ce626aea80d7b2d087a879557c8345b36c287a91089f374bf8186008e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca2d507f9629e4401ff66cfd7392bcb4de221afa3a740f90afd0d4eb1d8e8a831bbec49bb410ee8031790912cb37ac07fdef85c46847bc5149aa78be0edfedff5bd7a315cb4cf5cbea4002c8db945d8801fb5be727a8ed26d004b585395f85d9ef5bf657cbecb57453dddd4b939bf14bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71296bf5a877fe2450e33a67bb9e388bacf8623f7ebc4ed974bd133361029530ee0262d0db04fa44dce245ace1d4230cbd08bc31bf0dfbace3dceee29ec150322c83ee3017bcc2ac165d54b00af8174e1dd3265b73d5567dccae5ac916eff921225dcb5c86361f65687481fd5bf619df8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76f716db34d218c1e2b162d119bf5527ba51671a883bf197362e4568a8038b6fd044cde332f40d4a97db8c533fec45c8644ebd4072cfda4be16508ad9e2dfcff62567d78cfef545c3e7ecaee26bc7bc88274ddacc81d579d96dd5a9ecac3a918e27e76265c0260caaf52cedf4b276a8e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd2bde476be5973bfd97c2e069254df7f41b12abeb1a251dc755358416c8b3e2f646f94c2cac5e13472b3d5299b53e8cc5378a60c5f00874f3c6d12ef943b34c1e053ab46d086e6d785a9e8658d44ee05c9c4cb03d7e31b266f17b0ec22f227550f0c91b9d3bbfe555012fed5ec98d53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha527327bcbbd57922d482d612de5f86e3c2d972a0d50451ef13fd4fda813888a82840fb9dc593b99536237e74aaf1d0b6fc72441029d8f5e67ff31a07f71d81cdb4c6b10e6f15678fc616cf41cb4ef289d2adbf0c8818abe818086cd01633f9134a66535ccef04c9172ff4a57d13d407c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd10cc498145d31c2b76c6fce1f1159ff211ea2dfbadfb49b4be103299517fe795f1867177178df870fd7e5973daf483861a0e3e1db3ed07e2365a60f1ce1ca529666799c0337bf4979d8ad220b89b432ee7a5e781b4ec51bda74db1a90d8efeb84bf2227f3e9f384dfc765be30b52f524;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc72a73336507aeb687e4b21555ac6c75049e64a2ec1089ee20c3532e4784c0b8050fba2128f9cbc692a71dc60aa37c008cd54ae70fedf29ecf2b8cb6acab8e8208d0c873608be0909b3970f8bf3f26a0d2875429c0d489747a24138e92d89415725ca45703f1f18fd826928464cc105e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b14058e21d77c74ed710390ce48bb04572ae213ae231f500adbbd580b6aa86ba98a64ea1b6dc0390b8dd4ce86cf2bc07b3d0179422978f9bbb27dd5102084bbe8bd6b382b3251b828e10dd3918ac913922232dc8a949e0bf021d899c1ac8cd92cf3a8d5f1c62d12528a636230cb899af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc87c288521577e081bd89b803051ba7a8cac7091e49224c84e7ec7cc1678592d6bd1e06e90557ba1cf036da3d37af13691cf37de6a05cb3667579e6799a82f6cfca8ce8a03d57bbe96205a220d85360808ba6beea5618d381c40f3edfff6f3cbd3432b18d35f981dea7216045685345b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45409a0627b7b34b7392c02ee619179e307927f40ce6a7119dfb901ffcf6bafb3fe4db67626583e256f6252d3f71ee7e1e0a593a972b6f2b9534b0261d1fa7cded5889be51d38024e70644d298a53d5200f0ca7fc712a0ad35e24fbd59fb55d5b239f8ef49ea633f34c30fa6848025ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14266ce60e49bbd69d30d553fc4f23333439c61f38f88c4bc64a3a44957f6f7e14d40ba914205e25c1c23c8295893cfa57b40d589a1d166c9813cb29efdffdc7b1d7ec6a1a2f9883698810af5d340c3c8bf4c7acae5f4f17ca0ba10743a845f6bdf567d82c60e5bb2eef577840ab17595;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96c3bc9321f821f71d52f69c7f718a0c89f6917a26589aded7bd41066b4921118f7170e6089fb1cb169f6fb91b245468920cb5ac360c4aa27fa2cf8c630fe068a3c496ffb1041f775ee69eaa974ae0f98d5a9d1c43bf832dadb5b0bce43fdd55f6d3fbb160443700cadeccc9fe144e9bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2b8ad1353bcf8e71f9e48b02db01aad6c99e7fcd701992f2ea5947a53db7a6a05cb39573a3a7ad61162d14d04d38bc024f7f883aec500344d51955918c593dd3d6f279d725e34a70e75f91c28bd245b1516af81399c7863db2b5e7b00a41048d9965d0ba830209dd64a8c837d0b7fc7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81329bc819c3dfae3fc48472d0dce1483ef2280861d85632847fa27dde400836f81a82cc7cbaa12a597836781b84e33af7ef5c67f01d8c6a368a28ff40b5b1bf3ad7e0b81d819d87581736ebdc376a8c35cdec93c2edf96d979ed057cfa1d0bd0ebdc8d724c90b94a2e8543957299b528;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9af8508b856511ea738c30cdcf4aa3d78103d27963550190410ca0955edc736eb96938a92c88fc4fc5590f8d0449522770ba6253e3adc8d3d1096e2d65b86d43990fdc5a94c1ff8057187914c9bdf4f4221afdea17d07a92f4cc8af5fb21c23d5e590eb17aee93d1894fe41de8c338bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha01b5ab40c83048dcdae767cb7b03b4c2996093f618e311e076340358a00575677ed237fd202dfdd21ed4b76f449fee77afa356432598be4c4908dbc59262361cc61a277ebde83d08dab697819f5bf34904780b0cd9d54c144152a322cdff28c712b45657d4942c59a5ae1c49620e6e98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24e177c0604a6deff0831ca395630ae063e44bd237ef0a9ccc3cbfe87a71cac1ae778f8a2b7172e7b428f71847985b78eb90d4f20b2e613648a6e6716672886114e004c72b08995a1e9307f0a72a63324f440ebc43eabe70a4b78ecec5969d4d90d6a6f4a16c1a8074cf98bcd74818b49;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcc1e5b29298fecca91a9d66da89a1af27de9ff8af0be727ba1f13387d55bef0ae7c14c16380ac7da691e1f76ecba372c7558e231b518b89bae61b7e0538144060a17e12cb80cc20e0e70b02dbf2074ac7a0b3154c50f8294ceb9b92348a9be85ebec25e2bcca69544227c96ae6525cb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h299ee345e228b9b166ae8966471505e13dd38ffa21a38c275d3fa2ec9240a93e43b9bcadf81831340425e43d6454aa5b359e094128c968e017e7c49ca079d29e5cd1ea4bb430058d9f813734fec67eeb7b0abdfc10d113faa5ca5095896e95d2cb4170004109e80ad585d562c5c26e57f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e5da198f830249c97e825350f171b30667f7aee60e3dcc6c6e5477f41d417914af5ee0ef547e8c71173b480a19fcdb5640069e1233f973e062de46b346b6ede6365e28ab71907021616db3c6ead8d9774c2a81c9409e0fb4e83c777e53e8fa9be518995a54c946e87b1e7d4155579e1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89f633623a39267cc7cbd3e4ff167dedbc4868031365d1a2bbb81b3cae81fa1cba673b157cdce714f528ce17d42d9224643fd80ebf778e890f563d7d76d6c9e048f60f53ebd45b9732c78daea693e911ccbe5bca32558310d12692e2cf335a75be8b904ccba2dff3d1d3bb40726dd1e74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he66b81830cbda31162e370edd1542273727eb5a2aae1561c94170d10e45f5ef170785c52fd24b97f796130f72e736c34bbd6c9a1eba7a6ce7e2e786c4c98ac0611e80ea2bb05de01c6095a8b2091db539c7ab78e7585ddb1802935d165895fe1767a7acb826c33afa87cd8a59b756604e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cdf522b60a79239ee9f2b09d46fb4e6bf8f3de70de5744050c3fbb9854ecba1dd5a38b640dc4d4c2b642405e1f6c9c29505f50773fe06a338e2783620eb55e01a6aa39cbf77cd85fd30291e31d64400be13929fe8e2e37ab04b5ccc6a3e44d24edc7ae8d443e2d53649dc7aead63e1fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h829d12bd31c3428b77d215fa77724b84ea205c9c8cafb3e425b8658e99709e2ab10b03797be4ec539d4fd87ce90b0927c292f4eab0fc9bb8d9edbbe1f5fe5e84a291003be97bc7b35385cd49f4d8c4a4efba5acb4063044b4473f2d4c2cc671414ec3119171e6bdd991785af57b91d632;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h991f9ead675a5e49d1d1556399afaf18d5ed7e00c5515cc77cf9c7039e3aba4538a1cba27ccf752ed3b86443e464a37325a2b1fece9d727bdebce1f2beb45693a7d9122ed0c2d0c5ad704c31bfc54cd3a09cdb89e570c8721bb4dc3b81cdf8ac20fde6e298d493b55e54c8b713deb6ae8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83c5e01b7ea8e85981e4532da17b0fe7f38121057d8d7b464edf766f77ce8c63a79884f9ca3904ffca13e500be357629c2ac724620e62e16b08b8ac83d6a758a51c72af06a2373f342366bd8ec8eb8bed8bc665d29bfc8f3032b7269566f34d682b049bcf5ded1a98da0bfaa44c5a79d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc63bc645db250e096ff87bae1b79f956fde6ee67e05132b188946e839877a863fbd40cca2d131670a848fa351f2b5db91b9b4d172b8d93aa38bfb38c14faa4ee7a77229a3249ea41a8b7a5f7d5168773f32f5a4277e709e9b3d96f0c39595844f67d18630c5b604bbf783641f852f8f50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8f30d7f40ec8aadfe4c3872a40bee43b053f04baeb239838a7b1a7632bdaedeed36822254c89bee9f86ac426ff8ec667bd6364ec2d565c55657aa7488e79513efa3f48885eaac790f93f4569337692235c4afb203a2f10317d83bcfba40f3f16732e410bbda54d135d25d937f95f8b33;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59e38ccdcf311984f9d7c86f7640d6823f89b89cd681e745dec547c23a2f0d68d584ff64d11d20c479c55721b2a99b504d3bab0917b07ac649c029e820aab77dccbd8f8b0b87ee7e04827debf631868f9627f349dbe119bfb5bb521f882798bbd9058da8f07cb0a5f7ab25abd1e4128e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a4e6171954f1ffdbb498c16585bddb97a04ac60e11e2b13195f56683b7adec1e8993d2dc28c8ddf2c416b892d42dab5e75bdc7abbb21c3deaa977d540d3eaecfc945df2061866b336293412a439003129e0c88e5dea259cb8421e672d2c3c717a103699fa7d6681fcf4089d799f01bf1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6229901929a2ccf97ca2896f01efbfeeda0296d89d37988dbb73909509c0d3fde448174ef831e7b7a482eb109246e65233600e3c0f2a8383fdc23650aae88b8b9a5c281a9c2813a1ccbc42f1c3bf210f437c17abd3c547d2ef8c8278137f9814dd379badaff0bb3dcabf48fd10424de1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b7a190340bf49e01c54e883035d47d9162d5e975113588cdb2952ba446f63d7eb17ae7f7b22530c78625a47e9cd1a9a520647675fac703a4313331343ca036b9dd70d0f989222e24a759ec33c3c6bae8f9b8f2817d1e1356c606a56617875ac1de0c8c8700fa07a327f23b5cebaed673;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb266dcb1d2bb0d47b69ed31f73f444fee7ca32d35e1a6be768d427e78d48e452c419b49307309095724389fceea8b6d6d3fe4a90055a39f755a0dcec62565e5c102faa350ba12f55fe41ae5bfd8b453a6b6efa753a0885fe09138c9805fbcfbdfd29aad6972a9217625d8ca4fb8471a91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a80ccd9d6a47083199931be621a573c4293b910952f1064efab966bc098159009d79d0d9ffd9b031aaaaa0c49473760e274e90f9e66589230067bc6f2e641485b9a0710f8af74cb6fa60215676180c4ff379bf486f08778bb0dce3df69582c266eaf6ffeca3b583d138cf816293a8275;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h384d4ae2d8d97a84370e8b4a0a501ec959adbc9e63795f8334826e5092a7c0e7ff4f09797df5da19ca7f7a28089aabf69de3ab290113f7fa46c4c2f30d9c196249b85066c12aa154be6e718f9afa6aed054b40def369f14d9864655c2f2ec76d77aad13adaf7d2458edbd7a7246f450db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e107c22a2bf971369d2ba774f4293981768ed71df49432a3c86344bfeb534020316a903b33424e89898460f36a832b7e50ab8d21e9c3d837dcb8a2fd0a93dea88016766a34ef80d167bc630f040be85b44e1e7fb09de7d16eb171c2785e541090b238f47b59de9e57999350055cd3bac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9450a6f9b23670fe6d97b821e825df1b28a72d433888a4deeb33321239e09b96a109eb47179e1cdf6c045a0c2d7a8e79d8c1bd258042dc4a1cad30b92b3e8865b51ff77c0b28c347dbcbc69b2f6988f3622d533c4691a6b506ec0278a5746d3094952302f31c2e7909af2e01abcd5f84;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72479b81ba86b224677ad5fd180f725e680595fe0dc3c22ed8c898d837387af9d7e0ef9c36049070702eb110960281350b5660dd5a3fe3213052e2cde18677cf5cbbf38d9a1e4de3d521ca986712abaff97100742d932898612f518f97d348c620a6f43bfec12847967f60b74b363375b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1ef41a61c0c3ea25e11f41bf3684d454600a26cb1c9a30ce7826e884178684edd2ef821a6d690ee98132437bf47ca60666a1bd165d50861d03757a48e7847b98f7b686fbc07ab22791c56f6b8bd1394fea43a28504b11af18e25271e63b51831f003def4b425e5ca117eca632834eb98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h868af6cccb33dad2f737d8393087b5e62470e394cbdf055030901e73fc68c9d56b71ca680508c4d4a6ca4f9f6e8702da946e128bfdc424f600e9f0774225b536689cd2f1f9933d30cc526f26131d3dd4978d3650aef9db2cf0df9da1449924e36f43bb998ef72911f82516084eb1dcf40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87b8e6b7e70b2322cf710e4c6fb69d87b3ac79fa798c5d790cc131070965edd6abcda944dc7a8e34aafcefbc6fef2c100959cf6a00a632494932fa320be861671df5a4b32783482ade98291e4c53d796798c8ff0d189080c3a4b7e5bbd380c5462cf180a36f97ce64a3717a04314c23b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c6e6f54ddd59bc9269e4d965e1025cb4e2a27a7db03d50e3f8a3c14ba4660b6cc5366178b3d9eb31dcc0a19b4eb6fdf59bfcd9456c7f02d5fed71f421196eb233b53f0add51569b2b6d22c3b608e60264fd4a3e89bd0ecb315cca4d6f7b8d2dde4c5a8aa8803cd4eebfa6104cfa8e9da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c0a5cffedd825bd47ae1a4077fb955648e170e377739d2537ee23f9149f21d907f87ef62e752247d7f1fc6ecb991b6e25e43b98273ef707d25139b1f8f086c18656e446b9fa9ce4b2cc09bb2ccf090386b2b779267e94d35b255999a447b2b671625252e3f8bbd42c67ba8fd56f5a894;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haada64d32b0ec1391313455ce7d54e251fa294287182ba993f580842727fe3da54bbfaf1910f9f1f9a43f2429eb19b1bd3d35b841a2d3760dc287e692e6333ab2742d028c511d1ebad827b976d354bfa4e5a4518e8dc0aea00209e49bc12a18b0805310830a1fe2eccc718c655ff5478d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd10fe3c26a52909e431717fa8001d8f0b97c8c567b4cf69620b88f1969db788f15d5cbbfba1654aa4730d39dd192e9db8a2679f7588de8e6f43969df9e8c0857645b77f661bb0bceff9dc53d9d13d80d047a4708f59d29f44e0caf0ff69eeaac20eca987068997479cb468c78064aaab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbead60b206ee2a3d3c09bed1cc5acc8b436cfc2dce5d99f0ecd51d29a4c4705710d1998b67a28c4d61c8fbbfd561e421a29631a597340a04ef9c7df9cc119c7a0695b7d4d0055f40ccbd1cec42f18f27708cc4d3d3901fbbb6811149e270812420b9ebd0c781136aa591799db10c8ef9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45310a6e684f8711b9b59874008e92df6528b7ebf01a63fa1fd6087292edb4d26790c5f2f830eacf2d686b150e40c4dc31f1d132aadd9474fdd1dd41983767b898d63dff9c8964d3de71996058844c9d3dfc5b0c9d0357b9ba0bc47afaee87fbef458d0c6774039423d94ee71340cd925;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5682b3c49884c5bedbf4f24cbba92ca89480be953f4a8b95c1757f4c1dfbc3675469b0a8b94565461fcd80ddc0d50e27f532a1a29ccb42a4b854947c8a828839c06bb1600d8af4bfce925d6ca0c371cfcd897f81dc5b80acdcc2dbeeefbd3c5f7c4e41da937e7bfd56c9d62037dc4c81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5384e90238898ffc1638aa6bf3305af3026fe44517782a5e426015ab578461a77879843ee40181cfb41e0a38ccaf1bb2f43d2e8340919c21ac71fb4a951a45afb12b25e2f3c13f7fe3ef5719eacfbfdaa0f1c0de00b7574444cf7c2cc477c2bf755c81d0b42551018524f1e2e457bd5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d12386542df9e972d7839bc9a3e2c40a009a39a53e079b5921abb8f5b6b5356d786e3a8523ae6dc6594685ceb089af1f6580263512d26196a95ec47b04a14e55bc055d31c772ca7b86366a338dc7e974038fc64fae62ad4c8f7bbca5be999f7bf57ecdc2880fe303841d86fe4fc7db70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e6edf1db056a5ac92f2c17ef49fdf9a9b27429bc2c5c3ceb924684abb32ad481606783e09103a1bd15f90834cb13cf141370330de1d3c21b54f9c06ace5c19c17f5576168e34f79c6213904e032539fa001cedee7be9985d67fc6761ff719646e00bc090190e086927aabaf9f42e781d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4840326b29bd8321643b5127d0857e00c29fae5fadb91e9ddce10040dc9fdac7d2f3dca462f9e54488b7526951126e1d8916f7d2e28a4e1a858a69ca7a86b0f87dec4641a71a71e211461d3b0faa7440ea8aa55054b19c98a4654783bff6f6570b78720ea3d8e272f34d9295f7a7eda4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16becd731fdab96961a1f215916e6c1e914f957b66493fdab325aa461c50966b2f9e28690d6fa4220b3074e7d4038fdb5124f288aa8710f2f8b21a40da76c716a03ebea2a8250ca509ba284b4ba68a68e5eff128fb3afe9f92d7169edf7eba62cb5843c1132b3a114dfd6e78be7506ce8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h965c47f30144dc7451b29b497238d542f9564c0a572ba6a70ba791bf275629bd63fd801c05c335a628c3cc211e213f87ac7093c92484cca243070c4ff6454d5f4561f9b4bd5fb28dfab24f80dcd593d32063cc1a25d2870260651a4c5ac618fd2891582d7775736155bc45048bd5d830d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h423a5b7d9d4ad82f950e7adeab53f8c7e3452784aa57cd71a9ed2fc366dd4ff8439be975f4af28727b56ef5067103b29b522e9de2a349d5b484311743a9937cbd6e49f762ae3679bb46019da815bb5a4b450a4a9ce2d169001d44f7cb6ce0ce47061e172dc9e84c7dc43caddf2d57095b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68baef5b87887879512ef05a9dc9f13b769395dc0f9ef9125122e9bc92d9f24e4be920f8d002022d2d6bef8332fcec80205319db8741b8dc9d5069bfb9e5b9630f74acd754dc9a85f8b3ac0ddfc611935ffd24ec540898b0c5fd9bc2ff32c35de7b538f2dd1ddf1ed9e65f92cd78dd844;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fe96565dd08b988f4cbf859b839dba46f9b8222a43250e5b8b55a03f8a6009a7fdb8efd35bcaacb13dea08776125195d5f24c6d3849b7fb34476641586707fb09f2842c3b8d57ae50a384c71f5a5fb223bbeb7638992971cf22936b9c82a668a17ebe426b4ee8a454fd8a3cca806b9e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc81e9f04c32e451fe7583ccebec7f17d0ef403ff1c913a2551d8ddc21442553b124de0b0a90ef349d1c85e43492106f4c862bd772958d3ac38a799f43d5d8f5c48681446b40e3feb3e2c66cebf717c841e9209187533068d173896c71fd36a4d9153c00142d5edcbe1cc3c447fbd21671;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fbbf2174ab52ce8784331e2f37488471c7e6ac0ecde617a84b5cb1be3845f594af42c30300172dd99a0f59bd793ea3c999b3a8923a16f40d545c3ebeab6358f02c75ed97204fef5d5c6d68b1ab0405ccaf4876435bb4477abee15016560865c9d42e4aac4c797aa2f07a577a973b88d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1bbff8b440abf2c24b1171c9e077954ae9e36162e85271bb19e739118af872591215fd9cab507c9899b7335d8b8b4141e5fef5ab5fd8107e86e9e3671fdca931cb540a05118f47b783dca0cfdb92aa662677bc143776e150e03da2c4561648b7c151bc8a0e14d4d90e3460932e7ff91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73d3511f78e2e62b1c6dc2d3785a7b9aab05372ef57cf57ddc1d46a4bb3b585bae8fb812821c184f49af8ffefeb17400064311189031104bce7840d483af4f95cd89503e7d3031cccd0af2a53ca800d922ff51448d90acda23bfb82c9ac403821ac0068cd2a1773c90ca9c943f015e340;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf2f356e975b23451dd557cc8a551f5166076f4f825c98ae23378a88fe0f52c5dc5f3ce7d73da94ca3a20aa2a1c028fbbae360f4c7560da708aad59ccc1237ad683d0a58f78c828744b4a0a9d32feb518a54e75999ea152768c3546d98213f0ec4d9909d5411750492da19a52060a01a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0ee5ba90d5b19933c3e9333899909a10d5b110fabfde3b8c45c486d937da6d62095cd9c66208a34dd36b548adbc3ef90cb81f13e17f428292486fec0973f7551ec1f2460b802d03dd85f37170c227e79b2c4601dfda052ff6b020e8f399333b48807d043d8928615ab6b15e0df6d6f01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a6b39cca8c0670ad398d84601a82008bbeda9764d408adc5c1a2f73d4b463338c5ac3d6c47c5372464b0389a2438ecf55140ba26739c642800462148980a709ee55839107edd7be6184b6b28f1b4d92bb1111d8c0c39d3367b14cd5dcea704e0769cb1b4c971d5e8842b4b5b638681e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb4f47a78c7447059585591a5712da4121970f7744c3679cfcf49772db7cffac5dd481d9b30b3995cf3fee36d2212b88b06ef23964a4de2caa353d118716db57c300773c640525dbd06118f8589a94a64d4848670fea24ce24fba3b2966aef3a8f36ddc5da838de9faf1ccc53d5c33214;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4015c8886b5afabd49347b24084b3a9f3a6811b1675892c5698a0facce2e36669a74d4f540466995d9e3102208f056c5b76ca1cf5b8ecddd2e63a3cb16d08970462b8c50ed9336349245c380901aeec2d7572cdfd3911869798d4ead8737ba664b1d01b97a105dec65ed203668a5960b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70f0330f2fe2d2c477cf04c0b1ba1281fd491885473c2987e2f6ed2b788c68a0a86f7ff4c72a046d42c0bd24b6a0fbe3d8893d417b342bf29345249815b1c6e6b7b58b3220b4dd9464fc84b6ac995c04af8235fb3c8c86ac6b9a0a44ebb880162e53f0e7757bf9063db4f3a9adfea38c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88c4ae5e2fa18d9990ff38d8c8f2721cdc784de9166d4ac1f424934bb13d15d04594ae4f1e77f53adfa9ae1146a04033cdf2c1c92e9212e13f4ca5fce04dca7a561369b1cb82362e3abda3c38f344da84ed43264b09907f540e2ec04ca47fef9c33f3bb95ba847f5e039118b78c817dcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dbe6c92798f3753a0002a5695c117f43844eb08e3af3185f1c071da1c8cace15f1af125c35e1dd2bd0c024843d26e30461aabcee6c85bf0b4871d11a2e12ed04c347d6b5b1a71e08c2b46025f96eb22092905b65fc5aab0dad0c7cf766a89989113eb6465ecb8e0449c475f6b6fa8656;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5077b9a028d3b375e3e4516f1befa14d619ca22bc97198fe030ecc37eebb4ad0c8da6a7b608b8657065a0752d05e00b16986d4588b2ee0d084940bfa86e8828c8d2e8ffcd644e73b974377b20a31d5f73a1f7f548ac44e6902aff3241a2cfef627b112bd77425191bb152c26f3e7cd4ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d0c808f5862c3cad25a1f31ef022956693fa0205bf243f7c440fa9ee102822e7391aaff34691b7868ed2d4ff25dc4579436f73e04ea82b23c1676304b6312e509178b0b2055713472ae44855c8db4ed8553cd3fecfbe6ca9e54dfbf60b76ada919d2ea4526e42bffd9f9dadf7f7d1687;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaf8c8be55156321ff3c69bb59823826bb79838a4b39e870b0207c63282172960c21a2310bcdd9bdc8fa7647356eddfba5e5869227308f62adf07ced41abf6669f1346d9eabf156305bf841826ad789d6003c0ee844edb43d987be6b159cd5b3799d08e1364560e21ca448440e7aceba0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57adcbeaa8c364c422c6953b5ad6fc0fc445113829cd044a5d75821d33f390acd9070c9849d3391b347d6771cfd275dffae08d74f831f6e2dc28f046b4bb49c257eff6a42c38f11724a49e5ef477b850071a0433791eef47f2028db215bf31f2836e9f44f2a1d295c4317791b287a6d10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0db0dc9906fd3cd3708ebf1b32733fc248e4fd1032ecd59fb9e5e076957d9a7d3e3dda4970b5d20b40e253bf2886647542cf544f83e9e98127d9da5d21c1311653a6675905f082616f3cc4ddabe8e8305c7881bcdf609ac733ab213983f30c58085f3cbd182074a5cc1c6352ac4c11cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd75dfcd3f2bd8d3c2066ecf9b33a7e066ec90e84916b5ef2e916821b6a1507404bce564bb80fe10cdac7455c111254c7b6b2bf1824ab286d8f5b53e552d8724b885f21afbc9d94be74c0111ded9c99f288b2ab88f970c86894842a998e28627ae9d82e088ec25286178be522677163adc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a57f3676dce103bae8dd298924b3b64a5eb9d1bdf0d0603d37cde87469288919be8b5626ba475dab99d3e702de07f164503cf16157e5bbb7b0266ccdf9624a20bde1f6e919d3808e3aaec8be2343e62dbfe9a4ccf1936b2bbcc3a0df0e6966b5928b0b2f218666c23ef67ec6dc8abf3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he707d1c064406e01a349f54c6d13fd21d2607db1d04aa02938ce878be055754171086bf439bed93088f3e651da7ad3443700688ea4a7243a19194661c83073773def733236ce07fcdd501db4e28a592aec87e8743f0673ab8073ec62b69b82ad8364fc3d20a8222d820096e4919cfb7bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eb11bb8de078eb26be228ba952e9ac62a13a18c082e47364d87929be33d53c4d54e3782c7cb132da77fe90d7e2d4342ef35d0ebc6b97710d12ea694cdcc10feaa38c4940d9384f5e2dcd2d102fca7a23c2dee7530d966f6adcdbc69ae2569ddf73cf69e31e42950314fc707863ba760a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97e54d37c3a85695aa83884e89ff5b5a9ca8dd6aa4e38e770c3b6482dca1a26f389e2bf392c751311724121c18af8cc9b1c02db629a8b165951ec5303f0b1c50d227c1789e2e9da116646096f954731a45e7fef6e2a02d9cb9f2ca0fabbe961834c2e7f1a653f1a2c7f93dc891f311f73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2ca25581c5b7ec22d4bcd8bd4a53c60365e0aba493236fc1986ee0492fc2e9b783c1ff2c9b03b048422e13ba8a7a925742f4aeedb743c343e2940da29af9cf5913667b6daf2361ba5c1bff95020905259f14cddefaa7dec62fa3637b2d1009e72383b33f6d737f34e25940097990aa5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8644d37fb44a4a580850e7f8875bf576e8fb9ee8b0f6dee82c09f49d71fd90ff4877197b6348f6ce7ad4c647d3708a54894d5cdc39b74ce818088ec3d78b70602382a7ddc52591b4db08106ce12505096787853124ca264c557b2476efa3302872b6e9d6329d8e53b192a8e09a9456c6b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4de699dcce4ee035e870826932e0aac02be2951f32490f180ccda4bbd2af4bcafb20ac2c3063bc65ebe1124171b6c160ab8ff1351d0978911d2b7cc12d95929177923d06ad20401ef139e8900fa19956ec096a484446b0df3df1e91323095c177a315ae22223988e3f5f4e1013e56516;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36b79e763fd2dc67453b5b24fab6e5585dc555a57215072973ca2981ddb4662ec57bd66a12c54feeb40e959ccbd06afdd0c3869d3f906769cc4ca8cfd644bf99de2c5ba22507df2c402602ec4ddf6796c60b9292e2b46a8d9d5ea5fdab1db5dba1acb114ca50df9c5d12544f1530ec52f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0664025db08302db1c5a8e64fbbd4b9cee4d46f757b4b4090142cf63ad1f0626ec9510df43c7ef7a4470312e5c46e3ab16aabdd452f5b51b4d3a599140cb125168afaee8fc816682137fde7dac9c2ace9eae787ad88313ea387b0b0b6c84e05a9492b28201c4cea2119a23198a8f88a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f7f7b5a9f5a27d355a922f964b8a12e57d1f8d6928de95aea64e56c02286102096cc536c894c18942a695f79bfaec5c88168b239d6580f50bbe4ef5c2e930e3c4a0fc2985d5b0b23ef133c1a4a83814380a438d4dc379299b1932ec2dc18d9e5954add3ed1041b7c4f2c08b039da439c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76743165ff003a2581f1c9b80f95c51311f2c5e627c270bfcc756ed2150bd932cd35d6c758a0f8716359e9f1782b38df783e5858015908111dc66991428dbeb5d17d4c180c0d873a6f8e326774d165af209c51d911eb6c07a67f0f8c4e66a75f6558990160c92f74f860ab627a4873577;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5612c68a9b216483eb8926e827fe2909141415c126336975b6631f29b6bbae92a1cf6cbcd880ff77f9a6d0d2f3f56349b290b7e366b2a1ba61e75b94e30e440fc70521888dc5eb93f583b1381e423270dc4a4c04fadfb99a7a46ddf3893b7176e63ff1242e0b230a4543c2d8b80cd8913;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ca4c68a9de36efbb7888655e955d77df5f212f4877f3606c310b891ffe539813db42a103cec530b4ba8e9add26b04f2db49b7f5f3c35dec6fcc4896793b98aeb497355769ad351f5ab6d7b60f1054b131b0ec3de45cb806fa4a958e04ea073de0d487699ceaeb7e1130d51a8ea28cf54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha68a2dab7fa1ca2335d06fe5629cc2e94d8884f8581f99cfa0395dd1419a9a452292699517e5cf7f6a5e41e887092f389cdade386e58c767133edfb1c4cb01e736c9dce07972ffab5b862ad703ccc805339542cfe4922dd7d21376bc787f0eb566d173e556324983f7ad046ae81c35588;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1aae4c94fe5ada81c4659eca7f2d8c8272812049134e8a3b30d7b5d370d77ca9f811af8b0e3ce40c723a244735577e949f567149759b8b6bab5886fb8ae5f511833fa68d8000950d3263e860fecf13f53f4b4d1068500a093808a00c9157c37fda8a4736f930b9b78643ea119be9bb7b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e449c9f241b41dd93355bf1342b361c2494796256274288bee1fdb33307159edfc57940665c9f15dce700687ff1e297b39c2bfc622220b0fc1a5d8299a6ec06782c7f60cd2de9853d98f78858445e714d706a818e3bdbc2cb28115cbdacb1a702d0117149a5442f7d87f6061fedbf6a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ffd072b5007ac665af8c1b89385de832b9ce39cf8b79b24099afbcd1db96518e9b03e97c6f21697447cc8c43a28b5bcd1f5d49fafab2e1956e4be480a0a91df86a7f1a9af94e01395843fab667962d82f25a4704837c73f060410a163b9f14a06e4be0c7b310e3d76c1d9550c82a6fac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha96e5ced35752d127674ee659fbaa6e53f1f8cce7d80b831e8ab2b7e93b5041372025c890b81a282beda2ebdde6a04716e9a523a39ceb4ae02819e4809f8630a3a1ad7249053d71533b7d2bf0d772e95c11034154131b0e9ec7ae4ab82d5e07520548fffd3764515435311cd735078e39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fc8f25aaaa8330cda0590922ffd174ca9dafae3dd9450906a433d23e9eeeac1abe62d7f76f4bdcb070da876ecfcd3dad9ecef16a434ff91fead44e4a7f13a59fc36b944df3db6987951f930a2531273dc1efabfc1b39acf60c99e9b99d42b62757b6745692f68a24f16e8a8ed5dffda8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had33c7634df41cc9942f496e733c28c4a36dc993bb47dee37b90990854c7d889bec44b218c809e3ff661a6c08c2c9699890d05fd4fd1b3022f2384eca09a5867f25210d30bf72d3ce74a67571d3bc04fd15ec0ae2b470521ac847297e4e26a032c6df3457ad2cd6e6ba09a74d79600487;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26daae133d99aed5a934684454d6e766952e9e8e335104fca686fb7b71f16c31d2010c4fc9034186fdc1d7716c3bda0cf5c3ddd9a91291e458d9fbf2f74b36e0ae2ca7cd5661a61d555e0d9dd144e62c9e7e0ee810ebdd434125a47e6f3e5fa1efefb6dca60fc2cd491647661e834ce9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0b09d74f213f73cd660f9c0e174127484e89d72b15e6405bea225c2ac84c5aa9568b0846d307e1c91ebac2255303e3ea7d6b28e658ad639aa39e8f03940c0b4384107774dd50a7b78df6d174f71ae53bfb905d5c96b21da4291bd6756550cd3a89e1775a96b0ccbcb342aad23734c2de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he96b0948a4abf5b87694286890553a0b7a96bffa810199aa6a7377904e7a4b349835681491b5b15488bd99547fa357e29cf93daaf032d7eb28bbb7f266b68efe637b277cc65f1dcb2fadf7bfe961b20e90567e2c06f0abd71a2611fd93b9281b8b344792204fa52519c13a2d3bc2c2ef2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81f49d822e3ae0018c3b0773d9644f52b3ab535b87fdf6a9d61b35e9748132aa897890dc8660adf8e0359a62d23612c1c0b3fabb062d804996f6963f59a230cefa6b3f5e2ccd470892e03557a50a38696817cc5b79270c4d8fe2b358f94f79e9bb530b2c721f050f803fe80e9aa9a26ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbffcc3e0992397f1cdaadff8ed95610fe9124aeea106a3f9cb61ecc28b4861654f7e257bc86e01b5d55b6f37a1aea987142effd760fa6b6d508333500f3b3ffd7774211039758aa094ff80b9ceba3c3053cfeacd7bebc1da1562ec5b5a495012eaa154a20c21caff2fc10af6988d6421;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38cdb93f6fdb97a9216d54c695538450aca44875626b6e5140c62d9622912947bae9c78cc04ef4cb6462d5abd5dea8df9fa509852d4002099677e0f113150bfdd4cf94471172d01c8a1e6492ee40bfa9bec1b282ae69abbedcec3b9aa71f525bdeb3e9d57c2876a0017d7d89eb9819bf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1879c8de505f0b450ebcbbf19cdd23c40b2b21fce07c2d6f1e270e32c2163ddf84cd592d21e4d99b7853e3f6c5d8ce7f9647e67548de04e91f7acc89c60d28c3744bcaa862fb027fb62b70ddfd795ebb5ea8592ccdb9c7bb5ec07c1ae7753cbde1cf0d1e18b4245f6c12e2d0182fce5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e7741b5448f5323d5965311e70d37abb69e42869ad45e16ccd6a8404f739b29955ad33ff65a4457c4ce980903872c00c75725d6b65cec26b191e6066fac2daa6107047e40ba780a20223fc7d133c1f6bacc40af0cfbf0738702fcba2f60405e8e5610167a23a0c8981d23b7c544d8915;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h357617f5abb341fbf56804dedcd06d1d513cc6ebf3779177b617f25e6ae5d8752b1632bf83806c248cf13e5dfa18ff530b5319c108c8852d5d7dc101eb177b64cb543c7662ad5580ab072be78131a29c5ddd3c3853569398425e6ae75eab5fb2b8ea224a80dab8319ee4617a6675ec58f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha71a70e0cc6587d29657b43da30458e8bb794f083370ce5605f68fcf0dcabb2e00798548d9e43b155882c72e509abf353a077bdae05211d2bc93dcac030674ff1a5a1efe08bae772b8c6edfd8ea8bfc1ac0c54f12f799d5ced501a1a3ef6eb86d6381f8b1e0aff290f8401b0ecdc17204;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc842909db2b244b2f628cda9e7f92186d4bf007a87a0667669d5358b9acadd8b5cb60b7efcd835ce58341eb56c6cbbdf849d794295f234f815874cc22ee8aee5ada6e5f8e8ca4a0e5f25fe67765c3147c697f6b61e04e54c02535288e38b43c22ff30aa777dfddec94c91be75d42f1468;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6be2ec17706397ea87dc974a2ccce123bf0fdab235add437eaa4bd24ab120d073c9cc7fe93180dd5df88b5dc596a60314a9eaeb2d36e2e81a5c397d848e76ea238a52737b7a35dcc20155164026835eed8705968f196355b957d3cee001d425b1411e134c97c8dc1bc55a37a003958d3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcca005c20355195d190a06b86dbc7267e33340afe34fa84cf4cc9bf3124402202445f525e59b01107ee6a8dba0f9fe7b5f29428916695ce9effeae765a4e917a53590688441889a5959a7e96dc469fe7e796265c0c5079c126d75e627542d0df27437f9b6d88872f932802aa87f8f342f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0e9291e1dd3e42f9b557345228ce9909a56ed514de06ce3aee4a81847c8e4349d3457a98cb35411728f7ecc747991f4c628b7a1026f48a87d07418f851fd7af8cfb6640f357d03ee8452805ed11639291a3feb93405c57b9b402d8908d701361d3d1a71e1adbc02d5c50986a0965b0ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfad13a5e38960309082ce34823c834eaa67f1f4d3edf671db4a4ab7917eafe0e4b0d3b08be1e618124528ce1bccea026cbf04c58430a8056b286d187b6cf1f09ad69ab05874b02e94d4b528070ca34d8771eefab7461be05a526f3faf09f56194de03af3d39a07497f25fec5ce6330e39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haac61f6f7b5de36497d8ef9cc082c1cb43f7bcf269c86585c56c4455e44c083ec452f1262adf98346715b0f9444f6117a0b1259e762fab8010ca6aedcb83ae549976096fafff394c5aa59b4c9f29112aac5d6eb89606d96b561cc946628d4727bdbd1a690beaa6e367ac20280d9d3ecbd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b35f88f2164aedbac1b53c8badc04c62ebe786493f3dd0a5b28f5971ce57ec2e7048995828cafc3408988da3930f0410dba55a1056136e7a10458bb7dfba451a38fc115fd1c5af0a281cb2dd3448f1e151683ab49771cc17dbfd99e0ee6b1841ccd38836547ae08199c7298b44f84e4f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdf1c6b95d4904166a0c9a86aa345901187fd8ad699a22a8755417f4a4ae7fa87860bf0050838877da36fc3e61d11c735fd7600051f41e5184ee1b086225ff806943114aeb9784dc2bbf3bd1acaaf12fe874128330cb5d970793a212320bebef7a4dd84558115412910860a10cb1d66c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d7a79cd1579fca150c16616c4d86f18c997c9cda5674f515355ff8b4287cd5a6cf6fc5ce2861b9e6e7a920a778aabd0b964ac8e6262e511b9a5057e87d516c46384230031dee295822510ea1499c92c08ab46d95e5de3d4e6ce68d4c724a8dfbd6786709a38fd10a92c9616af1e6210;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c2c7bbfd34bec9665cb7a1e121b9ab1f7a1e68be3ea6480faabd33ca61d82471a05e8e414338e514a0b6d9b26343288b6ef876d4e30ab05959afb294745eca98c31b75c856f9acfe7dfdd80e9bc74345d528e31abcaf476f291013162725f495d044115584f25a953beae35c1fb08622;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc86e3015f62a7d9cca8c5bbfbf60b277014f36d6c6a54b006cbbdc9ffa042d70f21f39e6d73ce92ca21416fe8e8779a906d2a98d63e7b6a48ac2accc7f15875846362bf83623f27591e6dc95c0cede4afe7c70f64739ad5382198eb651484bcd045e9e211fb4c6e91874edcd24b4ff334;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12a89e864371d9ce3c5d362fe0012cc2ca1c6d05e7d4b3541167a42adfd0810f5b38053ef6d71e47f7e7350f323f74b579b84204d3e12a42f4784171341517951c55872a3a0adef52c98b55bf097383c7f3177b444cda1c9fc04f4537542e580346514d964b2333a6667b2acb59db5036;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f0dda25f009fe0ac7cd1ae8ed58a86658da2cd64522a8e2036d201c74a23de7c42f5281135920c84664805a8069937199efdc365219fffb7316dc8d0c3d7ec00b3ee16f3249812e6e803840ddacf9747e0babf659996fb32775aba3217e81ac2617cf79ec6df244ee7da1b10a6177b85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96bf8e6a789c9c4b3b7ea56c393df4e087e53ed80ff503e67ba818c2e48f8eea5a9ab429ae7b37a8bbe16d9568c9b088773973add953682c92ed76adace94dd6afae8c3e300cb230ff697e9f0fffe619081a5ef5e809246a23f97e7acb15a3ac3a2d0e33cc22260816e949548975f3b9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8c23ffe359cc2e6811c629162aa00f85c30f08e94f0f31d4a6bb5d4870a1d574f264c62a793a1e13441d987f13ed4d4cdc4d1640b2cf8b2819cc4f6e287bab08019453a80bb21f084a43d63c2debc8021bf02a9df6f34a64d16523b6ed48cca1b36f905e7874d9bc525a66c8933b2e6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50252824a760664c9e663926d32ce46356db40456233334243423301fa6e083c9e70cb72629268a65994a48acbfb2a981077ec922b1bb2e3d03fd961129263198a05b9cfe04c3c616efbd4bc6a85d69b85d37d77fe2e02f3b0e03f2c81b174eb7623659cf6b81aa506414c18c3158d84e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ef2af29e91db5188d38effd82f8bd3afa59e24c3b7b6def77d436d36fc83e8c1aaba983f65062ddc583224acdd9d099fecd3d467150852296de33701946dbd75d89d2721c47c94b949540a7e4af29fdfe3baa24e683a6180c12230717497b0e47f0218d84c4fef8335956507d10fa1bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42cccf53fd2237163ccd4f0225ae20e8846128560523c9e081178a39441817d720d3c39fc688089f4f2ae34fb630f681ec6d5b58964595412d73f535a20f062323e96da6c0f9cb7ad788912936b97db1703135ec10ebd7125f93bf572048023ff805ec6731821567a8636581be7f8478;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49d4d0a4c90b1d2f3c2722a41d9e90f3044e5b435b239be78c0f5159cab739fadc5728126748a234403baaa5209f1a95bca77d229c1994085681f8069f7284e4011b62ac917c548299ab51681faab4a7f8b041fc47db97cab86ab12e70f5d9b46829f1a300f0bc13fcf0e02b0fe15036;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60d7d70654c1d2be840068158096d845a5d4f1518190dd8e2b29256f7ef7fd919deb329586b05ef2218f54d707da70f41298a4a5cc3d2d1def7aef36817c4dc171a103e5f3986916b5b85c052375d7e87a26d670116e874f84cb12daa2bd69ca6ec60f0a93282c79edc83deedb099256d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed7ba560ad0d401a5e251c77036b033dfee9557f3f75077f5991d551f84c41d39fe93fe8145dcfcac0e9ba0c4a8d2b33a21330a999885a0e844b4deccdcdd2ae9e98df4f99a1038f83eb0d08602d08bbcae5e159b7ed1b98bdc92c04a711e4b0991ac3c37637609b39286ff94864b5848;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee61cb93ab3b9c2c30f92535c4e18aa138d9d3f164af433f0e581a865f782c66eaa4edf67a6dbb15970f8f72d86d00cdd6f1784852cf2eb668dfc9e9ab6e4f51b13acb5eae4b15fc90863191964a69bcf6267a485b031d1d951f893e6a03d876b9dd709fdee0b11c105ae089e674627ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1758a9c8c0d0cea0901570c2c4081c9e38456217c326bd14c25930423799ca48f933ac15419e9ed8dada1807672f603a6ac418fd1ec34bccee5728ea37f4540ae00c9b7ad93cd3220b2562832744274e4bdffc239338316fde294df0b7d15c245440fa59bda5bbb9df237dfe758600f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ecc5ba169bd27824ef83dcbc1463103905721a5fbdca16b9998d1048b4f606e7a7f8551ffee9f4bff9d014c02039e9927cd59b9b7eca83cc753e3c995c244350fd8404332780ca8de1f7e766ce78e960aa6ad32bc457a334a6d59c64730c425a96b7ac697319b1988b61136cdb9da78d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf200ed9287bf0bc7c77431940f9b3bb68eee553ad83d690713ca0bd9c72394a5d070c43a63dd8d67e46f01f907e94b8fbfda956d3089683f538f629337bbc63076531653e319a05de64b9a8cdfd1219ca042d6c0362691625d4c212a86055a1c3956b8b0df4a51232e296c5d0c23f2723;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12c6e867e27e9a2d411e5033a1cba6ae36d282e12ac975bf98e8661f2868fd5af05c70cde1cfdc0d5e09c61de4a9745498009da86ca9937c3ce6727d0c3d60cb280b98f49e8dfbc7746953fd34db7f5cfb986aaef5303ffd424326dfdedcb6c2075579b6734815c857ba1b00e6ddd7305;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e59155a9cdb985eab462c66d22485aceb689cbe5e340ca0e24c67deceb67fbdb7a22f5872e5947bba56647266ce9efd1c7fcc3de602df89d0e3ee03909dcbde72cea0fd2bd51cb0190edcdb69488d35d5a1c584f1280f406acef16b28a2321ca2c4120e3641f6a96b845fd23f158a1b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9202d950b4779876ffc8dfaa6680505fe9d2ebce0238190371588478a7bed0792c388a8eaa235e403426b29c458f91950d3e4e8137f1499cf372085394804f886da508c571516c6cb312658f781564ca2527586b1cc085f65afa483e15e47151fd8968240047b781a694f066502c8ec69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf81c93d31a15ec54b619a5174a3f7ce6577824da892abf29e6c70cfcc87dcbb57d604b826dfebab4a6d0eb09c799860b2371e605b29334b303e8aa41924d877a0642c59a03833263e99840a6ced422bacf10303c51797b80caf32d4c10ccecbfc18e9e1c6660d8446b876503d081c229f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91ecc5b13ee0f8879b12b334b9c304ffa086f5568b60591f864b5ab640204799524d2b4b1eab84c5db10965a88cc6340b3f719d4b82f7e7198c16b83a0d840a29a916265d7c7a218a36142f64a1ec487148e127e356a778411b70a1560293ae2645e72ba059d5a231bfde54cdf9af6fd3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae3fcfbeba5e84dcfc7685fbc58ec18a7c817919f8b3a8b9cbc6fe68a54e702c3e7c1ac6c059b825989bce8cd123a0a23b58554e049d058a32a2231718c0c59c0c89a2c956b17fbc6798d4e39ed727f0ffe9fe43b92f7a3844943a7d971a326f0af20445020f0ba82cc9692a508ea5c9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b47bd2df5776ef7d9e601e9ece6c34b78370f9b24c7a754345aedf154d134840432084109d7641ec349a3a760cb84e7c708091d42b4a65cad0c84f498d2d37fd8cba84c482dcf79fc406b0b730a74c4a210ac717a6d43704148c73290cd328251f7ce05515689e0e227e38259ab21034;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h880c519ffedaaf7abb233cd59301f3d47dc9071a89f9c02656fcd1757bc000a5ae9f5d5e4dc9798f85ec3fbece08153701914bb5f5fc1e932a84acb8e69ecb77ac23a622076b43b57804c8e19767f69c38c751fcace012e81fd9a9d4c5a250b900d1edf89eb79ac8c89eb92240e521ef4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8800559db448d2e7ab218eea6e605972ca37daaeb1a38f62e3bcaa39e29763f00668b035bc369ac786860f85c21f74b99857a7e7677db5fd1dfe070980eaf46b09986b9441cdd15fdef1d3e1d794d8384bb1c3bd938cc557e11a18d645636f22725c5eb06b44a63b302d6ce4114c37f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha48971c664024239b42178a91939dd5f43ae671052adabc02a7576a303fc4a7b26e0d60d850813a06ce2b92e41f096d5df961ab225cf95d3c8a783ba48ecc4a6ff75e8fe6eb63b17bdf45ddae66219a57b80b8cc54692f27336f67387a16a2e279cfe0897400f3aeb9ded871bd308738f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6debc006dade317dd39a69313e3bb8dc038c82f6276e5ba07fea3e541df8409b478431014dda91e3f1b4383d757976c18bfcf508670c8f259dd673991b66eee9704e77a0d02c20397864458411a92e2986dd3534fe7f5fc5bb4752368bd48382c71c658b97d07554a0e049ec574cc0f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h929095ad43a756f6202de95d21d9c1548847f40dd1e9d13a5f2be7748de5d307933ee0454f86ce93a63606e89833e470c4a333776464839f8e451fa43be4d37ab499786ecbb5e205707a0795efe6cc85cbc5ebe5cc7c1bf0df2b8bbfafbc9f79da2628fe0ad2d3a4241fe9d64cc260aac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68bf7dabea6e36ff8550adbdec41c04ce8b4b0086e0bce697d0de18db62ffc58b92929c534f23d729a5532b43158317e86d0c427d0cff6f299d18c40bf395f3aaea7d1b71c5250d7bc128234b1a16e2ad7701ef094cb89c17365e36075aad79acb4231bd2e5a07bb1b18c630e7630d888;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he860ce26c1c565990ab68a207c3559bd520b2b6f38d0b907626277f99f0e4590a915b131c1beb8dc067e092c1ad7a4bc3468593b6c63e23df6cc70602d295f03ae988e24b6dfd69ec7104028c8c6e6dc16c939752ef8092b21a333ca63bf125b661a26ec0ac565fb124f1ef376c1de7d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4f8aafd680bbe03e579da2090d1d9c3f4772c170a84507322179ce713194ddf71d3acf606c2282d5087a8bd418d65df9053d09541f0f83bce61f0d4321a67fe6a938ac0e7e33786d195415bd6e1e5ec98dd88ed6d80d4f389f956a57e62c92c7b2cbb891eb7d3f17fc63cf0a6d99a267;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h912318de9936c2fbd1c5c60de37dc70be6664fea1f08fd1c1b933f389c261dd4e7023d93fe9ab192c8891f1684e808a0cf637883fd154b66d6afaa69cc9879cb00797aedfbde856e63341d0329e0c569bf0a7906c8c0c3de07b299cde41089234c8577a518171432bbbb8f11308ac8424;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h128f19dac630550b7bbe4061853f19b28aa2a1bc44139a9c65e0bc2acef7a5dc33478ff8b2cb65f3e064fed40f3604028196b7b8f2ff86a0424a8fa5e484f368a60d4f8b136f6d2a9eb9eb768010c2847712ddebaee374c5286706ac4b31f992f61febcf45452d6caea1534b75f641609;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5337adcee080326976a987e78cf5d4c8c795a0aa7791cbe71cb293d3fe70e00e9b11d513879ca6f8a6b3420e531cb3ed6fbb3aa3aa01290109cda9da92a95e3b7ecabbee78835b3ffc5ed54684bfa0dab231abb815efbf49c8edfd9627aaa78c8c8025903d686a9f6c5cefb46ab01c4ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf74cbc011ff43146f8d8a025cea42a5d835604f42615e2e57578f6f71bb2c935d1061b7890190fd61029a8951d96c6b3fae13d32c9bfd54d3a6da6dd312179b7d18be2e78166813d9492e553c783a28cfd20bd9124142de086b170cafb0e2cdebeade0b1a2b14c00bb48d07a934457e65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e17f1e81529523358e82a76ed16e2a4fcaef5f1e8ac20f1e17bb6c844f70fa1bf076a3a3ae5e2a5f981f6042471a4d2f1a8eeb02c69a3736e81ea77474a7378a61b23548165877d961a680c2d0d71bd60937bb787900d530f62685d5df17ff8d0ec28be12a6b886fc9cbf24a0ade9ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c16ee444ea582e9f5903397e1d70e80c12016eb31239a6fccca7158ec28debe7bdcfd01af5fe7c3c530d15bb32e20ba8d1a7a204ae48c188954a91e1714434aa921e6e7ad0ace6c061d6fb44f4e35fae09d5a4e429a838a30a44ae22244578de12affe0d5a16437bcd4852e8f72a010f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c73b284963fbc374d42e149c4d2b16a09727a0b4593e516c08db3498b461b57713719669820f61b364002ee6bde35dd59f0019298bca269a97482e3b6dcdaab305f4721bb7a8846c0675e631dcd3ecb73c37046f9231b3d3c35678cfcad46bae0329bf16ab5a3bd3f4dd1328b5b70a85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24ff031205eb6d8b0519e912001e25f59dd99a3aa05b66d232e9fd5dc829d13c5e4c9ae4221c5ae4da1585b42567b5dde81dcbd01793d199a760b302f303387b58c0d8c453a7c1c0af8406e8f8556e2674abd4767c4192a778bd62dff70de6d5c376650182657828123cda55949628766;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb29f2d1e3882a4c4286fd2c080d2d1d3bdddc5c8202e6e5d1c4703db6b199232c50ad8d436015905c80a9d1a18312bf7ab4804d0dfd3b457a3d9e6553526b1c3431f4be4d32614492a3b7b3934d353526dc9bdf8db8316f6bc44abd857bdaccca2ff8a0ab2a4329e7afb09a17014d3a6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c0c8ee3a685b0145265fda49113b6ced412ee834688076cd5d45304d4bef7d8bdfbd62b881cd4ce38e3e70d169e55bea17b05debb085d59f81d7091b1ee0865c6896ef587812bab99fc1e67bed1082b1f55d56e4135859d97626ef0875132ac2d0882ea158b633ad8936aa989a1c841f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda540b2367d4e4d131dbe78328a732ffe64ea378f20e6cecff381ec99818da0924e7e7987381ca328fa90a4789f242d05655211025cd06c4b2c465da2dc008f989bdd79f982a528a4841886293fd1b3f83544a2bc04a28bedfa3fea2b388e330f523cf29a205bc3a8cc70dbd46608b7ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfc72bf038d646609278cf53743e939c3c124ae65acdee9e387b12170ed481376a642abfd1714244dc30cca9a7fcad913cbd144b3ce481a78c744d69fd464ad372aa914f504d833eff3ba5f25279c4b29714311541d00d7318d909cac3ccb41dd21d30877efced238423850e07854bda5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb60e424329a452c158751be6f699ca5cbfd6f08078c50b39ace434af16143fcaf82059b2c1394ece2b87dd334d1518b4f2c632a32f4b1c2c45873f8f3038d4148ae602c7b4dae2bf7c29fd8c0536b532e27e057133598f7deed23b2998d356ce941c6cc5547086451b4344b8971b99020;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fa2cb3e8d988a9730903494394618a82bf5e6901b4b3f969777a34dba4cf33ecf65852961e7b6a55cc6be989b9b0e4135aac4afc29fc3ead017659e382170f4f3ee48ba397f74a371878812589e7baa03dec63c90e1ed8d77ebd300b185895156eed22ca7fd888c134ce5709960a26ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h652d365bb7d4d7315bac7f9dcf4bdfeba2ba010f2de588878969766a85625b638e0c622d32c4428cafd5e5300d8197efd52e418ba518b78f0eab7892cc51ad1245b6e2fbc1157ffdfe17f0a6fc4558e1ded8af60401e821659d10ec5b7f781fe5a23e5c4b05a6b1e89bd48f9031d57b49;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a60d1033adf7a75acfa759104a5a555486fea0e54078b8deaf3c230a82adb63460f0fd09e3a333da4bcc56ae333af799788ba68012a4656fe2065dbb3ed536e898569bbb501c3a0bd03f2a1eebea85f82cad736da19d180650f553a631e81a20852695b33a847831fd64b7cf6024197c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ad508d7a030030970810adfb3e243c42f20e55e79cc5129c26a9ef0df65c42874813cfecc14324c7ad5d51cc6120721bc4c62a6117431d0c1ceb9aeba6979a71122d2c87bf6bfe5b65c8585cb9cd32d9fcef0d9d28f12842f789ad22c19525c1e7190482744effe4179493c557926a52;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h544471b6784b8e370cbb8198c1090b04a9c019271327fab129b869931472a034317a4ff07929fee8d6d159323ce2de7f83f1dea26dcbb1d8e21c4b137bf418a265d7380fde8c898b4452edb48695b877acecdf1085e66bdaf91ba68a2662d68b7ecee323dafbfeca10ac18cdba08c47b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4757de6dce2be378e48c98df50d2a10dc7158d45916d7a945a065b61d9b4ce4cbef0d82374434feff29a9aa1d1d3556a3dfdefb86ef6567367589e400b3bf15314315a608eb64504e6caa76dc4779592c0f28e68085dfb7758060bcaafe5ca95ab93e3e77307cf6db6e1e1d8df4bb250c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5b0768da13a6e8bd012efa44d1599a291f219edae7ec4cc82a619a244211aa7f6440f18f25f10fdf15b2af8996f68c3262ec6978db9b8bb02c3ef8b17a8c4ba2236b1485750654f5e7982253dd638663ae2281822b6c7db64854393c06b0792a7bc8c88b10b2792a18788d7a59d49505;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d805bde5369f9814400731cdca74fab1566b2bec0adcb53862e87afe1d8df96a03d4b1b0c8c4a3d95c72f87d346c8444bca656403ba2afb765651b07999b6e5f84e56b0c6f4df1fa8e67dd9227f59453e88d28afd1c7deebb751176fd5a045a9760da9dca9ac4ece254f9c6ca591f140;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea3a7fa3c7507817304d15245d92eacf4e3de220535bf826c104b7bf068abe55826e7c916075234df201da99434312712880d5ad3403f0f62b35ce2e13ca730af94ba6f3f6c1e189b6d64e777ce96367e2a5fe8faf3c27d934696edf33b1d13aa19714a2ebbbd7d55ebe732ae63cadb1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae8cd5376beabddf0a907784cbab02942ef1138ee72bab16b0ea1488c39b14069fb1b88ba998fd0212cc696fc4c758b82f905b6784ec9e65450ce2d69180b9aef7714a150b50c81a86ae82ba81739d2326fbf5babbb75ac46d9f19e0c024e3f1a94eb5bb73c46d82328d58f17e1cd9736;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb869b4656a59b5a10ab1341c977d225c505383fa6ddadb129849b6389cc4e0b7f9a969d4f80781bee1ccb47527e3165fb8b983c12f58c737ebf314f70f7567499769b2cae7700ef9a187b03983cfbd7d039662a7466257e62d50e092f5fc7470e04a857305e5b04b9caf69ddcaf4e89e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aa3cab44283a419b577c77c83c6f1a0a34d9c1edac52b993a5789b81507dd223d1286ed8334f3d760d49e94e123f664663e6ff4194c2fde878ebfe656a15152aef5cd980302d6377d7b9a9ce38545a2718301ea2e29819ff598a5c2f5f488cdbe08d1957a763bc2afc8e5a0d93c8f0f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha974c554d815f0e64240b7aa2b78841ed0078eaae35c5fbb0cb0a2ae210ae23694257173407f92e09989355cad3f227d8f8ff8881377398778d5310fc7da2bcd4c78f82b4484e5f6b103097ee528c3b12626c8a5d49a50e77e8840e657ade5825eafe0b669a5c8f5a7fc2c5942ee0b823;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eb163c1a46b1e5a3a34033be2dbe11560d28192211df37a16fc51d40b1c5bf1780931b27d0a8414c4d801a8edb4f04d3f078bdc0653903d5a789cd48ed7d85c91be5c28a50592345720078d425885af0c94fb46fac5af60e1358999c39e58bfe4dee98f6daddda665c544c29514f143e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3176bc9c3ebcd62ae6f2c9f1be539d3e665c2571c3f1d19827c08a18809bf78ed0a54ca91830968fb6ebef738ad465589e9fb2a030f480ac7bdc2e00a3453bd1ed35f227ae71c091ce55536fc7ac84140ac021a11ddedfb81ee5cfb86ec7866fef697c1a884b84b332dd693d8b40e3887;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2877aaa3b7997dd49221764ace7943a9ee55ca3e8143cb2f056c9e02ab7fcfa221d3a7b9eb9fa673d6e050dfc34da31dee896a196352c3cf0c31954ebe32809cdf22e4cfcf1960fa9e5af4c88afab956f3e17542091707d4e907da37fa6161027459b87916fa8411a1a0e44c376867956;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h256938dd3758a919e805d3d8a6c04c01eba07a69de3fe38b839805a6cd5b9069de70428debf3e15d2e7ff16b7de81cd9cc400cd4443113209c346351a8f8083dd5f4886a266080f28eee889a0ea9fb99318eb807ce2f6d460ec507644842d02e9f4ad7571ae2d873464123fae086f2e9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b4adc9eac7fb4ecdfef3425229c7b19824d5db689b7a245edfb764d12db97c4a624ee5012890c8b47621d1efd6ed1689f6fcbda23f3338361097119328d6e2163201a9c7a58bc31bb33f86d29d3249a46318ed2395aa7363059758e9f84fdc7e7c8b6e4bc5a13ad5ef1d32ded215bda9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82fc29562b6bef844eaf63e78355f3b438c6b9acddcb2fbe4e28525664d6bb05c4f8b483a40f6b3f1ccdbae40cab3cf4123451c568c01b30db3c2ddb8f450c392f2a90d88ac7a7f79a1c82e19ea9d5c377050fc1b28f9266c581f40b17e567dcec5140812bdbe79bb311f0cbc11e89a31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22f040bb686348f4d3900a6a97934a93567d951759f74ef8f95d9577847766d309a4aedd109d9c74dc2fa3947d58132a8ea61b21de1703727d29c32d78f9a14fcab0788a9fd11e93cf07a6b9b1087b7058d8a717ab929e7e5318bd81c6c196c5c0ae4ab605d61b3ec06f9f8b53539eb70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2a211d90c3310fe2f9908e52a44e4f0743a5ca853f52288bc517a95650b29a3c4833a16489565e0c285d6e167a6a9c1ec601073e41e733a756d26299cb0d0d209228331b389daf6c1ba78b1a138ec83d3fc97d24d5949dce2bd39a1cd2c04094b3a8447fa50bb0a24183353291ec8177;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d4cea8eb63381ece9031b51ecac2223afa45d6e877542d760f974f0b15fc9b87587dd036787e7a50ff802f5a175404450167a0bdb377c21a0b155d1784a841c1d89415ff760c995aa8af0c304dfef25cce786bffd9698e3825289ec63e0ef5dc9c42f5ed4d7f5592f1ebfe48584b43c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff8ff8a9c6dbf950a5ac710064294cd0fc0ed50d81fc9af1d36688d079412b5895b3205ce41ab2c8aaadacb947d2fd7ba5f2265fafc10fc7a8ce4046140954a35c16b549d55421d0934ffba59a13a401654373d8a466cd6e9a5605153ba4bb972e44bad232ee0d3d53c9fc4b25cbe6050;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b34f705bdebb3087b601804af40c598ed7f7cf3d36c82111612a8d782a5426ae335acf5947c127591abdaac64b1870731d2ff7586b0cb0b7615655dbf78a0f7fece99c1796aa9620f6ba7bd1027d5ce9d792f00419ee69e026cad8d4f19b2001b1daf304bc2f07d40572d12b7cfd4587;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8d6e3ca3009a155d5e12d8e1cdd15eabdc9d759f178fbe2e2f454920043baf483da98a3ebbeda418ef8905e5c490d7b99d1fdd7dea5138b97f19dd1c0d50c424e994ef15e444dec15e328ec475349eac8a5a6787d978918337793bd5bf8293e645be1bc1570fea4e2b61a9f54b3956c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef23c087888e0cc48b59d663d5b12b98f420ec3b554828315cf456014dee4b5c4ff3d2db9e751b50bb1a1b773923bef7a30921ac7bec1cb353d46252ae0b0803c8eb3de26d97c01287a3285a2643c1754dc6dd18c4b2e6465a6c4e88652b31f9053f419e5027094713678bf1af56049f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h865c8b706b02e9693b503a727e85b3e0d28c2d62d1e644db06243bd33d4f2f57bdb8a5d91d655f4ce6ca92948e136b336a219366a0b8bfb8c7d0534be0e0b7dae749d541af3962df54aad008d8d51ae02769b452843c2187aa8f6ea88b516d65c1ba46dd41c1bd97f6415d79d7c419834;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a422502f11e25a6aebad82714b5e7c20b0790495b09f33076b55b411b7a03628363c5dc8e3195a3fd56ef1a82021644c3b3cccbe9b63bf2fa659525da0c6a91f8cad2024f90ea556992e796161705751d94171f5fdf3921e91fd14e3e430303a298506816dd92a81f80390d0caa6f9e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a02e87e3fed998631b287870109e0946b856afd0ae085eddc9651f81071854efcd772d0149c313a517cbfb2e7f7f256ed90dee12bd89d4d0c8ca432768bac2cef1200b90d5ec645e81604885c9d9ba120c59f5ca3e396100c75c7136c5612e71c6a7d82cff1d093d78b787d23987929e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h800654479ae8fe1943362afd0f3ced1b27cb988a7a57a2e806c0f86949fe1efd97874e1730d9824229f990be6369e3a6be17e2ace7ca1059ff079e210a93f0744354c067e825fbf051cf2a6352be4eff43c909cf8a4acc870b0725bfc16f80979560d7b178f871655aa609ca2c0172da8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaddfa0e8c81f4d76f8c8121e58a82fdd5d03b20ecc7a2447f759ea976798235060bb54e3eff782bb137794a63501d982f169147058b0aac1342cb8ff77af38c578a80edfcc644470d0f5c3d3348f2017396522c39310a8c07b5ce64a4d1750a4a936cff833d87d223b331b39bedb490;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7e18c9f70154bc0dd6d93716d6621715dad8fb8f427117351633d1ce65cc12a750c38660547d1f48bca435936ddc3ee900a596bfd1a79adcbe32b4d7df95c66eb7d4c8362bb2a54d8f7cc2b1fd6fdcfe2124a9560be93f4375246cd8df832f1cce866f65157cd20e62d4df2a719b49fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6514ded8bd6d8978e6cc6a34332e16eb92240fef4cca8f2b84487bf9b4340b1fabd7f4998f5b35daa72136ce92e89d8581aa3f1169f30a68cd1de99a34ec7670fa1a7e09d58ee8cd19850ea547fd528bbaced56f3c69b53dba003b942922c74f1daca3b0ece462492e7b82b88e1ee103e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab35c54866fb99cf1c7f1b2437da260f98e4c9426565e65373ac650653e9eea51bdb3bc64925a5d5a84cd9f9054338666ee2dbef7a3c9c476871187ba1891dd81f5272dd3408483c0f83fcdbb2947aa205a4b2f2d03bed74aa1e729105f45a5afe3614abf59188b20d5426aed9bbc342;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he44058e12c424b57d5b039f5025b5d5506eb00f677aabe744574809a27dc7fb7720a68f8bbe224f6b8a1bc97c4ab1f9cdf8ad938be3fa92e496e3136bf1ae2564225b77ac95640f718e6eb3f83827f315d9eaaf89a968991d368335399d2ed142ff6564a27cf29a4b80e2c6a422f22c27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49215a25f9481340f496e35d531aca529e4d3602ef394e35073d14aceae0840d4aa51a205ec15fdc89fa858008e89c78a85731e163b848f9ad4a929bbeda4d2c5618d167499fa622c4e7988b1f538a15c15a8c0cdd9b18c49de4e9ab2fd51607c932620c0a6122e8531755fd8122f33f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfeddae41cdca84192b979311f90ae41970d65b8660a04faa33be0f2480812d7281e56e4a99b20e3c8e00647e5b7abb414f0319c2cbd3b0d0d7ab56acf894332f5b58c18a0c6044f01025486b58ef8b6915a3408a13cdd4559eab1c2ff81c4c88ef761798911ea442a6397bc991506872;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8737d062f9f7996dbf6dd786ec48e49a013c80466e21b26d4e57fa23430dc1122dffa06604d8c6fe6c1da970a5fc339376525732d102f7742eca2b5a3ddc240e000227b559b7ab72e9e42aedb0667085dcb6aec2a8b0cd45fdceb2e660ce096ffbf3ad0b352eeabc62d4abd7fb32fad7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52c234698f61f34188cb17ce90c0513451e4de0e97c2e7b1144d07682d36e3d3151a0e031c0590e1bed7311f43c6b102fe4c4b6384c71939182ac005a96698262f8c7efe4a19424795fe80f934c758f0b0b151d37028c6612454f1defba486967b013f062e744037b1dc882fd40241c89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd16da1d66a08c616bd1f8c2009316739264ae7c09b86fd7906f4e620f77f6477c0d5cf7e0e61d37f536129b1928535785dd715779904383b327a863df4a909b340e422990eba3b5369767bc45ae757940800812c34802220ecbabc345f13717ad1f441d7c147231103c3aed06b0435ed2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he62eb20e1a4ade5ffdde17f5bef9bda68fe8dfe5cfb5ee1b4c1ff9b455865c524a6aa771f28355858b6de5d4460631230aa2134baac820dc30fa6633dce6aa1a35f86b780fa41049591ce4b5b807fd991f94ba7c3998d744a0cfb0ac1fd27462fe813189515554df7f4542f376594e98f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5babc57216aa6598deab56b6da381fd680775277a5e98569c816daaa90015b66607d836b0f5d9b098432c1f580058f8d220b81634c072966ccc5fd2f47a84b213349d6678b3fc178e47613c70ca1184826621f79b6cb34e50807b306f5d6d4a0a77a1ed5e002cdf06052ffc3bec2e2f7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23109d15bf9f9600da6d4f3e08fd7542f2ec3fd2d48f5e1420d3ff293eae113fd9ee8c2e7a9712b4ef4d821bad4cdcadbc3e37e2113f623d614adec40a7e3bec7949ceabf78f0c27cc1fd5c5a790af319a711d6525d95e36f7fe7aeaa951e4c2d09a05c99b56b586231cac410dc9158a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63a9a23f1b40de6a05cf6f02221550bf51b4888b7f21cc96364360946bac7717494a42ce5fd00197cc31112ed01f86dadcaef399fafd5103744d6118602b8ed33dd48e1cbd717dcb89603b385f6a683b90c27316562d991e7bf9125b4e579fee8cd6cdb76bd84f43eacca6984ee210e64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haad2ff3fe5e6abd8732a3c9ead54a8dc567714b54fc712b71c550b55f2436472d1a3e23f2ae9d329792e549e3d5d7332f8fb73aeb8ceb58b4945a66ecdbdb82cf3ddd66f8173717af146873d1f11fbe7f6fd265b7ce696b4e37673765414949c6946685e2adbe5edb5676df87fbd8007c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bbb919c3f9306dfa8134bbd960a237415c011d587072be6e7e0bdc6ec346b921a7f2c1b94ef2eac422e925f234561224a9a7b4fee9514b72bac22e52017cd10546cfb269bc47f7f70895711b2dba2154600fb31f0b4eaaeed6d33cab9232fc72dc7c5f2a48c2cdb3ca726ff56694501c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76f0ca62eb366cc9a5568cce80eeadbf8199ed298438021d482c962ec42f7c81a63dba1346bcbbb5ac0031c096823b13f6a1fe5bbc75358f7679172951e2e41501a3fc33f5501f90c3c111d956f30b69e63b1d3aa1a31ea8bac18b2d91dc545f4ad6e4707ba2618046698d6e4d4ecefb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2445d76e6b11cfb7bc51022bed0a481d938afb5d47c097bbbc41c07f121fb12e9f66516a5f3705f8a662aa58a1aad61d717b2709984b865a9cb4fb78c99c790ccf18124162bdca7057a9c34bc0a49f52076e4edd57de66a292a84aeea970acc3a57671b8bf92efdb2be1ecef8db0752b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h486a202dfffb158226e88b4edef93dcc37522e2c4db6762acf079c2a79bfd5ab1a074e0d1194203d007cd0b17ac5cb8aa44ef0d28b155482d85190b73fa32353711d1c137769a3b85006ac5b9e66a78544d428dbd70888da197a7238e3775505da2c34f9f2a2b087ac98f01675632da3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ac13ca23f8cb730b1a0029b497ab00f6f878c464f153b759c6310441b630d5874f7e96372ef2c94932b4c32795bff353198d218e7ed9d9521465d004fac44880d6fba2f5d126d0280016f00dc22b8a2001a5104203084cc71a6f289aebf710bce5a2ac59df087319d9a3a767f856edfb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd25f45b91eb6bce9d87820d006f79809d8d4d94f0020cc6f831e16e3cf9d8587a9252935ef2d0bb0e11677bf84085824306a830da6880c38001a111ac771cd2e48d4cd82abd1c12cd3c741a9a7559db7dabf04bb79ad202ed1456eb8bab90d3cad0036c2b2f6097b7faef0df1efee5596;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4284322b3532242c3d2d9f8536284cb4b5e706999716879211f9bbb902cefb0f563a9075b5f9c1b8004aa0bd265ac56d7ef8b5e9585fb324d94fca627b9e23c79193b9d9a0065f25c86ca45f997126ca3ab3f8409bdd715dbbbe0fc6dd62bae5a86fa3dbb671af9d2e079e7ff55471e86;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa7747c44ab8674ed5ee05b2273a0f5a07fa9777f5c533e7a130f650aed021c95aa8124db68e7bac72807c0fab3bd277a45e428478a4bcf4d7aa522a139d7a2f2ed2788e844e7f8d49bbcfcb188af909bb04aef1ab8c6cce910e208d39ffbf41c8e1ae857478856f68d358f757434316;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccccadb7bba1c108572a24dc8af294c9577925294ef9e77956d055b5be8173c514c69059e656fc91df1e35185de143f9ced4e2c5176fd493c0b34116e397b754c952e6e5ac3e868db6419376d6494d78e5b94f716fdcc7883e9c319678b0d613823ba883895f988fd6e26a9eff298306f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab37fe934b6428e951a724ef58a40664d6e49308e470da560604d6f3aabaff1f99a4af1cbdb26c6a84224c744f8f05fb672f9d718c14712d7a2932f24289826f1375ba737d68351ef686a4c82621934f62dc029b668ca258aecbf96b492c7d296a03ca14aacaacd92cb8df0036e2fd7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6bdeb6832a9fda3925f0327c056239d143be2f0ca4144e443e96b85a3f8eef4d7cdb9ab19bbf2e08dbcaa0fedc46d137c538cfe5088b3303ab0f420e1e6c3d16f76692ad7bbfc1c41cda02b1e0aca3a5f8b0a1738088f49cd84c14cd8c14b9230cc8d0803710734663c2620d183f50583;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42bf4146eacd387dda92d073e2f35641056971ad6455e1269fd58640c85d4c6300a78deb5f7a0ee127358dcb245b6dc19581b21dfe6c8ddc37ffd1cd790ddb5967f1e60374bd87a5694221611a538e13ac842bcc86c2fd8db1e1cdba77400f692082e590ed93e145cb2a0760c076a0d09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefdc5df67c3c9f17e014d1c26e33bd9f9293c987aa2827a2cb51a9fea02a6deec64c62cb4b56f99609de3687c3bf24731e63aa8f9f8374f13ac9848d5691c86dcce1f094d1c35b8caa06bd5ce4d07e045f4089df5f90e8b7716da5c76752f72aeedbfb938dd90ca7c0a2f190eb5cf4785;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6216b8556eebd41deafeb22e59a1de1cf844d64eef0a24413655a1b0dfae075f41ab589c556e0ffd6d902e247a51e439c52ea5ce34c43e8774ea2803fd19d6c75e0a83b0c44ad7f664f5c82a3d5668ea9cd08e4cd2c8bcf747c0fe4b0f45c1f6a5f8e8ea2995269a7a42cb1cda476b749;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c8dd69029ebd64497707c3b08bf51240edaefbd3c662fadae3e9b72fa35f3074f4aa920327cb7ba79e3bda7b248cccf8322777d17fff59160c4a47c4b94d8dea0da7d7d89b7c3155259b7eb4a2869271e6e7c18333ca4e5a3aab417afc854de2bb94e3d9016e972598bb364633997ed3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a69a9d4843692fa5aaa3be150259bad144a6027e81b02477de906342e087aa0264fe593ac23fd2d06cb3f63845e48b60af4c9dc38e045e00d83ade6b67709292f362cfc1970e72eb7436434f6e386e2c2b202bf2ef848e40bb7e858b1bf665da4e4ce662420a3727e8d22c0b4d6e1b5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d7e917f3cdac315879826e8172a4a1a2b62a68ca462f9d161d4dcedb85fe37137950114eacc6355db98f5ea49c3f3a480fced5734152531c9273b4386ed57768641124f6491c7727eee3fe2088b64f4c14469c41e658c57d3e8661da028722233fb19e72b71a1f79d6e59849b8268957;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81eae09d5660154230f31bb547a7e88815809d4e62710662d75f43b117ec6364babc482e58d867914d38a4bf46b725f0c994e918f9f83e978c1a8ecf3ec9b67d3417003a4ec64f3f2815500186151d0770b2ddd17cbab5be886eb30342a4f2f5b06a5f62e10a9b38e39de8779e183fe72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6c6c14f3d5bef5f8620e2011cb21731a4c5753e0cf6ac4995b6f9b4f7e1ddced8fda246ff3b1ee8fc4fda0ad288f1dbe50a8ae87118eab05c2f162d5d12de2faa9fe74f01f89e212df64b218c72d95edbb76c5bc2f96743244ef2060dbe42d47ed8b63a9400b4892330e0d5f9512e3b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6a32af11d961a222a246ae4c96795228ba7d48066cbf8f50575723568f3497dae197ed47e9ec88a8b37fb3732e48523f55a6ce16c2a7badcecfd5601d528f6e81cf5fa5f022a95bef5f435197248114853973b755a98aac7f145bf2bfa61b45f647f7d61ff39d1d6cf17d2c6d2d6be0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd118c8252d3a8b5919d72d515579093bd84ac22eed67ec01ced71fa3be035d2b1afe23fc05ec2fc1d85704661dde6e6098959379161cc167d4eff87f0d7d72a2d8bd2ec914e181070803a669fa6e3b768ebbcba9dbbac465b5871af5136e76a851e966b28c3d59e35421a083ea75db3d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafa3cf064cb57d84ca89ba4481191a71874d751d11456b811210c332ad6347544b03fbe2d6ef5b292caa32eb016052a92e5a2c8dc1381f88e537ef7d136eb7183ea3f6a5eea8dfc03d64a5b35e0f27ea834f66983d3bc637b2880cb22163bf18eafe172b0a76ee35f47908409068634bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72641fd9dfb582c3288d849ca4811218a0a4be9e8d354568d0e264607f61aadbdd75bbb9d2cd1d62e5636ea657b959f3b989fd7fbd7504dc6fb424ca425bd52b2679ddf42b4ff713edbf1d286aca2bf433ea427b79ca18dd82db84479343896bc37e65254a6be55611fa9f653d225d6c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbb8fe80b5316c9d53da2d701625b33354908ce93f37b12beff2e1c487c7e149e5d1ba1d77b291e9e55d22110dd779f99470caf9058eb7a25bccf2b7bc68fec87568947560325dae63c27b15c05a732cf0b7d8ee3f54272b3ab0205c1e3d15416822738c6f6274c1bf352b879491f18dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd7df24488da651179c321713270b9534498fb970c90050d85b775a618d97edaab2323ca9259954cb24caf8f43ed0d45dce4f77087e649f128063be439cde62b8ffac68f96628269e386bb4747a8a8c7858ea7390043d4df0c49a1777f4bf5c4a925c9e14cb153ea070c9159a865b6173;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he43de2263fbe9ddf02d54570954ebac10f32d4f4bf82f24bb968016bc3afca5521155a43b6dd8fbfde75f27fd394cc6427c14d2404a4a49b2385a0bdaa65968bec98afc35335da67a0784fb453269c13b5e1c01b9377178aee5b88186a44f15e82491d3e5480826c87c94fb1da37ca48b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8adf057143301a4e972c966594342f87060c95b949475cd896bbdb2812028f3ff3fd8ddd1557ca2e9085772a96e99022e48bfa2b181482fee78b7277483b57690921c2dd768e9c5e0f40f1aab61fd4fe04d54d1104901dac53415b0eb1ad55153095999f19b6c28e3c5d4f96a0bc718ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd78c47bb54d6541e037109c008e14d364abfd39835e821f876337f05d3caa1e7dc58f44d2fa187771610bc0d993ad0fcce29bf36e9007d3ad84743e5c15be9400f732c205db6b12e632d3b76eb3821dfd03d79bdd9860b7f3271bf874e35d3d91eba97d109222503de4ff13ebae110fb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5397fff93a6cb413df9e5531df164066428de7908980702989bbd6fee1315aff63d688fae9b0521d6c1211dfb0d2b6735593cecdc2d2db986009b5b640cb7f0067d20388ad8e189a3211d56383227bd48380542bc8c075a81c91727cf53cb8f6acd8e44989e793a36c1eb6146529b4db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he24d8a29ce48bd7c53f2f16f3c3b58bbe229f6d72e1794c1ee1afa0e266748afeea9b67fb8a3ed0a24a107a921c9a91f4d663b632be4e5c7911bb03ed07c5eb981d429b436badf7f7c2e4aaccef7b1f67840603e904d621eb825b7282a5c248afcfa33704a26f16f217dabaccde4e455;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha525d75c24dcda37fb1b3997efd5a4877aa446768eda3bbe9ab8c8836fd2bf049cc718263c1a906e9a1dd0f877474f7002575158d171040b737347509861a4af86e318a8fa2f97345968994d106f748b564ef77b874ccd001fad57c24896e33533d589c72c45a62022f208cfdd8c6caa7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h855d8d1361c9e15d86c089d500a3d9e442cf303528f48f82266bede19bd1032e8a3071aeb5071c65126a98a147e687314ef8a268caed96d00ff5c072d8c8372dd2513de98671c43b64a5e05e2673fa1882a2656efc3c11e866c666573d1f5c208840dcafb6cdd59acb302047eab152cb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa0a9c0b955c7c055628d54c4a7b6da640130582a5187cd49b43c65aee0eb85e76a015d9294b631f19925bdffbacc69b14a7662d1ff8d1a52bc151f5ca5d39005de135c61f41c20d13fdc3d157b1c13eadd37e85546cefc6de1e4f9a71bda47b55014fd75dd4e12f6c79760099e2747c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11ee2d1dd5ba4fbb707fe092c11f1bbcedf3a2b5175aed860437e704f49c050e2b2a14498ab3343f4183150b7da264540bc04b3ef8f43f1c87758b37715e6820461af0e124ef8410aab21cf7f22f064e5d856c5454041f3c8b3bb25f1cad0d62ae4f1b47da9434954a70542cdc37723e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee29d11d61177cfdad5530aa1894fac410fcf8fc73df665adb7d53995ef7b8efc6af3e2037f32951f2885f9b82d55334f5b6e756b6a9e7ba7c9ad68e2573486252e6643a812d1f15ce08b8d6f776d946859b08794a398a12d129b7d396941f93ee95fb0cf4c82462520bb13ec612a15e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7f68234c6eb4752dbc4f0f9b355336765978b391c9d89c8cd96918e1685c52c5eab7292daeecd26c8a09ebcbbeb458203d0436b714e366d275169f5fb3c04d01d3b7a8d10b1a5aeccb67709705e856f666f4b3727ba460d9633cd1a473a9c73ac492403a09bed00bf67b5242dc3f58f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5c9356c478e50d3aafda8a30d971fb59213617e3ac0e5294257f16ca1f084a44fa8991235dc52914ac44697433a0586d5a8a35f48ce5cb655d237c30b10b5e9641b5de8acb56ea01f58d40f04f9fb18c59c084bda6bade141874d5c1ce2f4ca1de2f27169e8b5bc053e232bcb53fb1a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h227d28d5fa40f74bbc221f5d7a1a1420f0fd18cf5178b40f4a2b586c0b7f1149b2ad5369c663ef2fb51541e1acd3fff2fbc1f67da4c2a91c9c24f974d771ae0ffda8361e3900cb956ac6fba976d82eb2c76dc45a95128500a7246ea703db919de2cdebe6a378dc7696b66096c68352f5b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heebe81acb923395b70327e1e6ad856c9813381b53289e67fc5e9566e4246f8bd04847dab729cc30532e7cc85a1ff4dabece1a9d418097ce348fd0ac46322da11cb56f6693fe79f51289ae83bb2b8afdffd5b8df6a5afece26981fa3f747d03ff90eb2269a5b4db2efc69e1dd0cdeee8f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d53c9e08d538b235fe8c09d91754dc8f369eb22f9a2f576af5851b1b9eb1b8bd0f9061529e426739470fdedcff50b7ebca9f358be8d37820dd47c2160c3114069674acb82cdbe7175b5f32c77e72d6a03834d149028ca3a130a543841c799dc151b5857e54c4435e172c69b5c0b6d19f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h152f5b27c36c97a60b889b682bc711f2d0f3e0a45d4b65c651750ba9632864345d64078422006417a768bd1483a38d02776871d194cdd442ddd1cbd0d5d7fd8fac96ff274cc2ae5de1807d712ee53e6f6914b196b9a4035f99d7b3d4a79222abb953e4e82810e97a51eaac6ed12559d55;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h886c61d0c1e0463b6611b88eec3c48995f60416154dbdc392e1e1a9e16a6567cdb2f23e32090f316aef49912de71abf9cb767b065f624a22b23cfae80b120ea49f0246f00660d7981d9599fafc1c128ac3c8a70fe56c74275cacb592e578710f971d5f55764ea209c9279e329db6277cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h233353fe07250e4061b160bb772b66629e4718d75bc92c92b0ca84214e0ff3c330a8432c5bec5745ed6e584a30f32dcaa7b5160f015c8295763693894a6f9b17f7b04bbab51d83e1b09341fc0a7b798557c522983e106a34c71fbc25c3fe89652a333cf7e01105d140d816e88ebd54f87;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22fcaa25dedae6aff7e5fafd31dac9dc5897979124281fee70087bca61f3b3452b9cafbf648f923f5c4c88fb1602ba1778257658175994bf00998f0233be5faf503b756b2c56f35d0640d28618e5b62bd46930ee0191c048caeb414caf0dd41741a36454b57e7733bb685f51de4ba9beb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbeaa6abc649ffcf643f5b1570a30aeb21257c1be2cb0d1c1bdf9aa181a99873aaa55c352066786d6adb106b89390f2f8a9b29944f562e370e053235ab150bab4f66d07d7ecd365deed94ec812ee1b6a2047c066ed5bfa42f42d9c9c08afa5f87a18812363c59aa2df10ba051da9476e8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f121c7b94ab71ba17f5aa464dba43ccba7d1af76b9c2833357f3baef2b757ef0caf7745e5749329d48f719298e898637d115cdae34a32843b2ba1342d8b169b47042d436abc6e491f2abc59ed603c3a0fed419c099de18808307cf0cb1480d56829eb834c77c93ac506df5909d0e981a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63eae7098f3580337269bfae0e3091624826a197be549adb56138a9a767eb0bd62b4430b6a9f8f0a0dae249dcbbb1fe491fb7a6b760886d93c10d2e3fdde81f8f673bb6b8e6f009242c01e48cc38b128fb9ffb2a11f34f7eb8e741e5eca0a2ec5c2085db3adc96de0128cd92b61a329f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b9e754ca0776de3d794d424ce530ddd7c89575e258304792a9ca0d19bd2a06dae54cef8e6cd050a7655fe46e99e12961501e7a75465e237beeab57acfab68d972f095bfe376369afc69535b8e8f8ae2cb98a762cf7a7a13c2d8048a8d8dc459c4e3d219fdbb831d8c6f51874633c6383;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e0ca19c99091a0ab7d30ee0c0b0267e4fa30c22ae6323a7b30c6616033490e07fb4051a5f6c5aedbc329789557daaa119b69f327f27a7ac6aae6a41c037cd81c452a9f4256c8399b69bcfe0e49d9360ac290033fb67239c5e00157c97ab72ba515fe0943f8e0775cc4d395d94345b535;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4ae48048919fb3d112115780fb1ab6021548ee6aafc8c4d601d76795748fee1a52376967a247c50efbd7fd71d0a190492b9891b9f7a18e2364876289873be398b4559f75f899f45be60b1de42dcd70c7a7ea8c254522051cf87d783537e67353ff938dd8881399fda8d3861a9d10ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d53f9956559598a04a6c70a5dbe6cf2cef384792c2a786ab5f40cfd488cd0f6082cf67996e920753b5ac340c9d50efa4547dd96963310b6c5e64f41a512c1c12edbb52ed9d7f16935f3434ddefc65f731d9418544c6ce1a46ea58e1e610afdf5d3b901a1fa53888bb8e7da7bcfcf8740;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88ace13392b93ee5f6501881de9bdd812502d95ec3e19984c1a3da595cd00b3f45638f8a09445df0e7181ae787d07852a3c62c9e7e2e73e6511b56c8e7af67274389ff73e2f85b14b52965d4110cd39f2885f7ad69d6bd09edc602252fcd15f0eef00dcb3fbee82fab9eb024e7aeb0ad0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae4a1f2e179ef37c4ed47c16dcc5072e2a970407195271df1d977b8c4c644e328a038a2ac60b5ee189c7169b248577489eeb04ab14ec5a001c626e0775c0610b39e598e86518212c7db1c7affe60247a17eafee719f24876133692ce5cf0a9aed24083ecbc3fdaf6e2f92ff6114a55d17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4747686675afcbec8a3b81901e42d119447a1e63d5316a669354da53da101c03f09bd7d451409757b26685a5416896811eecee6bd84375a5095151f7b1dde523de3d12e8193a90fe6072f3388fcb50ef39acd10afcab46527b47b3dcb38a3ac45ba6fffe28818ec475e797d380d168b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf56e6bcae81be6ee449a4dfa95277d3247d8f8eb43b525e668aba70749ebd58735698df93b586e37226e1dd667cecf8e41dd8abf89b004c2ff77eba6a197b92a75e1ed635f692bc47e36ece59701eaf405dd70a189bf2d6f608740185bb8e30beeb10af858810e2d1e29552ab6f57027;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde39d04d1c6450cd3390768650c55dbbd15110022a1880fa84dd8ef565a45c2becb69585ab6d741e90b7cfb2814d3b879cd010066f3dad71c0644779d6c2c750f4d225e1ed39ec1b5afddbb59c13aa9895edc4fdafdaeed46b65c0bac007cdb0402cee27278e1b63c7853fa087c720c1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f27808e407cb68250d92f504c2538272911e3884e1bd1dffa576932873b3727d2b9d0fa4e2a31446289eaac5c97c94d999161fe1e6f8b7747a4b9575c6d21194cc4a4f85dade1522299aab3139aa1815c3d01645fa7f11f6a3543424f1fd443eac2a8a7cf429ddda1df8349c1fdaf5a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h245baddb80f94c09a0b26d12fe37715efc476e3c08680727d601c866eff482b00ee0502a1edcd829e217166a08b62cd5d67b70c300ce55fab53585b4bb448441b1d915eecc71339b37988767aa222a216cb6bff301f20ed6ad6d701a6b72b0560113791fa9248475310b6c4e26f4f180;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd09e13b997bd28515ff2ac840c0b49340c62c5998cf24d081a57149f0531f836b7b22909d205416cabe6e089d62cd6b73b4f9652a2cd1929d241f7a2d7bbe9c458003571826a91c8a1af42475b3f561bd8896d0e5ebf8475b987b3ea9874acb38d64c11ec27c3cc68cfacb943801d34d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89e95d1497bba48a859e43605c28ed2efabe15c37456918260f29a5fe8c68c311de0184543f1f5a0e5d7de28cae3002497585904fe0931b80146a55bf9bf90e245f8d729d4fefe7f40e982c0eef918decce790951fc6619e09e4c69fc29effb029dbcc8f91b3b20dfaf35918575eac4d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28db7a8b07b368f34337e236b9ba5e197a8c9e889250a88db0f5de0cdc7e298d10122c540306a8cd1f38be01c045e012deb372444726c799548645767b8837a194a8431c14cb09b757632b24debaf59daad33cdeeb2e2282f609acffc97fe2cb64394ac4c6ce059c958f5e066b7fe64c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b9495114816d44f7c481f1cd3b14b84247ed9d38ce39104eed8bb0e84c9e8e5534e7e95dd7a1e0114c41472400378339856f15a376205d88eacf0d9a306b14bf40c654539b9291b261872d590062a198c63f60ddbb0860d0ba19c8fef25e7cd4cad520a19c32bff8fcda70cbff096c3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b57a5bad3750280ba626da11a09a404b079eeba0753c444d0024701a12a01a51a99d8a4945130f8eee068fb9e5f60904623986ff22f43c7868a98f780f788fe77ec70a4b0d7db137b6a070944f2490616a63d7ecb5934adef07f41625c067bdaaa9ca1ef7c0eff3a859928552ab93060;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebc6d4945f145842e10485e4c3b6a5263fedb079837d4e45c6544c95ba100dd1207c503badedb58205e5d2e4559f00d4e90831a5e3214b6372739c5d3c4a9b21b83e39707a99829ad9accb6c2678aaebbac9e64f50b440d44857535a148596505d67a2f8fe8d66b3c830a7d9350fc8bf6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ad20e4911d59fca0071301af76c09e0057657b61a04ad4b1a3c7b5d23bda3ce7e8a459617ed2e4da0623abc34793df6a83a7c96925cd5a7b0df4ee7775a0a4e3009945d415648cfbe02e692bb02033ce6b2d0cd0cfcb89fc0d0570b854c8bf3f9f625f7c3a762919924eed61f7b01b32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba948ced9ed0af112369c37ff8c46987c94526498110c2e16a4a2263b1f8730c10b9b8d285bd713b0a3a081d0765923276dc8c3a8c6ebd9d2f1502c11a29a03b1ef7fcf334d37de9d872794e0eb92c017197a801833bc3166afa75212d3ecf2bb78164ae09f77c2e347eb4602b968ce4c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45ea3e518d4c7f32c26709863e429f611d26e7ee91105b5a759f8cef27eb555a254fb2cd58e46c6867342e520f6511d178bec249328c5a9a9f3defd9e6b68bca2a861ebc75093c90aaf44427bb5d3e43adad0f5906c553275913da4397aa715cd925343e676b2398d5631d6af9a583b55;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf63dfc7b9ed6c84ac43c2ab19de9381d23d6d9943324bf048362e8f0df5f6f33d58067905c9921cafd4f81e06a863fec54999439d41fd765c20ad6aa5fe80669f0ae8c097e99ff407a859cddf431d15c5558c260ee8d64ec6e2398b10db8acb42f26288d20a5216d8f5c2a4ab75b78116;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h782f0d69e9351d705f10f4160192a46b369ccae5862a60dc8bff5f6cf17c8b6b1458d73b937c6ad8ca7821f08548b5c1eb30fa2d7f6ee50d43357949274652b7e2effd7da734e8f519a51e7c16160bd5885d82157ce08d52c01f11e3b54ef2c79be79ccbea4a52801605f3e79efb7974b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habbecd89268b2241a77620b78d57ef67ca049d618fea577d362af5b722efaf62433200f10a2a66be4331c4b5df87ac53552f1e07c667b2837e21478f1a45ea7a1cdd12182c91f995237c0dbcaf50930be02e675d66adeeeba43b3ff080940c08016fbe9ad2e4c3f6921bb074748f46a0a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e6102b9998f9fb1fbb38870af3516b9ced6711ce753c0c49039c0cab1042af52bfadf2c8140d165825f5b5a0dd77fef012392ff019ba72eda1759a1a7054a337e331d66e08f6be47c57a83dbd7172f9f76430dc405bfb6a0b9d0308daf4d0270ed275129af39c9d12a10594b5ffc479a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0361a9e72379b8933987ba3f6971d2edb2767e1fa382fad313af5d54899c15222af7974e23b63d56ebb693237376ef718a27cd0a04b15089be01cd4604f7c06fb1c636c1598910a92fff3ff42aec7125f0e4d3c583785b090beb926dba91247e9e5c8401ecbb6483f05ace22314f73fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc12ae169e7735a0795dcace90dae3588eb0cc69b852373d63d43816d0cd0dff389749123fd4953b81cb38e1eb964b21d8433ab3da39a30a4d78b1bb35bbcb13a559c78c3ee81d04e34a8712623e07acd98da1158984a3647653c9223d1b45ac5145abcb6ec9f35aeff93361c3e4895d52;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3838adecb445ff3c3c58a75bf6b7c5b705184ee390f12ec870349981fad82202b251f900772b1424fa56b6027c93d5e80b60171b3607a2be2546f4954aebbb03e0ed5846ffa0321ee4b05206cfa8a53fcfed89e449c6a5c27d21732d549dfd66b5c596319c44202d0f607b4f05b848f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6e9cb28911c69efff6b33d1530500d545945b171cb11405c9e89b3a1d66d125048ec96af52b65ee983dde2c0f5a31d0bb3888da051098e205d3505203b0ad14770e3a97dff815b402912db1f4f37eb6334dff189f6cf3f9227f54227186c89a911081be9fc7c7e1cf64d265d3699646f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he71dc89e452b6824ca0e5d13de730bf7ddf6e428585734d2215a4a2cc003e754c97e7970da3afa3735db9c6733316724bd934503fe99f14e27cfacfbe8509ee79cc3dce14904a37c390b972b104db26e694a4a69f297c5931ec02a9535ec814d23f021298418c3d175a09e054c9c97b7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9ce1e31fbe35254f5aa247796129bd448325ad7930f7799ac2bb7eb64bd0ef33d89d2798fd9fb45b568a351b84a8b22d42c32d17b99534696e902e43adaf6440320aaa1c78e99c05dbc54a8c3202a0530b08b501ee48523a5af02d3f6fbd4e40f17e63f6f30f36dae47a840e26ba0df9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ca9647ea168c18f900b02a3f10567efd7e23052e2f7ddbce5eafa7a7bb5ac920e30a1a04f017038a331d6330972152071ecc21672cb1b103684e416d82553f4a4f68b294c513d332a0c75f9d8b35e1c41a6a1e2a8c10824da447c7bd5d9242a3ac655bd351285749c3f47f62100b4b3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda4828a9404439c595e920f55239d3321b01747c9ab16802584146d36f4b7114ce22b932d8f807a0bfd47b1e7e2a07a1cbe706f3c54685c9de163f08669f91556da33ea1a92146b8ce30dec52352ed1d9cd999158702e78cfdf121d1342a448610a3c89d91d21d4c2792ae3ef820c1c88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd10e65e29679b839ba9a83a9f8d46513a0d2c4770c0ca78e99ba6f5c74cc366c69341b07ea04bb1cfdc69737971730dec225c6cc45487ab3033d86502251c81c1d4553997898af7d7b475016f42a7d4d44dafcee8e68dc1d195b1ac5d6c2fb414e76eb8453f55607b0019f27d9e48858a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15c21d83b3eea3e8fa35fcdadfd5f741a8c51e1807760091fed94b6b9c43c5ee7526c5111ea535612b4a35509df3bde04aefd4f00cf62b3e3f2d1d1eaa51daf26838bcb04048eead57ebc399f840e66318ffbcb6ccf8e3564877d8a8107f82d27b954eff837ee4c054805477eb94f0293;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4974c4ddfac0839772985554b21ccc4bc954c49882159f351c87f68a4caa4c1e28615a6ce96c92f7c73ef834c769f61cbbbee238081a94542030948a845d4a412ec3d2c6a7e1e52d410df9cf6bbdc53e27a494f794ee204265fa0bfa38d0a8268489098a8557ac74f3e02945951fc6ebc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h564ad7056bf1d57783ac3231acdddd3d2fa48ee547858f1465970c376ec84a9f7f15314ae0bdbb52bf588effb307a41abcace66f586dc9b6233bfe8a86290aa0529c873f364881b62f3a1941a79b5fd75144298a3d6e8d4bf1c13dd58a66a4e686908b977a4f735b0dbbd7c332f6dde5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d2362348e62551cd2cb9c4131c46641aa4571f578460f60e907961d49b6b5e04f0e956938a12d752a6b9553eb1d7cc8486c4f514f45c5e2d814242ea14ebb85e20b24a0508d34385f8a8aed64f84ea9ebec3ee35a00fe6ee7449cd86d9c99c51986aca435e5a013bffa56a0d007d9458;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd63d501660d65fac2c6c5bec18c227e8d48907494bb65bc1dbaf0883eb14edd21590fec1b793b09ecfe112e80fe7def12e2d308096ffad803c6ce23a7bebdde1ba07bf4f575fff6fa9e49d02e4d1004279f4da59e4011dd9725bfb054d629ca4b368e69345d5f1253941e2a7a6f3b6bb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8262a8339f8c0ecf539b2fb0e733089abf7ae3b0006eaeb35ecb41a3fe2a31904e66434cc0c55da342df91b0b0b95ed970ab403c977f25514b0fc73824e817da3ec8773a299f641e59952de812e181f19cbc93ec995cc79e79de04aa569b4dd77992cecd2cf28104d88de40a0e0690f53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77514db4f227eefd95175f563a41ab39afc043cf2e9d28b9397a27ac6275fa5fbfed5ddc490892c721120f7b5f8ca8d66389d7e43fff360a81fbc9ff5605faf5287122b02dfa7c328858c6192e7259da41713447460b45ebfa701da570ac33e0437765451612a2bea644999964770b3c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf93ff04e7d5042daed0c610997c638e645ef8f719a266a8bc97e1469d192040e8da54089f71f0c929cf65835bec60df9e92f846e815f68d766d3fd052c78c96334104a3803c8d6604d7c819d036b7d571928d327855694de1c39bee7f70ce68b56fc5434299a5bf6bf667edb3c987cd4c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10c49573a870fc799410ea0e7e121cd51f072927a3f31777120eb28ed9be3bd01fbe93ed08c58eb1a41f307182dc3fb65efd97b6d005b66e41a1b020f8ea900bf48e85e41f5d82c24c44dd0ed26d9e0c000ab221ce22c971924d1c8f1a78b737507fc986798ab038caf427e7adbd507b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde722fcf7e1f76e1e7086ef2de720bc48447cf6f045a687532a7663fd4b8ccb383676faf2d2ed7eb2eac10c25a307f2c8312e25cb5937e68d7d313fb5d28ac7b4d07cf2df68c220cd7a43da1f54a092bebcae04876126b32b8d1357b2837e8dd4434e678daf1b5cbdb3a0254e674c0714;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ced8b475f0b8027d466b09792d087bac3908004b0c32c7541a6b0df263a39b63e7f5211d103a39b5c97fbb4fb5a86a9f5fed6f4176edae1d247646ceddcded8647b052c6b4644847399050c575f15ef29cc4a0d97e30355d0b233172497db1799d871aa2b16ff71abab18ce6f36bc9a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87cc0354c62328d84fcce856abbf8dbe762549761f7d72fdace6bff87f3e580b536ba2b00b9197d921f6a8efdc8d60ae664c738c3d4f6a0d4e63c9b1e46e054497a20b06db4c86f510d8d15712d99b57e2fc6fe2163c1c38c99fc93c247d1e235fb7562980c9135a78305f267d4baaee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h508082cda7f24f2f35da39030c8d4a67689e75845abacb7c600b838d16722839a3bb66e26a071403a0eab09de5fe0f940410fd9d405f09c162e1d7c6010f9474a2449f3616697995e8e79d6fd977d5f950c0e092ba099eaa6f0fcaab2116cab51dab098f39f1316498a0484bac547207e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee88141e3e5208a6f51f8e9d3ec0ee984e01a33d39d31baeffede7343bc021e8ae147f69e74395701555ec1ba14cccabd563850ab85b6c93ad9026705c7b4dc36e9c6756302a5e7b869bbaa971756e5d7696f8a51d91a50061e807ae7279eefbfc7b61ce41b2cde411c1094f0c9c5024a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heed266bf8d6cdae1e96fe7f1f3870a7addefc4fcb3f5217d4d6eee4b5ed880c69e00c7782003d7054bc066ea2fda837bb6b1611a9e02394ed14cb81ea9585fe667ff39f60091f4cf04eef417c22390d5d2c8aa0d5143d8d306d000fd2f8b54a958cad912852aa2cdf6f4f5d1c39ec5932;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77db2a76ee170e87673d446cc8e7f46c47829237fa7b56c11349aa7905c513839d7d35b78145368d28bbe27c38a6ccaf64c37c3c5a70467ca1ef1fbd1fb19d024772d0618c5cfaa83329e53a2f7645476fc06fafe5303d69976ce2b38d952bfafdd5198606b2c06c39c86bbde615a7bd7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ad9232062cf3e43d5e5a0d9681ca78c0d13e21acd61eccf71f93c4baf935e087e4e5cbd3926e58935213705d64bf62cfd2d1d91b9261fa8481c916f898ce0429d427b9ce659c69937c64610ff3a1752fc8a98f4b24263e40bae8dd4c680b43db474aeb1777d625188091b55d784c94f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdd17f34df0c386de5cb69f758d28edaeb6f7827f935abf8e2198ebf6a06126ec6f6ac75b976988df29a40911a8af58ca72bb6351cd745f9bcaf9dc4643cd179a0dea251912e910a902bade4a47456ad029eba307fcf435235c750d63a1d31677f9384f8cf2f83897bf53dc4669cbb078;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf541f99af5bd6ccbd1d53325a7b8ee0c05b6e1183b62b55cf050aea9c257d87070a8547ee5f6967f5610346d47a18fc99c061de90350c11b97452bb653755d2efb75756494ac5faff5a13af06b2092f919f2e8eb4048c7640f5c84be64d4c4e21e78f0041bbd4a049152a0a5790eb6671;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69e526dbed252a97f3b8fe90877d4b5a83bd29b8217f36c51c9d950c5b06db04a4fc842594123a88f7c7de6a8d1b00e7a1380a0803d1032925fba62af9db4e9cf5caf682b2b4641bcc3882e853f9e56a0ddbc175eee8e92a9f840ada84678d9865f271e5fb2ccf107b283cc38988bf9da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aad11ff2e8280af1b50cf012711a1fc2671f83836719ccb19a92093441a372a64da4463b7885ee299db62cf82c3541c0483d9ada4e5ad77030be9f950d15cdadb42c92785ea7d200901fb52988dc1c80d98105c53e6b44f6e41b7530f873044ccb627fc9caf49f56c3867fe3a3846ff3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d59c70f03ca6f7fe5aae40804879f78b9023100aa4d1148824b00e7fdb583abf216c1684d083daab11e559ea13e389f663adf7636a71102a1b7cfa80e230a6de69ad9f845dc6a65bb3580af2a24d388ed72218d24eb4842cbd6517eed1f91919814b6c73fbbd2796995676a0ad066a65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8389c57b50421ab615a5858f50387c5cb7de926074037288b4a92e3456bb779c834a797ce7756dbab0baa4e5dc4c3989ff9c0d2cb07f732297feba3bb7391b3d1e55c0bdb613a36d6937ab8e2578247c7cfdfaa3dfaa11c9e19ad7ed9416470fd7964ef4af3d008e300d2dfbca27b183;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a10ebea062abe60ef99969055d92cf8c8621c402399f14b76dcdf3fdd6319ea01c5e3efcfa044bca76f8ce99053d6a0f16d930518b26ef905c9eabff85d5912dd01a06985d48eacb4f8b9bc9cab06502ec03558c7f8585b2f6b2eeea7653fbaf27244f3e6c73620398933146973355c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95164bbda8e77e014c7121da4b29e2c70772a5430b72ab1c9094742c8b2ee228f2bbf5932733bcaada2426db5211b4b8f27a4f256bf362582cc9cca51613fdff3ed026fe2a60138d1e35e14b9af69619daadbd59f15d3fc8ddb2abd126c5fe9de56a83d62254ebc36074a877290425439;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h227105b6d4fea0961cc3b950c3013f2a4b0c5d3c4fe84c8e183c67a40cad2ebee7ce9852e7ee5de4406e6eb4eb0545f75f91f030d250b9e3be2bb872fd612b7d9e76ac6cb4c4e4fd3ada129e369b56a2d4875d642f1befbc7f40bd33459c2c45189810efdf8df4604c0e1e36bb21f6d9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30cdff4d39589fcdf9511775be472a80b9a86e61e3a02bbc6591c397e1cc97c2d4ae1a58f9307777b65a32e4ffaca8b114ae89617c2e933589c3b4c3795483ce6a1068606f5cec185821d613ffa2d3c758d8fa9a244b679f798daeccc8c84b9a5bd27ed3ebdc00e7b4c92e6af4c10d87c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa12bb46b2bff9ca70a7c4d921b562835168de77da7d36b86c04d3effff6cf60e9ba7485c7eb22cb6d90b5f0fc3d896768840347db0e1dd88ba3c93f1479d9f596afea2c190ae4ca41e5cf5f080bac6c471e7a64999917a6ee16554ad16ad38b22e026a1799f9551da4164e16e5e9c37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h593a6fa708abdb0d97951a03c13b9bb788e05cede99d70ae1934a576aaccd66440d1aafcdd07bb48fa5b3c3f002b3b62efafc98fe02d3bb2f0e09c9c34ccb2211c7106b3a49bba2ec80b1b30759a8d89ab6de8443164df78cfed8ad1ce9acdc40c4a8040fd4d50605ac6a1079118fe053;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3873ae7e078a4cf0a3364c4b991b3f3bf6a542feff90a88dd8ce05ecc6445afc40e09b9a0ba3e5be29be208b71336a1020f574b3ff79148f8a9cef15e68e6858cba3efd682b8bba114bfbeadcd2944e867e578f92d66641c6fca354c9a3ba60183530ffd138fc4807e8a173a60864808;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26a29d5adc9ab1ca38eb66dd29a192a1d55a8d341b08e5e55699c870ffd0eb3d5395fd48c5489eadc0388b9cbd75aa24959d7cfbbc0e584cf7cb011e63f8ca64cd449d2e9be383905c6ee29e96b72cc2daa8a6b481a2da3596234d5099d08e5684a86a9818a1453a549e72bbd7067c31e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f0e41ed7204d321485a8b9341a11b42fbc774b23751c060ce90297a8a2141a4fe50727a8785c5e2994984c7a1501fb4dd6633a7cd05f02a71f8fef242585a4dce6f04aa9839262273c2d3e50f0e0913a6ed936d6b17adf30076bc00ddda87ab95c5465f13bee3a939349139db1c329d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc30c7b9b6cc1fc15e09f0cf4185aeea9a27188b0688e68b5739df0a7f9af8b54fcefdfe663a18b560237d0435ab58db42308d6c435bb2b1ec436e0642a840ed198758816103e30d8c90992b9ad79a3dd5b989e2d7431722eb312493eaeaba1cd9d465e30374bf05c00d453c8cf538e5d4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he47b5194e13a4fa3be3aa85c62b7a3a143a0e8caf3b636ee8bbc1d1027adcc346925030c9b975ac3d006a0e1a7f3bf90c20e01768991b69f9177a86f55a3eb1ccf22aafa8f977fd7b70461d6c390b09e34ef2f82122be9c9c61975b40196860214d083db72861de313f9bcb5b60bad1c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc390e71723fbacf1b23dfd5eede3a1ee9e50016c7e02fd6a0bfc3739acc20e65c06db34914f50a83a02d13483ce9a883f1ef93297d2b960d50dc50b6a38e0873ba4d42bb0041bbf1e86ce145c80818da9d6503dd77b7ce03a6c00f45511c4d407dd0b3232cbddcda24c6ec905ede8c9cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97ffadeec3ab570639ca9267fc3b7b806778ee45fab5aebda33fa1a61b1edf7832d38095e05cb34be6f3d8ac8349464940e853f5161cca7b4e58850a6c1eea1d58fb89afa8e8d6efaaa9d596372be25caffb31dd8d09698413dc1d749d9ffec78131b1b6ee408dc34bc32577599023e68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4218510e993b709e01a26d84065792672a8856418840ee443070273fe8d0462fc3a0994da697ff37fa3ffbd430c731404ca4dc0fec1b6d2447ff373c098db0c35645fc51d9b1c208896d44fc2f63f5993ee95f04d5cc23efdb2b217275efec6c78d5a1c42244b3d6fe188cab6e79017d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffccb1d5a1c324474c5bbd92bf0bbcd15a637ab7a470afae45d152939f8478f0704335d6f08a23c27b4a30ced4bce5afbabb9bc615686feebf4608471922d7e18fcd558d00d5667611a3c6d6951b821a82053dc9a63ccba6b93500a9bd7071249888e2906ac08160f338282e2fb5f2809;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf597a3ca135fefa732c0d838d59c774831316ac0695380333cc83a00a88ee104d243b5a68a89554648b7cecdde755eea2fac31a28e0a6cbc9cbdd6e55a385330a666c9cc22a19b19fdf10856f12154a617227b541abd0fb06481b15686bfbe9ec8a782c158a21a5effc22fc82b33e563a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f423731b7843c7c9c51ecbd94c537b6e3461edf2635c2606d29419862861d8f82c75ef634946a0b4e1fbee7c220d0d0cfc59f148b640ffaa254f26a1be7353b3acfd0435f850d29cf2750fadf788cd39f981061d32f1e85fd77cd0c1282d933365dfc5ca926474e768a075785f5f4f94;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9285a337812334bb5dbc58f0fbd425e2005430b69ad79ab479e08e9c607669abc21a2fe91b9cbc510f47c16e0e10f76af4098999b647c1e76c9a88f4380e51c04074afe9a09545250329416117b756ddf7a4aa2bc48c0ecb3b7e8d071a389bb1c229c9b4a643fe1f38ec02f0626d66d74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54a16b45a6e4b41a4669850493bc0d3284b118480997da36cb1e5625be38d62c838452eaa473062a3374bc76f7bb4846d3240672ac16bf4d9480d5e6f0b0b42936bb59ff7e05f0670435bb4f28afee081ea1705d5071f47638449f9c05c615c1e1c1ecb9c9dd9ba6a59271cfda5ac662b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4db51f1707f90c31a9a85450019a3d3ea07c2982363d76e325f5b0887936bd990364be4e305639216593e15194c7e3da71b213d36227c0803d100237fccb5bf211134ad0355a59f13dc03ebbc3d52c20265c054d1e606b85d892e3c728e5c5099081dfbb950a470c5ea3b48943a31f330;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9125ce8c0433e0e6677dd2e6d126e6d791f7b95b08e905f6f7200c1b3aefad5f3e167c41e5d596f12f87c5aa2bfb8903e59411c872c043b586b617a8155db2177949c4a23ede0e737d65313d715ffa35b62c89a34528b46aae653c5dc0cce649120710c3c7755853bdfeaec222b1764a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c0ea54f54aa2d5f727a2dc296a06a94782342630f100f3d70e3de0bebbcc6d1c402438743535dddc928e5d970ff392bc38e8c692e59f2f53622b4e8fb461efcc30e7d8e65b875278970ae3cc89dc4ceeca37f14077604f4144e9d2f1808670aff5ef6041d2091ee442e37672bbac4966;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18977aa08315fcf44f1513a6ed63f41c7d9e4a7fffd337ce1a328db965e9b7043f7baa04a12831d9b4789c373ddb07372cbcc225f5c76082db68fc8d6b9fc0344e954043125d31dfa58504000830bf73b42a6150d8645467ef61d70e97cd1d70328de142641472703747f7d566598b6b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1265bec58a9a1415c42da1b130071320648627b0f0477f3e3cfd54c42f1f9361000976ccecab33768224557fb4b101ed45f3e63b486b33f2f43bfe32151358261ba75f712506fc8f195da5c16ae2430cdc1c79c3931fa88bfd8adf37ff3d1891ebf82cf5438755f0e3cd6428a1c312a1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha33ea4f5c739a42ac7e796a8cc05c0f8f10e764308c3e72262a6a337c9351d903eefd08932113a329d747cd6c8b323adc2450235d6f441dd0bdab3a43c649c7c7228cde3d3a99d8f9126c82f91ab2010a0b9012eff8cecc9e1273496d366af9337f3c3bbf9a0063840d5403929378937;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95317abfb5e75effbac371e5016578c566f2d1a8f6bb38ab44d8073926034373e0ab73c62d7da043780b6bcf1e75b9eaf0f78656186b8dd71782197ff4862ce18c915162b7471dfba31d3887400dbd741ef6c8c58d49100f4510ea0fbf584a5ef1e2dcf6bdecd110a597126aa06ffc9bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb69b2faee7701156c3cf5413e8afd48bdcf02c88b77b6f69f237edc154c5f88c9b361d0fde8491e02044bed4ead27596a7984956646919a3cb9d0946fff84f718dbf07eea2157a8ef24bbefe1ae2dc08e6c6c1dba4cc848a94b5fa306bbee04dd8dfa39ca57a230b0dfa97f27855c1d69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44572bddbe3f66e5bb12f757aca05bf5fe055aaef31dc40311b81dd987700a426a2e6cd013ad4a5bd8289d72c2d2c1e1d23e85a77987bc4de984c3147c5026efc67a6de69ffdf469702b8fe9740ae570f24f2ff76302929b3fff1e867a450b40e3028a93f090c6de2d59eb79cf773006d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa1cd65fa537023f27f7d497adea221bae37d9bc203cbfa4f022b63318c0ee2bba3ca410323a26615f65ef5855fc39bfb9a8ab141279bd4e88bfcdf2687f404b4f876d2e1099e0fad9eb9708ea8fda081d4881eaca7f5aa55e0de34ec8cd973c9035e5089a0cf2a5c151d73da847c2853;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61fd13b9d29ac44397cc6b9eaea4ad13a11b1d47e40b4568657617bdfd1d33ea588c622cbd63656601893825c314a8dfc8ad8d638e0ebe8a3030bfd71e961254d67e4062c223036fc20475c7331514d563fead8d2ca0d68bc3c411cc69d0399b69b6e64d765fe903437f6fb2a27554fc2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdb855e441357435b20a75bb03d700fb6bd59a4d690f9a8c8430203d0a1d2437ada398b3765bee5a5a9b4a56681900004f885496daaa247bf24e23063bcba4c29df40ffa23d966185965ed958d30d9aa64d818dc598071f9b85f9fc40809e9c2436bea471a9a3d14518112b9d29a2271;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0bae0332cbef6a558894dcd6659942050d56b641aec6aa69eafd24b51698749ebe38f7616bfce11f56beba35373ad4de0b5e45a24f2a5de58a8fd53158708c1bd987c7734e6195cac4a64be72602278af6e6f76ec9dfbe8841ee97727511bbd829ddadf9dd6d149fc578f6d9bc082cce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f65cec5ffd45d5aabe62e7a2a98f1b06f20a400c2013fe5e02ec6ff28d554ab09f18db8e98c36ff1f95a35381b11791254280647b216cb4ce23ea282b4e3bd42280d9d883f84fec66e3c7aaabb0d0dd8368a76105d78fe88bbb4dfce390eb5101bdbfa7bff34d8ad790cae12d543160;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d116946b47ad854d71201ca30382bdf059a5e14b1c8e8d0bd39f301da4e7f1247d8f0ba37de49f43ed4d7528421815bd7157ac3312fc36a5cb82206bc75b86c61b5477b485a91f14c40b1933d92807fc7873a725f540b1d3f57b2e9b9991859911912f26a8409bc2e31b386657d27999;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11e8debca7d80602ad29c6f28113b897fc81d9c7eb34e74778111fbbd0e7eb94cb608bc26238156bf047105e93f7ab0f2a5a7ae07269de733deb5efec6ae2265061ce9d5e4d293730beee289b91ace5409b36005495674a03bdaaf6b3dde9c635b82d4e9aefd122869d30eb8c8406e1ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae03f1e4dbe3641823b81a7eea5a3163cde96e182a32ebf692f8e9d05ac77ee4feb1dc2b1e4c7e1e22dd256dc35205917f855ead6ffb50383e21463fa906fcf2cf29cb900637a650eaad580d5db91809dbd5f71fb60c0f050a5457227f315f6c93592d702ceeed525e186b43b8463950a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf880916297bd53e5dbf5c065b3029d28fb55869b0a4a8931f1607501c88a9486a0470b01335606718ed534c85f99020bfffc4f8c06b8a02670353c4b1aca9f1c8a6c598f2cd321ee5fc21e6d1ebbc50f0618133faf4e11592d5deea278b4630cd989330aec0f8bc0a09c4f8b2beca84b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27710832dfaae4dcb030b29b2ce711317f252fb026d3e93e6be30c105e0cbad45719fc7d0aaedd95f7ecda78a8906c276866fa89b0ccf651551ba462f4e7ce0ca1a31d468d5b6abae574f84eb45501487dfb19da2be9bf778d2369298f14e30b0bf8ed4b95f2edc97c0cceb571e18e25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10badc9c9b11e24320bbbc350153bc2f7f19798501c10cd6d99f60d94a8fb5c64f2d76b52d4096dbac8951001dda32bc0b9b03ef230952df4c7591e2b4e99bb592c7689782347cfecfd6902c9c20196c55a21518671b590119fb5c006e658791f32d1c27507a2d858b4c4923e42f61049;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h715fac481f684bc4f12048db10d0934588779dfdc78e829ebed8078f0ebe62f2081dc9b97191a7450172714cc9845a6a234e7f54d0b254f1c19db8f0d3c9efd6a0b992297a7330d45fbbf3343d438099778fec71d7cfb03ac0cffa4504e89b63f4578c942dcccfce7df0b7ce582a587d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fa7b6d18d83661181ec94be75efc44b375a190d9f01a8f5a079370da1021fffe648ff0b69ea20f1172f254c191b6484002e243a55024676cafe5dce286c865c7a7fb09f4f4ac8e667f133acf8b9ecd4feb0968b6db62fdf577794156fe7bc4c96ceed78f35140cfcbec8d24899f0967f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2996b89126cc1ed52e60425ec13b720b3ce4c94d638c23e387cb5cdd9cfa0cf74bfc9ff82394df66d3d546891cba80cd30188831320a98897cc9ccc15a0c7093e5c16ff3a45e5b1359f71a970a4e57441dea915387d3093f36df6388006614da67ef1bb07d918a29a6031f44b54f221e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78027b8249162992017738031400108aa8b8c506f989a0c4596c07f77cec4b56673cb9bdde06894e1894f502b8558113621d26e3fbf4d51c93c6493dfeb84b8360f4f9ab017126ad6ce56f208f6fb0e69619cff7754a0d26adf494cf9bdaf26e840d3d07e5a698b6899712633204aa388;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h377f855c9f3168e8d098ed5670e57fb1172f0fdf98d5801d52dd2c7440f320b171f7e68e7e9af29bc8c2c789ea560002aea99ee310423240c1eddb2adf6230fc483e1ff78571c0c07faa1a3cb6c0d955c4b3bff053f9c31d50e84a623272fc6758898e81334f5affa09196e59d368ca5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1136220caed3f775263b9c4efabca50b771fc6211e1be17548213fea7396f8095335518a9269158e0a92a9c268ee8513eadb14fe0437058d33cba02105259fec485ed77c28bdda776f9274ed61c4c7f8bada8524bc7bb4a789ee8e4caba670b0b1ec4970bfa4647bbd79f51c214722e63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h580364e3cace3dd3787882056e0788fc9fe6c4e13a4278bed7d127d83335af56173500261c169eeff3704e00c9abb29fc1f0623f8806d1d64ca5f03ba6bf46bc96f9b3b49ce39aff30984fc5bee92a611d85b23bfb9ec90ac464122d5e2f72ddedd844b52feab7d555f4912f771634cc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7a63687292fcacd2a07315e6583e291fdbe1a8e86b38c0024ba5a043e573e850a034ed015ef1550874596800ac89e8b31d7df810e2a363e26ff0fdb51d0d5ac1110c58008b036ef13eeaea1f6c3b72b6f41eea19c2ded0ed04f86ceb497840c2ac32427d789760dc42f8f72937c89eba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf05e02bd7c79c542a8a2bb70494afacbeaf53900c7ed5cd0d6e710c47b3a722a37b212e341bb07067594d329f95e51600a268edd38dd1452515be3e88dca5bb66c047d1b5c2c1bde7cf0d55915c88d371506df1850c32b6f5cc1d0c0989c94ede260344176633742dc681e2a4aab5f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e9273dfa2891bc0195cf64b0be2fada7617560ce32f83130687a2d8b22e91aad10e806e7bac7084a679a91e261ec5aa98ea41615ae5c0801c5d9237f861108c49cb4bd6739d847b955acba3dc82461beac1e3453971dd0be15db201e5596eb55dcd2bf2315eaea0474dbf2ed208e3912;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he01d0da6aaff32fd8c7ff920a135273c3296864e30afbd151139180b04d9e4e077624ddbe7355ef30cf1d23afc4fec46378ecfc05adb3a957597c3954d29b5554f7f42d8670a2b6bc580cba468f27fb697ca27cfaa5e056343618b45b864a48159622c7f46ae418cdd96511c734e2de5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50de72218552e4cc7d3550988af5540fa45982db03fe6ab3ed4325432680d4ba1af429b15d64981c5d0de67eb4bd06f4b115ff78fe4ecc9e5643fe99b1d8bf79d0dd394d465783e968bcb64e2daf502be7f68f30d1307cfc9148e564665c59c7ffda662e662c26aeec264e3973d9b1623;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a208524b074be67b3b3687f68c53cf720090861392e2ab61daa0b47a1b3786d27fc5411ac87475566102b60e441498fc2382f7642235899035d74a5837b1ae5ba8641016b31fa87cc8b23a47cb1a7505bbde56d65fe00fcd8418e2472b20f14b39e5301f8d76320ce3d45ab947d3c124;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaaf6f5c3f0190e0967826a7d4a398e58c971a6ec8cdda32d52591f66d752fa666ba1cc22228239f9caf65660be956dc628833e905205fffde0bbe9a7406225ae6afb434d75afd0a025c3ee5b9e902293a2cc34ae15c99329d7f20f1800c8bff36d91c79cbbfe28af9b7f989c1e2d9726;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb69481a0fc5aa4a8dcf9a534a85a3497001209b6d5882cd7dd72f66ca672f75ccb1b264462f4603b19cbc84592da15936b93833c4a546f3d030c5a18fb7061ebbf046155fac2bdd89b6759422f44a4a0a2c59f85613a622357b77447a5863ac2248178fb27f1bc1b622171bf0cfebd1ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55db7be559674afcf11087955a3568753c73e6c7968034535558cf9c66ebb4e7a0ca4849ba1a7dee9a5f2c70ba6c9b54d8d81a0a23d35c80b1ccbcbc8d168e365777e50ed5a7fb4c147a234aade18b8047a744aab7fae2432db181deeee5ba6816e3e479550a598b2f55ab18937949ed4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa336a6a43f1bcca175a6ea949a894460776d65dd1284a9ab6c55200e27511ab6068fd14bd0e2acea398d7574ec0f2457df9d05d7435cd09b4984c2760d31cfb6ffdd838f8992ead8ce84b991002d2ee224c0ac0ae4ab4349d7425aa0fc25e8d0841d258c221cd696c61606f081017616;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbbfa3b24fdf37cadda036068583a02cb5ac923c8e678d5fa7cf012601b67e3cfb48aaefcb75fe748b6d0edae80c3351ba0dc378e2f33063fda5a318669f241987d290360252c29fe5de0551bb71ac107ea8310f753fb5a0520c81aac59dd6cf9d2a86e50c0e82d8a2dfe5bdd073c2472;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2808b6e415982bc1bd70340eea2f739aa63eff8a9a80327f13386d4eb18e8ff3e47fc86c59bc105804aa6dda7f1532010234c2fa81c64ee7ab0505d25cd09015ff98d50762bb08b220334979fb3803e7062f151a97cd7f4bd64abfb6ec9b29c11aa02dd90cf50abb78e0865387c217bd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c182a39f26941248d40fcc5f7ed6ae9b7c34956c7660ab1f5ccef9c003575556306c3b687400d4d93f2967a57c4bdcb388263252c2bbe6eaa590bcc5cdf64762b97deeebefc1ef6de70934ccd017a1938f20c03c5248b40230d1acbb5f1f2476a185646fed08468ee83c9914d251ff05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd35dca43482757e4f0e023280ac46f642e388c99d1fcb7c93c3842fdc0f4ac665454f5d9e4045c8340c07bbf5e412601923051c2e1c0e00d288e08a1f542f8b2949fa21a74d491283f06445b8f41e5be6ba6e0039380a5a99db01935406de9163616405b041df764a35817f2fb01cbf3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb58880aeb4d5017d5b760395d8b756627ee5cea9d711e34a74b87114952b0f4d949aa5dcc9835b34ac06e285678ff65db892a9f19caee24f6280a9f5f72c1af7882c2bca9d9889045c75e6a8c306e82b2543dba6bc28a66d69b9dac271a3d7fcda711a44078869ac32d4480f383da677;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aa60b70c59cc0ef6e3011617fe8f6efa2c79ffbe9620176d7f3c93e5399ea58fd153a8adcbbadf6d0d6f37d5cb2939d055d156db136fbefc33d456e6f967cb763b5148ec06e73ae891d33850dbd5a2cb6e7df19b0d066ed0be0dbcc6b92d0913adb742fd3e7aa94765a224d1e298f89b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ebe404c38b777dd72cc16a121c23abbf290f63a378a1f240238406412ca82abe0a443e79298793ec91b122bb8e033cd588c59abc0b37ef9b7af6324d5c49fe7e4e1b2b34d1314be37ba76a6e3470db476131e8e915d893e910d5ef22d9e32846eafc563cdc5dbbe064c91fba05eb41ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2052785e1ac665a9f22105c91b231b0ad735c2846639bdf3197d2793230a4951e09e81764f2a28e108d4cd43fb4cee6e3611c7f3de986f1dc30b1a25297c4e3225b3e81a642e6472003a00370c2d99ca2981a3f8bc3c0c641edbc2f28752adfd563fa7925acfa38c8ed059d38c70caf4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf70ab316b2b65dd3d372449b5bf3cece463be67476cd70a0e05ff6e57ae1411e3bd20f405f5e93ab81673706516cc2150985319989508be3b703048f3fff402f7f32597503f21c91efed75be13e4077158c5a70ce6ec7ee13275240ae8760193f6e953cdb44c830b0924f7329cef1385;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2eba6a3d75625e3e07db9f9f3714ae1c5e43cef0c3aa27e71a3e496c99d843f353e6f10dc6f9b6e0f0ae50eb7a938b786cf7cc74e3c445e91ce85b396c99ba2ddc6886ff8277febbbdcab45de80ab04bb71f6f854fc9cd193f5a024d889d4b00352aa05b8ccd61f1c675421d612d7131;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd95eb6e2388f8e083301f8c96b537c4e194e18f05223eba62757ad5aac11649039824321c76372b6ebeba193c2fbd7415338e16a6fbb60e06fa95fc8bed12c1bb0e87819398aec6cd6b5e53a05301652b7cee0185a653ebab91442c276b537fed4b858b595ccfc6c29ab041953cad6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7e1a2a15021b98b9a8bd9b936163387c05e26e29dca1e381e32d82e136edf80d91c497fb94356d5be2abd73ce77fbc65c4e8dd2f2307b7deec1b1671b88d74a9c030b7eb7e4677224abf5812b07b460afc79b214e370d43ee09d2ee9e27c8ccaf628300b714432de3dc79b94b2726023;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18cf575b5910334bbaa49d1bafd18b74585bf10949433d57000402f49704069f7dd0b0e5760d991873f15d34967072ddf70e1ae4e2efd5821538ea98485de1c704e1272738cbd04adfec08da41c4af5964e0ba0cec462246aaf2234824c16411ac81fa3707f41cdd11d2cde395e5e7a42;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ccdf25748b3ee986bf5437d76123918b853f08973b104e94c733dc8987aca2764d3c424490f4bfa963feca6359f3292f8a4fe1f2749445b48320ead5361280a7a46a3c9d01ebf3d8114c50b3ed158c5fece86e462d188438e4d265c508573a0c003be71fc08ee770bbdc3d5d50ab678c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ef145ef647aafa8daac0d501c2c269c90fbb884ce4104008eb7ac6ac8d8e8698a57a4b62020c4661c8011d535988c71ace398c3bcc3930a5b42f30d5a81b3b130fb28b5498909dd3d85380ae642fe62ce7b46355445b0d2dd31b7181689882a7c4e3b86432373a40d835ceab879b0a76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac7b63b3639382478599481d42ba8a770607a1a38995978072634dd9dd3b54864e8815e67e96175e50e7eb0a156d7537251e7b8d45b66d117395d0f480844b8e7fbfdf3351d9c75d20adce326bc924bd7947090b25eaa61f8acf708cfa58d8d2e33f4121054f82c491850b18bc054cf12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fc2002c72f0c628dcdec1c218bab35483fd642ec5fa91e8f2d82ea891d7767b3e582f4613b81bd84fb37f8306421edeac51ce7e4b9dd76036e5a8747e7fee3ce726a8be3c6c9d1abba651635c377264d6024939404f24560bd7ac0e7b096fc2dcb10064f57bfbeb90d2351a0aa3a9e50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0ac2bc5bd831fa2999f098ed1732349699bf01a0a6f0b0a56095f9e60bdbdcda88ec5627679ed282bb04eba3a0d8b5b292c1543a6a01471e1725a3c6baa906d4f9e9148613a9e3f7c06e31bf083545ee0fa2678ce6fe6e778c303be12164792d3a511932ec2fa5c9eaec798d26b4e8d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2c910e80cdd5a34e0a85b92070f4c929568ce0f98280355d45dd194405f51b9eeb1d6dbd51bc6b37902feafd508c7eda9fdcb193dc28ada4842f28ecbfd8dc3c94ef8bee91ef2437554a1df633078ceaaa6be94ac8e4286d708e27397c8c0db7173f4ea18dcec085a423cdbc7b7f3790;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c320d8ed6ff46dc7be17cd909c9c4c4a15296c4cea989298ce07015659eae211aad7fea365cd80d62d06b2a78255a7b3b5150ee4e7ddd0ec930f6e06d15b630e91442d11097fe785d33759d5eb2cfc56ae2afcaab0bad0907393277948984258905f5fa2f893e209ff5161461366f659;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5593a9bd1e156d2d795c5ca6b538fd5e639f3f5d8cfda22cbbe4fa38d77d9760b8d24a5d50e70b30aa9d9f19422ccad55e10953c759e7c1c9333ad321aa5642e46d45a543b389e6de1460730bf75f5aba40ec7cadff8e90f7defeb71ac4a9e7d9817e3826c7cb9e32a1140ec1ec5a1754;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1f5b9f988b02fdd66b16889b50c56d105ebba966b1028ac2a5c9d86d2b5724e9bc63b5bf7bf97e0d20988059746756490878b05b7e2e32bc3116b91b0b0af286dbd03c24961f5227f52bd61f85da2213cbbfa65eff5ae9524ff3ba57e9b064f5724b78cce4f6d7bd34abac27d05e946b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h280455fb3fb75a896b5ac2628b2db66c19d3e5cb49e81b3115d912089c125f8ae57dea8397be4c9cd1b76c0fc5e00ec528f1c430939cccfaf4b87415006ac0a0c6964ff5c0ec4e9d257d42c564ea5a1d38bce69f4f65c630640e77518af08d845e754bee479b7921b428376de92d8783f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a82332764eb3cf62e30df981321a92d6ce1f3b5e3e35526b0b791a43e8e702c8773842b69add0a6b71e569b6f85dff64cd8accf1b08518f1838d75e471d63640a3a52df838eaea778d8674d6ab254b0dc896415b519b5f7c8bba45489fb0780a94fe54e319802f817debe59721e70180;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h525f42d6d180dc6d27ce0207f6a6b2bb7baf1a98c87dc336540a8585f57b135807e50eca95ed9811709fc51c31b7b40e0c84f38bb71079fc7f26a57e16edb81a5c0205ca9ba1c700aefd178ffe2abc379cb6995d9b302937fe708ba2f7bd9d77d8e2ef375c0f7a89dc9a5f28b5da264bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6f0c61e2391bdab6fa2633589fdab35b46fb4f5ad2bf469298e869addfe7f02045b519bcfdf0902a792e7cfc1e089d4fd65f8244132e485abb11fcb85f2724574a5a4c22c1988ea24de27f27863f743dcc96f7498deaae48e1c44b5f5d626101d728cb2c68c5c2ce5ceaff9e27743986;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc76fa76af893e7f2847eb7ac087d87da29c450d87e300162f14b2d1657171a19f794d05b1b2eed8ac02d1e9a7259662683d87c91f22201a07342d8ed48ad3cf3cccb35820b40a6b9aac66ae79d636da412d86ac70e62d07fbe7377e77a5ec8a637652cb7e70ff33da33bbb2ac161225fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bcc9bf9fc406cf708956dad2d74a9ddff36ddeb2d3166248a087e0aeff964cf5eac6eaa18ba9f17fabdb2d672190d056517aa38e0db628a1b2f49e49a457306075ddd91c53a8aab077f902f00dd1694f51b431fe4f30adc71c5e5143c5ec70e18fe7ea219012538eda67c32ccd43c5d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44d98f637ae14a8f71104bef28f2e030d48155cf170c30f4ffc544201721b25dd2722d5330afcef9e546758f43115811b0d6f35bb1afc65ae9780a687d605f6b3d154dfae00e612cb8e8c5846b38db8a50d6bed23e1960709b0eb8b8756b3ecc9e1fdd40cfd0e13f87422a5b53e40dbe2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed209deb3307d94d2a93e521f1cb939f3e25852d28d86d1fcc0c78ff25152fe4ad9ed065f65301a13a33d360a5c20316c5b9703c266c621fc82a78e5a435cf637b3337ea58b05b7708d1d08e0cecbf794b5809a418bccc56bf3c8bde67abeadfe3eb16e49e7634597a4d635c4b36cc24a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e2e82316c4053f828d31c8e806e63b3d925187bb3abf21271d025af69d16d23206eeb1d647acd970c428e221690f71d064d060818e57ccaa4e0ac278511a35375446f174ec2b23caeac0a6a8e7e5925ca19f22dc74c22d91584f9069ea8d797268f9db4efa4731723958a4a0616b1971;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fae152a53d52098ce5ec1e784cd247c2fb67c2d61da2a8ac638c0e1a7075cb2f19ceca08331b539dba7c66506c599b40ff6683b1fc8cc62c0b611835b8c36e5dffc89f48153127956553655e9b4d33a0951bf7577ba155321def7e21eff10e796c04418eb91902801f7cc23602326cb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcefedc98263e5d951fc7bb422e594ae71827a6fda36e589bfd690afeaebd2f63704e1262f15deb16dabc4319225fa5808d7f8a2d8139b0c4ac7e7e1bcfb8db5c84c7bce17f81bef1831ac7c9d3a587d40b1ed27ec08f4eb6534ca63b98d5ccbe21529f9f5d9ea13286f1a9768f1775563;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd75c5248b20105056307f28363213535ee460587f55c8b7dcec1c3fd82b3d1b24b91457fe5bb933e304baf0a12e3395b0f5d6071cf4440f900c12a43bb42e24101c8f559ac391b62532c8e1c213b6c2ef61740c1cd6cf5746f633af463399d1f6c14bd233bd7fff48b2dc8fa243675924;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c9956f21204b3b7128e54b9607c9fb961e305e7aa756c206837196c86add1f60669f142db6978920170b20cb16cd88e8bffbe61d5dba95277d848ee18eff697436b8ff0268df108c37ec10f79d98a6ba3942895c6ea499f6e38d823bcd7bbb4bc630e7e4583a8307ff55535082a29b3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h455c3dca7bc2c4f4997e9ddb63dbccf1edb703296889d8170319aaf8d743447fdcf67f6047674e25eb34d6cb1b342b2c391a7c2d2478193e6c501e3da428ec549d22aca5cb21ab7008868b9cea15c8e2b0538488a427d24c64d03ae4d85d380441e95878660e1529f8a6fb069b7a6a790;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he432dc93d67fbfddf6e3e4d4ef922d5b6c63328425a984a4c89b8920f41fe1790f3a29e0188122b1dfe1d4f842ccdea770caabc2ea68ab4f5c4ee7095768dca5b3212a33dbe046dc8798345c9eed201d5a912bcd61e3b25372285cd34617233876480d31f02aadf729e9b2f3d0fd7a35a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h654420baa9c0f379899c12206f58e81ae681eadc98f118b9703be0aa19214923a6ef35b983d00ad53743331dc3ecc93814144800e804bd5782a4308eeec3c4bf8596498d7a625b91b697f74bb656f7a7ccb6fc9717cd30e2ba5daf8b2621fc63b5631d5d96910dfcffbdf9b87aa93a9c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d56632027a863f1e13409b7198b5514f16a37acf4657c7c3162069ed63f1c34a3c7608bcebae106528cda01ce4644e7cb7271cf9608673aa8e22ad65e5590e2f7acd75b84ae6795720ff5fb323b58f7b792af8027902f9abf01204f9fe3744e9166ad67fee69b2c8ad87b12684e2a228;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h794f0782617ea9913d9e3be16bc912666fbb1f40955dad584aa2b95c8e3c58ece9bde3088a99d73924501c69f5994e22ba8b6e77d17e31a076747cf5a28ced1eb482f140cc9410e3f4b66d54073a16641c3e2998c10230cbc246e551ade992a8370068ca224cbcaba2250be703af44e70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfa30340b36dd29b0158fc4a9cb1a1cd99954ce33b8f14c95eb304965c523d40d4a6b3c1efe8eb5bcc23a946ccf7d99fdf59dc953cd459f1d7780827dbde87e100be1d193de6ee20da4e411c9c1ba3a884ee035c4394737fc9c628c38ea14e1d4d73f6333695f6e35de099b2d932f8f57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa79fe24e85a9a1cdf72812ff5f22503267d5012b0d4d6789912c3f941505e39306eb5a74c6c63117e25a27b00b7aa37047aafe96e072c6033f35a028db175996679ee656fbb58743736979dba48cd16c95d504c6e571dbb9a6dd34f85cdab6f189292e186e0d5df3bdb568f49318cb61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91ec106f82ddb02fe9851ee469f5e9ca3768cc5f410f5213b8b1c9472710e0f62d03d0836741ff748bc46cc1d761569fc3d986122a0802de5dac2b5a1a147d565bb613be7b422dc061734fe004330973c4db3e99d6b25178debdd04fa8bdb032a756bb4f19d68a9a398ac49bb0249e0a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc4c7ce4982dd0732ad8389500c634464bad5de38e59870ad20deb017575ca9418b37b8a0cbf2b3cbcbbb31d7cbe3dc29b896299a5dff6b55d8ccfb508754263c26a1f753397524f03f299889f7749f5858e4b6a8d1091a4de31b2de2089ced02eece3ee6bae2a0be7c737b1e9fb12211;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7507200ca1b158789976f28a97fcedc1732fd372e02249179db6a473f62a5770f07209011dd8e96d4ce5c6ca6083bdd348dc033cc5c0e40fb787f7c8ccea25f4d304705b7dabd3c62ab06a208a54a5e62985d0ee54990ebbdae5d9db8053f8291a88041ffd11786e7cf126a4a8972acd0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc29f308a58de85025a88a0ef38c4461f484f9710630c0c792c0b442579080240f9dda244f2333c7df06f7ab361b7282afa49f16cbbf65d4864e75c29f76493d4023c8180486d10411b1771ebf55a555f84bb3f5f8a9bd4228f898b3490d823d0edecec15bbbc62a4d7b9698be6dadb64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h645cb5cfdedc24400fd46a2a332876a6ac1a9bdeb194babd16b54b48ea72dbecee50f1b159a14bca3bfa4511892ed9104e7e3dc48a109fa1c43644555eb14390853a25bf9df56604b2ba865e683ae35ceb62f8907f602601a1d85a44b740b6f28ba61eb645c40eda96ac394b92f2175b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd09cb8c587d5276ae10c0603ef7b6a12e02cbc56c58cf428ae9ef35bc17e068ab49d58e08a9b3103efe87484ea828ba9e1b78a4d2c009d9b9e564703502ab54d1d2b45614f4c71fee608eed82f645ec576c493d7ce78ff06c498994d266cc2d714be77e5791bae7aa0ac53fc7301f8051;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h147da74326ae5d6ef210798fece3c28303b742c207ffa893d60fd61c8f9d3d63da2552bfc88b5e2f2ebe3fc2515867c13fc5aa20cda108716c71fd93f34ca5ce3d76eea83147e3a4d7b2382490675dbaffc41301f6949923526d1876653ad154f5fa8fc67668d05d9a1efaa8e5a9f9364;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h536e26acdddce8e0c3f1f97d01b6e3a22ed5ef7c24fa9789d68cb83bc6a923987e4f270361786d300495ba608d55e84a916ad7aa68ebdf683730de546a1b4f1f1545f429303441913420738df0b55068adbbcba50bda8b9b5daf4c983092cc94fdc188392816d5823efad9fb3348c8026;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e0fed057175a5fc42d4405779832b930f7a9ab6f14a01d0fbc23e264db413969b557a8a1c4cab8393f504f237b0b111039c2fed35c43027e9d490066f2d9de2b9d8b80ecb5fec039fac6091ea3ad1ca6e79b9d9641d0484d7475b7e60e33db1f02839414cde01662e1c973350e3a8d77;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3abfbdc61a816018a25584966ced98269e4fcd597ced6e47a1288c4dc8467a7587145a9e4c858748c4eedf8fa6b4f00eaefdb664150797d96c6ce810e32e077b14abb51b544dec123bdcf17c1bc4a6cdbcb4f4295f45c22561fae0f5ef0fe495e0ef592cf964003cd3b20116bcdd8339;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe61c6832be75994b0a31dcaf258f532a02d2c94db1807421e727904f849ebaedd693b809257f7576e917e5150b32a48b1c5848165dd9be49e2bd1ce1ae60c283f2bfeb021083ceb26ffd1239d2c0ace8e57b4eff6a99fc355fbe73f418aa732554734101f59abaa7352d346b01219879;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h913a1d521b9664df498140a01e2980863a3d35a7dfa112f3cea4e219b5c1c46e1e1b249a65a929d487445d90baee4ab260924076af9a1f63ccf1efba181336d44f66ce3f370985ce5443ca860d180eb24410f8e9f9e66c3b80b2b5549f3f43700cec0bed7406af38bad221d948d5c95c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h973718559510044216c3c3bd01de35f8b0d7b6cb4cbe3830824d34000c974823af2c8a158c9af3b6afd8ee6317c8d9f164a094076a0945abceb24d37d386a3f01f7c0de2c5f26afbd409a9d1e4ddca9c1eed53bc227826f0a1edd2700b3f6e7e4b0b20196e093015d5f49a6b3dfe4bac7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf849ca4d04e9dc1521756540c800bc6c5e3a1d252294b08d18f15e6c062b2f0caf545cb92b4c3581df7dba691a24e51d3f032041c096542b0746782cb8d9d93d102668ece1b558fff80a93fdf36dbacbb314001c4e1d2975846d885bb0f775e81b0fe98c8fa95070e69abd76f78d0bcef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3b816c7c2968e59afdc1d145f74328dc824464867672ba643b9e939494fea0286140e53819c3bc4917f777a971c33671c6fffc1cc69ecd2fed6cce543238361587f9000dcaa7d327da718aed5a6e2361766dc0bff70d5204c20ef511d99e21b2ba24b405f66a9c0f2bbf96b4d34fe54b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1eb6f6151c85007744694fcf254413525c27185fd6ed05eb4d8a43c18b5c26690039166b41a35e7a4149e0256ed14748fdf967eb7335ff26ba13d8d2494909e5beaa5a6e0abecc90855617a52b33a76853d2a5b1f2d624b7d8ccb685b31251f336ebc56748a17c735aa89fa10faf16ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fb8529f554625e6c0cf4b90caa316beaeaa9c77e63cf7633c5c871be1a47f5379dba69ceea0645a8fae3df68aebd5116d4ff82e9b9453d926c59c84bdf310b657f2e13989f242061e3a0b2cf18c08ad1f96e1b8933b52eefb48a5f5a772c64b49209da606bb02fd54ea5c27500563f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3ac8b196647301f06220b283c0d4b5cda6bb68525c29f0a0e069a643b04dd9d9629789ebf12b6e6066a89a4903f0ca8ce84c8b5e95c436ee350e77d6c67aa6369902524397719ee3288d7a864d1c99f92cf9f25e59e98da8ba203ae49639ccb3cf87fa67e70223516df858ebac80d551;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75d55e9c53d9a304a9edbb1aa78cf78db8226def452283fcdc115bea55763cb210c413f5f0724d8181481f1d8cc6946066dda69baae5b89ac9b8edfed234fdda2f31496bd67f3f1f759c3bebd58d311d69245ffe49a89c6499f22c70bbafbd7facbc4654c9c2a3234fa8f45c8731791a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e8b09d2efbc89f0550c0947a1995f4d29f162937eff09268aa1f0b083979a7026cc0c2b7532495913959b1484dc75072015705320397f6d823eeb580bc9c6e759941dd182fbe4f0320183a02a04f87356b137e8d63154f684fa79bf7508132bb821f609d5e6b9704a884fb891dc007cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1487c79f5dc34325ac96dd9e5c6080e8cdfb2cbd5e34477c0622eb699f6d3df69045d259faa328fc169efad1cb8a8207ae2758b95c5463db98e4ff0b27b28728d9373cdb977cf36770ae5c05bb531764a7a7865afd692050347fa27038b061e4cf3e183cd7046d0aa9ba05120b59d0b2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf48dc866cf4187db02d2019efdb62a00ebcb0ada9ff4bae8f5d877cb34f60f3bf9d822f1d6e2f666c897bf821f30f085ea247d164b86c282cdb22eadbf14087eaceb5e9585b444150d88387d114d8d2322de0d45e45c9b38412599a3225aa59b3bff24d2e53c26e5a2cc3c0fbb7274210;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf54bbe44d8046042ce26b124c025b734f30d953a60920d7eef780cd20a61b77d67b39f130d9aa0617f151a71cca81b863daf305021f4919a26485ad3fccf7f22ac9ded892f99114ebf1b4dd8d6593bb6e837d68220c5eddab149b92f31aaebcf963592d206ae0c53bebcdbad43a1d6c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60f68b9e7fe965e5f8e9eca0cc8025d1e387b04b9091e6a65845b0935d752d2ce8eb950be48fa7a9e4948f5c87e55d46abe4a1296259fed6fee360f3dfc23415ec70ffbb159dc8d228771c9ddbee4e580c72e4d80d086fd815e03307a7d348fa47eb0eede3f08fc0140d7bde32bcec03d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h484c0ab24ba0050438b13a19e53e7dddc45fbe312201b32823ac4fe89ec1f3a60d0ddb160f19981f655da1da7243729c5a37d3d893f7f08b5495f1a5a8af085244f599a110d171edf28f0ae2330aa5aace62c0ef78b9d0f770ac868a32973cf369cccfe6650052da98c2b34b5f94a5df6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9e7a4f5f4ea2ec6bbbcb101d15d966debb7655a828b423901812f4957b3611664a924f0f870487b421eaf38ab67d718e67f51193c125105863065e66f0de4b79d6c4d6e291f4b13928c251458e703380ee6b0cde58ba6d86854e55c934b7212104db576ccc20bd6f1c0603e87581d1af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39e09e29d4ee7eca9464e6ecf30b76ce370c6153f38d4c2f9c87fd1c5f099eb5851896a993d660d2a81462cdcd55e952380f0835c3e6dc1648e4dea6f5054c54081394410ca350f10f9839b7cd497d67fa595c4517e4834ab4750c44fd1b8031ed1c6546afacc5e8194c74412ef194159;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe66f4293f0233aef6026d72ca08cd389b12d2cc35c5ad96ef60b852ea7db1cf4789c69fb1b782e6283eb15b6b0f162d26b4758fcdec818253e263799445baf79c97903e3bedb807d162e515915b4ad1072d52f7d5eb8c589871e39e224705f01712aa4b96433d81cd602155185aa30c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd82b6469769dff017118fb74b552f84c45c28c8bf3618be7ea2d93078550eb89514aa6179e7842670622a8dc6dd88a08b495fbefe3b75b3bface9ce5799a2a97ae502c5e7f7db19bd565a02d9578ca3c21f4eaa62f7d46994cd40bdfb1e253e682348261e5de2e10382c0554c218d3ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafe5434925ee20b7e9a721987129ffceda8aa73dcc05b4c16f589d345aa5b843496461c912cab1a165261b50ec2b86e2fa5b2d92c3a11cfec1ea19954ca9afbe20130f6afde7698e1c118cfa4731c13a88c1dddfeab64838fcecc01f69c62e43cf9321e0a06edf33c9c454cb6a30bebd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3c32d18b97e3346aaefb7ed30ebfb92ee6a3e56f17b6163ac165920edd1b94437495f5b9841eb8519f526cef6eb37f41db8db222f9f20ad8ead072c62ca4b5d46f2095f4b5da9a4ab15494495ef62103ba46ce88047475a67a5dde41168660cf498ae966729d05211e8ab3d99714b11e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e7a4ee9b25ff8fd1b6d7ebb642ea1d9e6abc6ef279fcb792cb509c4ad8fb5dbcf55900eb83f6417730b9ad4ccf2e9e1c6fea2b4d1623df9bfe43e4f634b9b8df7ff5134a37ba7e41de852c4c7595768c2617755782c714c0067eb23162c7769727944fb176f464d6270a8f7fc18d95ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h574d1fbc1f20d08c3a053bc096b708ca7cd3288f2a908180f7047844629da24feca5819ab0c1d90beb8033593987ca2a57e3c2f80f44f72bf123910208a599001238e8e106a256f25f9860b92c9d497702ce226ffaade0d5372e5326b042bd3ebf4a226ebeade5e416c47730675bed459;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cf516cb50234f052e61b13cc3d2becdbaacde3a79e9f4893289b5356249b34995239384e73751567ca8944454c1bf1f6366df24d505a53586d3cdfc2252550c39bd8824bd0d27fd0bf3e9792ebd214610141a288c180e98f60a6b9be8ac61410781c5878b49e73bd5c5d5ae72caa0d37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b955c7e4167e502d9d71a7a987878d29ecd4d4b613577d745fc06204c2d96e5f28d38449977f52ce026bb84a1862bd1632412eecf192769873487d9682c312efc083df4af495fdea91d898fd2513dff4a3e8c72fd1dd250c486d29d1c32ae0f5294d9f335f6861e1f09625bc4a33bdb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed5f279c7aa97f9d74f48234279ea5a75d032435f0b9de42361019295f2d1f46a8960a5c6d85ae72f3e5894327d61c63c4cd77aeff4bd51c5585a604f2c29743aa94a63bcddfa36a8293245fd13d79c30d86c0367dc7a76bf9f69a3347dca0535ba4427471232191db01e4d1dcbececd0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91599370ec0cee27260300cfdeea78078216df189069069a4eb0950fb1dc74a602e8568fe41adf57958d1d7db2a0a16eeb29254c0792191747bba02d694c6c8bbcab2fbce886ef967059a652a33076dd972e281101186ef8a353b3ffd2f46293c5290ef6a30636a7142258f13434a371c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c76b4c3ff576e24a4844ae95837f67ceaac4993d1e3ad6c28193ff3f0b8e246e2e699705d76464c99f80686b3f67eb11c6d921417a5c13cd0850efa84953ddcddf759ed80129ed7cdeafd666f12027b5f0981d97b5bdc99b7bb30c14763d8c0b3b20364489aa639e34c00ff92138b7ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfb33b1e0847e018000242762b7bc7edcf2f4777e0774d0c1554a5d537056ae58eccdf317b057cf233ced8a8598115d4a6b49445b13284cbc11b753a993b162b5d3bc391f508fe76cfa1f59ee4b7e529c826a3c2ca1806977a26bc3bcc1cd3be8d116659d1fc7d9616ed054ada1b795f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec90cc7ccc611c9bc807fdd78d134beb50126bcdf8304997c5dee7418a9433240f127f323b07c6b1a5c2c895b8c355db8f1ca64d681a72922d6dab481ff2aa13faf70f64ad487c1b5e3e1a708453f7a029162cf450a4f37d55623374926aa6e2176807d34f9f121743b10d1c733835e14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40f83a6ebeebfecba7bb2305d8005212dae431a644ae9ce1626a0b87689f294c5f404e7b19e2baabf26bef2a5a1b5f31f7353c0fe20a78c1674b294326a84c1da7595c7ac67ce723b81ad41a1a8fd1101dfee468711bc9857d7ad28bc7ae8f3ad9cefb6737b5a235001796a5bc9be8087;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80c2c2fcba5a5bd5a4e562eba765f407790e9aa876bdf3a95c37207f1163cf100a131869653392b459e448427b2a04d5c73585e7607d291ac1ce1dc70cc2b991fc0216f59a6161248bc67d06e8196db5b31c777028fab12eddb9473f3b84f5df541ea6985324bc425f3b91b0c8ff77553;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ead57b253d35a5f348441229874396d753c2a41421ce0f2a8077185b752453785720490e7b1d94c30c1b271de862a2bfd76dc2e0e6116128786adcaee3ee63ecc66b287665907f492de588fe8832aaf5096d4ee2f7c3b2fd7f85ff3f2ee7a59d213310b0be9a0f6cd0d50adc4a395856;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee027bc8da2b1b56cee9dd17b22336511c2002ee275a03440859630db1b7fe7115d8e461885c618ba863a89d5ab600d84cd723feb38dfa76684dcd73f1c64fc923db404bdd01a6f123f302ea57b641e9ccc5dee140047a3a91f748b2321438f40e4d9931e5457e001e8e0989950c664da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4aa5ff04323bca4184461ff5f4410572937b8f910f222ff0484947f63f7a6a9367c9bd7027529ec4cec66d0f43d3c9a8a30c164efae80d6148a60fe8e9ae2b1b837f9e8154b235b4fd108b17f426a6cc52b9199f7d27efd4539c3a767e18167ef08c49e409668f3ea9adcd99e9ae02243;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9866c716644c4c9ecf6d82caff29c6c8b90428ebaf278f518f3a74c3c99d5fca4546e8823c1f43f0530c39666226d630b0bcf6bac9549de58cc665633e1a83fc670110d39c9ff5a3da9992b41750ec8d2bd4f1c8c70f8d6c555feacad0f09e6c1ae1b20151412173c9015a22a1849d248;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d55c847d0aed53b8c6bc108487b92f162ed46c9815d8d93a529d3dddfd80182bf895fbff093e85388d585aede7b6bdd41db824066f520146bcc64ac59ce54be9a95466ae2d6381fe056a32733a01052a1bf4802c31df9f90c89b569c01b59bfa216fc2ba224facb62563014734cc17c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h311f10956f2a81707d2c7472b974ca0796594b5af7e2eb9d00ba1c50c9a7fb6eebf199d6f9481e75aaea39174d8c2151a9372e3f926afdd71a52614768f5e48909f0d5db815b40e3e2bfbb85742b72c2ac526002c410303031136b49f389a95991824324020618ff7d0e0c978ee78dd96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f653a65fa46b7905bb13726b01f59df5bdccc7eed3212ea5f11e0a7a5af92fee3791eba47ec5eb490e66bc7daaebc0b5721addc0261e57f9b4c58aa4e0e7840f0d545b55efa8f0abae53d327c61d9eb33f1855922c3168e74eb000692f57e91f9a6ff9469b38294ab3127e8cf8728e9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8253dbf85dd8e80e3534c7dcfa5ac391d4d18691e193809da66a01f6498d3fabe4c075450011f9a526a522810bcdebb092f25a67a981730cc35377d13d871d0db3a868b5b5ef73ba8cd86600ecfc92f2bc091a8754d2a3aeb42e52ae4f84955296a64af00b8e133a55b117da301a51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h353e5663e1c91875413d58ac33f4cb9c045acefcbb354108ad96dcd4437715f7800a91e74670ca0fc5bf67bcfe4b7e5fb14c8a54d51a740dfcc47ba2f7792ba2e902afff2505eaf16b4fabaf3fb118f65243d6b4a9c6afeed5bb6e190a490f8d9f004888fa067a67903d95dc107d1b5a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2992f635b0f63250f73b75d4ad80ae81301f00e6b60999081ae2d90258a76ceb138e86ed59a4b2f15c116184a936132a95bb4ceed7eef0f4802a95311e88c19b7672e97ea8a0687edcdea9dd9fff6a31c8ca95346c6d2628c21e013a7bff85d4d3168253efb60bbe8d34ca44c9de64a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac5114b9839544be36bb4cae6aaf9ada65ef3fea03552311c8e7b533b3a70c0daeb3611d1bd0ed14850686f5532a8a18d1a981a8ebd15681008b53afa240b4d204b3a1ae620447a3bb5e91cd7d9e2babb367238c8196539f73dbdab8de45ccf20520a266973044ae898fcf15ba0013b6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h837b31e10ba16eb9ddece64cd85e1cfcb33939565a1217aea546bc81e031c7ceb6cd94e59512e0184b4b707ddc19f34541f906564dacbb1291a1119cd82d5c29dbef121e49cb8213cd719b3486519ea96d02ed1e4eb026267c4f69b77dbe340fba344a5f8f2253293be42114990188fb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9ed4ebf01b02679ed0b59ddbf22c985a14c9a81582c07acc08e6bf5fc57c9ba99b0a593e773d529b98fbe927d0cc9a3e66f9f22d720e1dd4d3be8ffaf329b7f97429f721c2471f3783be0cc4f98bca51dd855536dfe4e5bc0ea4f8c1162f6b9768c092d1021cf89770d786efffcd4813;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84d830fbccae8084ae0f2f3fb3a5707d940d3c445284e5cc840b11d93fc7501920ca842267c6cff6061f91645dc72a54a76e27cb2f20ce048a026a2e8f5f4a645c9dde67e96e8555ed64253d374d18d7f94ebb112b75c88d530b0872eea7809af4016c77a77f4f0020eea38952702b904;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0de9adeb6de8e4dfb4c3714729117a7e2b45e37a7243d6d5f522fa0a69f51109bad1dfa3336e483621d2ca566ad8828f2437ad907c454b295cf5fff689b58fc29a077533a68e2076b37de93631f3c1d72a3faa50036635d34b79270866ee5a9fdc6c7b423866a84583e5b06033ea1ccd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc28609c306b6891811dac8634a8973d5a2b4412903265d13db264482a9685bd3f1f8a88713620d6ecec708b4e62bb5c3e9f1055b9fc019136af23418b3a717671cb0af7f8d30c505bf03ce4dd3230db626722d0da856d133b387398e3bda3187107b9852665f172f5904b751fbad3f3e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c75b0bc81a04d301e129e8783cd7b8a9ab3d30aff70b506018171a9902114957ed9219dc3bc3104b916277f298a4163669583a5843e385a849cf54187c3dd8f368f541957bda346d26d283b50a15782c049474918597ed4152c60a246101c9838a71c8232d81d31c3d240134c5191f4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cfeea747dd60093c4a5205bbebf49fd9ca7d8934d3c8e69676721949c8163cc35b5df9bb78e67253422978fdc88c53ead7003d4329df0a77c55ed50df7206bd91ccfb02c9da2485e5fc5d58120c29ef8ce39e225cdeb0c050d232904fcfefc3c9a29cf48f5d7735a2fd9cf1985282549;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8b554b26d9d435ed04b76387278ab2dbc261eeca63aa996e582031bf0fcaf535feda3f8e563c312f491e43bd631c5ed7ad942d0d9b083d97f73408cb2185467d0546014afd6de3cd64a1fd22cf0385a78b64a342f300fab51605fd6334789252cea595c6ec3b5810e77ce39c8e95e800;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ae104e441e863a45b7e5b8e8f7912bd8684503b7a9e02cc014e8db4a2a46baf54d76d79596190879eea94880b8fd95bc88b1aca0b2d9b844fd73695458dcb59a625601721e5a3494439ec2b95bf7c4d2a95525673fa98941e451af40629084fe9d3609580563b7cdb6234f3a62db9a54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd866db9931e0ee62cddd8c57d4f31a10536b6f0c49fa5296f13aae77a0397b2f3ed4e8bacc259250aedadee2a7a51734138768d065f163a370607cf774e50b56eed1e60ec1f812d93616044b605ee2a900dd4ceb22aed1038f69fe29b2d6dff9062939f722893125d1c350339e78bb560;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91f3251d40e4f861ead86d4713fa30ed51c60ac6866c92ded43e3e3d9c4e2645e51539bc3134d73b08bf9bc2d8983665fe3b39719ec829b8203bdd24b239f94cd9c562c12c091a98b7aca0342fc07465fbf18ed12402a67abe6ab9f84a09f24bcadab8292bdf44e70252cf92f7a77114;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53cfd019e5b6b3199c73c705650e1e392eb8b07b49ef812e45427d58782ca7cca14306b07ef445cd62a76cd047243d8eed1fe8d59f0d7d518dd9623a3ed9604258e179be329e436faeb709627bdb1c643c7b4e0558844d3618826784fcaddd40e573f646a876833addde75cfa45e129ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8754a239c6147a6da17e16957f04b5fa2b194d8a357d67059b2c1a3a992c88d8dee4fc3e0f7a4f37f49e3c69601c0e5651910e76aaf297b5990870e29577d3568101e0e48c676aae0c1ded336c33bcbdc161b9a80bf771a185ef84bbfcd5ebc877f0d2031eda6ff53c0952b1416f054eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47bf74110ac5aac7fa939ed2c0d0fcb51431dbe61a4cdd6ec965111d3b800448c24280869b069a338db542012a86a5e60d2a7194f512d64c1efc9b0fa9572080d82099eeb903c52d304a63be4b26ab561878910c25fcb76e0412c334e2861ac0bf453860c682bad46c3a586f807a7f89d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd3cba28301bca6a1f683bca17a22856409ef3ef758d9991ac3a7f181ed4803c5658df5c7c2fec728cbdde21d293c149961ef97529cdc009da5907c3f7330137cabcdce94e207de58dac11b8c55142946e597be3c631ca7a7361cf5d2f3306753b37cb2b1273a20032b6cf6a05878514b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22768c5d761388e9c5772476cff9f2c8859ec2a856ebb5e04a10b36dc7f54444c08c630ee2803ff87b988cfaff576e9daa2eaaf7bd4143afe4cc788c7b0816041955d1fcb79f81bc959dff82ab58c4712c51acfa08da28269d6978bb8943c2e5b183c7e80ab4af481c5efec384b828a2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h720a1895a55cfae302b512200aa06fa561151f714b94a2770a65002b5b1009e35043b55dbab461468804e3d39c917f5b5bfcaccdcf95684d52d0761767b27ddbc7d8590a2a7f3f5c4f95fe0e546878392853fe938402fbf4ab0b1db1e079d7336d9a6c9fa51155a26538629789526d9d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3704f35563050d60e85d38cdb3639597cc8f5ae2ce61851d1f53b6b63b60361d1c64f3d706102a840ff79ffbf9991e62cf943dc74bbe6564124f2de58cccd90f49b1223ee41d915f201c801cc8afd1e8f11387932eb01bfd5ac5d9898a45a04225b31328e29f5fc2239ee457ffd1c37c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3485a63b4567ed2517e389691f30ed5f31433cf07421096282e97a72d00c44389a795775f95c5281d38a65b4fa8a8137bcc52967a76efd032a8899329bd2b977aa4a7b04427cc13675550548a70a3dea4abe145a6b5d97b040ba3e2ecdd1f7feaaebaedb6e5b12aae00eda6014ce1fce0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1628d1687a4dd159a60913b04aacb2c0f5c57048c8f4317051a8d6f53ef5d4032b7527464ec5460ca721861cf7130bf371092925cc5092e03716c12127dc6aa923a3f1d6784562f1be6f946cbd789b8fc0c5958683e368ffca221f4b70d0a735e0825ac18c726e6cecd6ab18b6adaf09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd55abe4dc0b9a5a13ccac096e2a5081ec6df0967b325253484fcee469c7223dc95ed909d26d7176c05619f3a27d2c0d06cc663a6d0e7422aa2729d593fc9288302f469bc451593f942538c2da8377ee2af83d2aa55f410b394cbc19f1016a204497a235e482526f80bd49e490126bfa19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5fcfdc2103f00052a46e31d7ded531fca23f5ec59decc65559668b011eed481c1e3f73d7837c38732d4800e59eb9be9c4254cd8a2c0e29259f7aa5dbe615ab5f178732691c88a74fc2be85e0562acee5a2902a306f05d49f65914b75c7a7cebc500d6671d14c3baed847bb8d155743d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c7145840677f0e45848db97230813b3f7787b2071ea315cf96ade92c2acd8734c9c887f94cac7c977b2626f45d22e83861c3f528e9708b0cabeafc63f824789b9083d921ea4a7b26ee7df9e946e7643bf1617396b5b3b213f648c8f7943e5dfb46363c3bf12cecce8828a3a1725bd72b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8004885e22bfe897db8bca1b8219ef9c74a2951f66edcc2331e20056599438ac703c455a30484e0a454fa0f9141ceaf06fb75c5cbced47f68bd305bede6257c44bcdb50b4aad39ac3b95bde44d95a3080d52bba05fcbdb4271a15de9aa204c1af784e92c853c6880873777c4c9f6ba52a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b95c1ec0ee5fb960e481ce9689048ab59e4b52f10abf228d3ab6359c9d45443359a3a03c99024a6b6def3095b196cd14e0da2af0d7c8a1513d9f1dd9a76970b8d8863be2ddedb92de0beac1bcac3008702edc9cabad27c69e86652bf3ab4186254262ec998994c7b6c9da0d4958ae7d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fa679ec5c9e2b3c9e00602dd073ee8d0f72a9ab94fed99ba3230c7cfc4c68be552b709bf8ef6ddf7a90661cc3212ddabdb86a1ff58b4ecfdb893c4c74ccf61030193cea335af665fffd764d89a7a27d0dee4d8d9e6b400038213d50c2643e92c9971c6463ec2935e3567e7a019cff2e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ce131c84ba7c84c49f29853b371821f274274905418fbef3bf582f5556a5931628ea82f85a3c185b9b22f81ab8c69d3bccec164d7af15452d007b94e33678c9fd96e198637a3ced8f30e3b0f9505886b928807a2908fc5eac6562f819f0b0bd0e2b8687c748a5d059c0818d4156be531;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaddab5e2cf0e2d5becbfdfb86f4280cbff584d38480bd2402e2b395eb600b3188bcf3f13e4059bdaf75666412be84a53ffc0ac70bd80338da72fa7973c3072c63ecdbb384ed976ae11a2f47666036be0441cc3f8b4a1a5105e12790ab7bf22eef9be51e3b6e928891fe7539e94c11a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe6109eaae53e89901aa665f582f7da47944b229cab40e6d8cadcfeeb3eaf377e880ddf4d6ddb1e2f458b0e5f23c8229c66c1b19dbcb833f119335e1b3059915e89365ea8d97ad6d7ff0be2ed8cb58fac63bba40afaed80d0d2d651c523dd00af2646fd0b2c9a5fa18cb16a2601635183;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eb477bcbb2f80dc7d6c778f8cfc5b35c2549d47b87862ea08c29f38cabcf8d4687affae3f07c9a531e6575df18bbdf25a105956c795e597ba4ab1692577b04636bf38b091974445f438e0ec21fd9c4f264b4de80d90a067d29c23d5fb8f528ad5f4b59d273218282acd5e0522d666b3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f951ea7ece49c9c34194c59404e7ecc0836e9a0a3c13ea93173735d2f6e68d68b88ad749e4c837fa2d0ac0a52d98e1677fd3a7dfbd3bc52521793fbf247cdd77fdcdebd6a09dc920cedb58600cf815a6ddf9541cdb14afd6a9d54a8941f5fba213ac6f47b64d557657815ceeb3509143;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89e35e68ac0a46ee35c5cc1eeef2be21113a02834640805561501eecbd451cc0de9a049300adeffb9aa9b80f28b1944ce23f611b892c227d92d126bcb4a592dff283f9836ab94aeb73322b155023e22c4946eaa3baac60842e5f6c1d8c30316fc1c4c62e91b7a9d75d555fcf8481e6fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f54bfc04d66639931f5c3260f29401cf30854f3589367431b21d7eb984ba99dddda7b23cb334d10b70eb0352ff77f768ce433afc63df0b2c60cfc2396ca25817b9e16c81e4596a74fc44f61349c6784a0c315cfbb793238b051887494d953c0539fc043f72012ff14a2252e40ef73773;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1add7a4c859b8c1953cdfef2282d78840513c2b7d6b3612c21e9c87a28edcf809009bfe03ac5e01ba9d13102393c5c996779855a3d60c9476c9f7dbbd734206e71f94ad5591b971de2a2a5fd611f696df0bf5ba9d7dfc67eae129df2820947d56431f44849d3e1a27eac99c0e2b13343c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4f68c3dac6987e87667e1fd3d1c41d47bdd8f418f4f8d23abb865eb2dff665ddc76675456e2c5de9a77d17807c2d61055cf251a89219452d10c61b249b88582801d2a70adac4067549e4c996efa29d229a2554bb2f186891ba9a38431b11159d2141075a2f33b9442839c6f710b93f13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcc3224ba36c57f40c70c4bd1df0105952242013fa7730064124b92f7e3ac626db7d1a94936562a848444ac850e03a4b3d4aa8432a7ecdf30acac82464dee4497e898d7f06d5805d77f2ee58418b78f2951d68f322ad1e3822bdcc963bce78290fe741eb12317ab11399d8c2a21865cc1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdae434800664694aaf8c2f3fa32ca9d83cde7901078e9baaead6cff211f9a9a708e63cccb49fea31201f93e9dcbd8dd1a4a7dce60a7dad3dcacfd218002208f425b43383f8603607c32b3a613b05eda2be2efe031bd96b9c28c02f3f6ec39d5e06ccc8ab0a4f858921e1831449c0d2e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h931b5271cb6f73d72cb9070b5fe51ee047922414ce2875c73b139759a20987f1e1e3d72aa5593a075ed1f24840895e9c610bcd454cb5b688414db8046db57d50672d0b2bf1a5786c1f1f5c81a562cb70a074656f0489d274a4c4c237d8b0276b042fc0742797b89ed78198a6b1f15d02d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h527c5742410f93195859bb6bd734c104ad52c584e73d2371a610440e98e1fcea6851513910b3cb8a169c1dbcbbfb1afbe63d65cec3491c3b3210db02b231febb4cecbd25d0f306d54d25a85a52deee0731e2a805497fe06c59f0bb6b3358ea144b83210725c8049f59400ad36a5b81a35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4faaef3c1fbca5b00dd28f7ea7cce6065d964ed09ab663b8a05a1ac7006c4f4351c16a097657806a9503669900b218862d4e9a8e2c306047307171ea4db6f7eca55add5ed1067f2df6986f99cebd21e1dc5c6a679fe509e070b4ca187209faa013855ff7997a625c6c2d5c031c5eefbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h937ed675e32fc6a55fab1ca301754023466681f052194306934fe4ff6ce7c47944583f14f7deb628244f5b4cff20e6dd32acc1e9519804129455afde66b0d2d76a2af2f2085c0b54a7bce3d53ee29b887a70c029636ac772b819e247f9ca9e3e1d121c24450d3735a8afe76c04196f042;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd2aaed7ba1a6d317ef81fb766274102328a944947d0e6c86725174bf8c249d83ff7e88313fbb4b73359f0983e6735af45d588870811b68f3c264dfde5972fea96b6f8198c2e801c8927dca2b6a20c4fc1e9d9a53c224330a205a2cc051e60841fa8ca795413619f0cfbc0f2967b00ede;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ef712b91be23636ab7188ea4aa5814b0aa7d2725ba43b9cb257783e2270240963eb1497ab73fcc56373de43e7cb6987f4fda0a8bc090afc1c9944739508ad2f1eddca024862284005fb87a3b1f371d19863a907d54e4e4e0eaf428878c347dca19a654eb6896d02ceee1f2175a1f308;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf60b403a4a9d8d40e71a52063a37dec80c91c9bd33cc474a9fd4a68a780682cd8f86aad6ba90144ef280c52f2785735daf6b2ebf89ea35b96abb66df1204361c53ef45cc1b10da8730e2700f7608a481e62b8d3f0c45597899732247a6e426bd0060664e57bd20ce33112fd1f6d90b55c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a7c51f16e3a92205790ada442e49ad0f1d60978585a2dd3c294db4c6945b6bb75b32c05012c01c6bbd35d38a0a477ce47fc6274f2bff3a844ee2a092ec3afe9e48ff45ea32909ad0bb17faf0ee0d33b9f50b3cc9eff498e9a8cc2bf9003f410c15f88910a1fbd49fd988a5f8583ccfa1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8b7c3e5ee6688ca81932538e63c6e5000ca6fca05b89aee2707623534b40eb4ca6988a293530d0c23bd63298a1dbd3a0765d5d4378410a825f7662c6c2cb397679f18c719285421b1a544001d85f0940870ba2a85b0e1f61b96c8561d6cb70b6aa126d8f71faaa70f8c8fa72af6a598c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0d1c9a7f8894b37dd7ae5cdfdfd3086c71c6d2e22ce65a87cef21dadda62946cd48f7e52bf1ac64f6c69b1de2d62ee23423ef0b1db7263bcd48f2378b20e6a22c427d2285de6bddfd80a24a2740a32040d3bec2388178126e84e133aeb50b04ad391e2745d0678423e136b421eb7df45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf949d4383b62bc208cb1ce9cdead51ee257bdb377aae6beb3ea19ed0108b97d2c6d47483e9a9f1274ca33aff4e732cbb06079ca76d9ed3e671beb3a3892230e5cec570489b69b957c907a6dff094d703a886a6c98c46994ee4abaaaa5e67b33fcca0fe88c268a06bc66802cdc38664b0e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd26226e46b553cff89c898a0ca852a5c1c043def7e69768d9724f579fbc9b664b5ea560843a7536cf966892d1e1b0da7166f42e98e16103a3c9177bc0e46dbd94e4faeb69a6d5951c66a19f29d4f58df2736191289619969554fbe762dffb9afca73490c9221aa79890e3856f334518b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97aaad947c5f2064f12381c361301cf649d991e627da0b904fac36d2cbfd21a1775d289655e72d87a5f6965b5124c2bf006d0d2f14e1b03cc2653f9e6305c8107905166f5a05482b803945b0c0496789a45cd2b9294b87ac357e25ae316e3ca2f8a29bce2ed818f0ddf3227bba7e223de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1d58f261602fdda1bb80f377eb623a5972cce80578d079c71cc441f15ab4b13fcec62d409d08ef0909c89163e20bd74cb273b3f5345ffaffec0e7b0c2ae77202e5b70acf066732b138fb323ec874b0676600b360dbeedbe1551d90f5e6e6ae7d529b59178208050759ed5e5784ae3cce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he24732ffe5773865ad3d9cb797b0417b1f1041bc9a0dcf2ab6818bee4e7de9b6cd95f322940618a215428b5c6e3a0d4dd1e44d3d97c4934eff6c1312e7314d61d24131fa14dfc0f4e8333b021dc2710560849d55f0b87c142c2c4976dc23cfd0db464e51e912d09147f961caa6cea7a5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h135d5264ae59efd48d21ddd5c5f04c43c7d5bbbf5cfd26eb867899138216351fac81a7cc73be20499c6516f8f173d0a93777d3f0b9af354f5c7812bdf31b752964f821be5f47de7eb1a92db390cae15754f226b3883a52d75c16d952ad090997aff2d749d42f69c2cc02929119fb56fd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d1a21b3f6039157ca93fd56ee0e8c38e3a47f0833da3a33838052d9754f92c10c9e0b79e8b54a32ea1c25700336dcb103de74cc0ddf41d2d8a265ca7ef95c989bcec928790e39eab1a44a9482a830f943cb1b090a05d96f706914dd55297db8768e17635efae4a959ede68b70ebed394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d186c70eeef41b22dbdbef2aa20dd82259a68ebc8ffdebfeb955a02ea684e7a39a49daadf1197ef6133f080f9c98648f911a10ac96980023d8a16a437e451119d7ced122b6e22cedf5f624366252067a7e0c352a188a4808244d36e58ad25a69fbc1f04553802e336c8a5d1ddb89e0d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a20278cbddbc6614989d47f3ea2941c2cc3e90c18761fdb2d14319a887e952a0b3734dd5d89ed95c252f9f3e78b5aa04f6a1b43e69bc1727bd179a4291531d39fa2ce6ec9f73774d373155eca66484ed3724d8b90b78e67865001f5d4032d0962c62b331e480b6f2e0854d86f00d7c54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e9842ea34e3af3427ec8694aa358bf4d5d967f5ca1dbeb2a1d58d85599efb350198c003684d939bd85f9cf711f56e6af9f3b2e9c455ea9c3e450e957580377bb36d5af5ca7694132fcb350a66db83307dbf8f82456129230cfd81b457810efd05c45d0cc3dc00bce01186eb5dcb8ba82;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29a94abc29546c7f1668270c23aa7983255a5d6fcd022efbb4370b39ae55b14c3fe8961af67f88cc0226e6e6455b80353ce73ad7817bd8933984f376df395377ea9cf1d1f3b49d91edd5859835197945fc08298549dfabf00d4fa9431a538a1d43a60728b942f757e3032bfc71f1fe87d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha35d2d0cd0a0b41669c9bb9ca5ad41bcc476209a50a9a852756b8e528ad724d1afb1e5330d7ce3870a1fa800db2847dc69890ebc2eb96e1ecc19ae65d46904fc5ff8892b1b989dc5e64a9d263226f536b981b3375547eca975f90f868c74a4b50b33fb9c89266d98a74a60233c18efe8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha821c33d43345b8f270ac56c0599c9f167a25191420c3d08f39a63262189c55fec9643201d4dcac1bb70dce782e6675e32e0cd5cfb110cfb69cff510abb6f454e5d8078970f8f71ca63832f4897d27e3ebd0111f0d9493a3e2bbadb879e5cd1f0168db753d643e62c8dfb228066d816c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c252b14316aea7d2231688aaeb4c6e281c0fa428a28f7b96c7293df55e2045e546a145b3452ad700c1af855af15ac4ac7a367756728b9f762cb933f9a738d09af11e82219d3bd05eced85e6b007b87866e80c06be19789ec0ff88916517e68ed795e62dba920c95a01d401a690cc6e3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4599260d9755f00c024d6ef1ece0c8eb0317db7d500fea53077d491cdbf630d3c8fff09ed202f2d1499ec84937ac970b1e72ebb2e227f92703d251579689f2f9c225d3b4aa7bd51bf343b65353caa16e784af0f24eb4db569083c0fd33d0e8b209d8a8d21fb483da0b839bd79a2693bb4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacf9d1d18b151d91963107c8555d578f36b972ad855a8101a00abbb388a6dd1fe962b5406ad2405043352073f8eca23832dc71842959780bafa477cb359b3b4f28988503b02cfc09a1cfdf2b7ade1a46b4f74399898ef2d7a331728d12b588b20cd3ab05f5404e17b57764950d5c3c458;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1034f32ba96c68043d1ab15b754877437cd592d06478bff7d6306c1c3ba80195d99ab0dfd40360e316e5c0c9c3f711c35c4fff2571765d4d59e50816a46855e29665c30522c1b488cd98f18ea9238577cb994807ecd23027ea853a88ff436e155d833f7155a97a56d52d8252d2f8c7008;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf37de910888431ddc97d1c3ca6f4d5e875bf8bc5bbead40bb2aeef17aa97c96fbd503b2c5231bea4bfc8ea9fe1dc32bdb01c0600b08d60fec144c03dae2fe52676dffd535cc3bc18f087eb6d14057cecb61539b6f21aa39c544b7623f2abe96b2b26b93a24f06908c5473ada5139614d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc55c866cae67f13dfe29028ece0273d4e202525b9490213a08f3641003183876762e1b1c3ed7caa76463bd513e47c296f8a024668164f908aec869c264b69a6a8c8cfc4b0e9236252ccf547bc6242789b00aae086becd0f8bc4d0dd0e754771fea96b65d4c92c64a24241982817ce4550;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fdd466a9cb3c46875c7689127dec350a5937efa53aa85317b4f768329b70f3ea4129e743961f37ae7b197a120dc3e486695439fc44635bfea81be112285983deca7d5b3f5c8f544a67ef7d8c63337176a9fab49ea2e5825de54fe508edd13ecde857833708888f69ed9a6bd08907e1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h550876d401ac2850506097ecd040dc897180e037f7189027f1deb242c34a8d764b80d578cefcbfd01e923b7307893e8f9c3e5f9f4c7ec35bafb5029669a0afc259774b700970bf60928f4e3dc30095fd20d4fba6ed4d4234532247767edb6c520c9994ae9d821bb2083d636dea0540bc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a5539ad110cb7042d9be2a1bb59cc282ef3e66e6db3de87de480101b79b36b6f6bfa21ff7ab0e0c3818d2ced3cf22f2c22cd17db0be1f175af0fc80c6c4342fd335746cf587b5b049e1be84da06f21faa05e8f2b4a207aafb3e5d679d62ff3599a618863081e8e595d2ce921ae5dfb81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb29f207bbb51fc6ff5d088df8a2e2921f6498abbe61cc1255570c23e5f052bad5071ea4215fb30be1d558c7fc9b4c5b62092023d270b89e5f96982d08bf10fae5e40f589e5acfc520d6a7db9903df3a6e1232b3ca16869ecb6e3f7d9dea53ea3f64fb8003603648f5a430b91585e1881f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0e63ed4d792163ea72f6b5e4078c662ee79340cc5c4a302d1d84374e010afb1c1ef4c0aaeade89f3484d07670d5b447dd3edf616ec330a3e2b5ef755a6d9ab4bd61db9110c616c26c25e6aadae9213a4ed191089cc2910a3037ea69e2e08912d73561b02550ad8c00d5f1ec56402ac08;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h691280854f0cbc37ff792a2aeb886e439ffed1d616832551d94462bb4def503d02bfc0459bc3cfc3541ece23c58023b925dddf8c788d05873c5472cb2f0fef0d38b86bac44728a21c98ac3652f367b30a721e54f9d694d460d0f5bc18529880e99d025d0457aad14758d4eba6579f5a03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec6f0fcd06c9d9dc269a49397bebefba912170f5744a6cd5c758e5a030f0631b605778e445d9a1b6f52f06aedc890d06ed78745392964b842d0f2c1ee089215420eabf56fd793bf769dab0bcb5fb68a2cec2527b6d417ca76dd4d0338c2dc60b3174032cb065af113b711049efa6b30ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc098f780cb4faad38f640f5f91dc9eaaf195b1c3fe8b281499f6ef1ccae30b25ce7e6f9561b0d8bef9d1e94f12f118dd0adbf3e7752903d68b13d8bb762cd93f4304a67b51ab6e253bc0bed81de367da419ef601cecb1833c7cf4a12c9964ddc458209ff1ed4d987da37ef6fc4210f28;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd379f6bac85a4f1c1560d87ff35f500a4d25367664aca496d40e4895daaa6b67d8c7124064a9509b4e916b7c10b99d30717c41c9abce4b351dc6c6f8c3c4f1fe96d25419112a30d7dd26809306959b43c625971aac645c980b058aeb365fb7bb8f70b71a256035232a60049b322cd9e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38f666190099e38485f9afaa33d48837073b1a003ecc93e36a8ce4c1c88f3267cf3a54b6afcb7a0ebefee441c66203961ea3f2c4ecad21880bab397c7d965d9141bd0b0e5ac2c1aba0b43fb57d945819ebef7eb0e167c0a84fb176cefeef86747f9a653bb0691805a8956100146dd7463;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb748cfeb14863a5eeadfc60896456884a91fb69c1fcdd9d99fe029ca578a62ff83259adc7656de1d3e152d833d76d721c6430fcb74bfd5301ece6bb60882e2cad9142e83a797811f4fc33661aa2e6591498565d2132e108cfe69bf8b74a0477a61cbdb46241b48ab243fbdb57f2bd071;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7604e482b99ae6e48e84d93643f07713d40950b825dda2e4c9c2b903b0fb7eeaafbfd4556ed795c26516951d4c88b7a422e99c920b35eb3e2fe49e755624b2127dbfb7dde39dcf73eb8d668e2d63ec63d05055414ca4ab2a7e1a0813a73d4482b7e182ff5096bb5503312078accb7c2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d46ec98699e24d82dc6e77c9b8ae2298386e2df0530730782fd228fc68170f54808cd34670c66e47984ccb33b915023e105b370a931dd11a229b36ca7c2980d5f6707f749cc49519ae58f51edd49d9865e8b1ce933925a09160bac30ad060058ea74114d1bcefc2ad024ed8583ce604c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9e94b0ba46933582036c2e40cac7887ddc49ddc70eb4193b8011c35413eff9e9b24432e274c00d19e54f54984331ba85a4a61ef5953dfe395be976a4f6beefca06b0ba9fe45ebb07e986c3ba447b868cf7fc94577ef57d758c18f13023c964e41aa900543a0138515b24d182393691de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66026cf4d53b3d6b0d20605f93709f9c2cf3d9f2a771188c02df8bf3616ba6fbf8048b8b661c48141cd2070bd778a526f65d2e09301b1a5c93482b0abd4abeb492c96b9897c3a4c6e529252cadfdf6324e991af812b48d16c3fb60d6c2b0bbffff6850e646fbb05c9b43adf7bb2083810;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb893f08fdac76f35cafedaa02f7ce4661d11e6f0ca5738ddfde9688e405f5d3ccf65c311a44ade1f54995801b2f57234511b4b17fb951618d13150893b8a241e58f1888cb988cde0bf0f50fd99adb0c6725522a67870a41595f11b036b93ba356031d092a5e38c7fa6d44ce57900d73a6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda8dea8e785a959831d83d25a08e72d61a2713c4ef26638dbf71de0b947c202d7e38cbd4a70dbe1d221719e17654924c5cf99ae263b7e63e643bf3cdc136447b7e53550b3578a84845d08e888a1c4767cc4a8bfc7a4c62744ac0efae05d1f23c7f7a4a5f3083a5909f4d4bd2fb9b5f6a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9487389321b656ce5d0194188ff9cc214ca5e83f72fa73de3f73f30ea52792bbdc8b87d1ba3e7c52c19ae681c182496775ccca23e0cc99528fadd2a01e1697725f1da5ebda246227210158e01a53321d2e886411bccddacae55e96371a9b2baa8f6b5741e9df8c28e7ff5e7a53b1d4a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0415bd73dcaf25f689804ab51c0c3cdb0ea1231e885ebc43b9baf3d5747375da329b5abe1aada7368f85b24e099fa8bfa2424a8b6d8f52c7a30d87ce925a8a23c4c47aa11eb5c20d5b6c60178c16d02505f6d85e9cc9b382e246708f7835ba7225ee62097d0e64728f13b2fe3212fda0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haab19bcb5a4ba201af71057fcc5a2086ff0831ce7a6f9c8e5379c8370b7002f400b38dba90ff6a4fd978ffe2dffbd2ce542a4d77cd4eea38c17b2863af7d9694e0d06707e3a0071fecc3bc892e49f80bcbf3d03ca4790b4fb23ef53a59be7ee87f4b932e2c4cd5ae3d0f526ef3166e53a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9934fac51a730835fbc754712c77f0ba9559555447ccf0532309f1e7d154405eb59b2dc84139bb6e17ed7c731be019167461b96d0b201eb708e05596be83293f10a0ee5260214a43a75d01bce344ad048eb982af2e66a2bd429436a84d292bdebc9934a2d1641555c91f64bad39f686bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1ce4eb74da0ccd50586ac8a1c9a4b6c2f50650d2f608aeb734d0edf0313b286ced728d7f692ef8b23be778d719537b3d0698c358240a56141807daf45e88ec3ecd75345fe0803d6ac8dc30787bf5c5a0afd87dd69ff5ce9a6155e61418fef8e7f1a63531cde6d4a6a86183a711103526;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he47b00ee8d3889d5073171d03846c2a87c7b5f7b4238022f6320bd39cd57bf4b7172bfb058e4db2ef2ebd6c715a772c39796ed523c2dad982cbb6c0af94fb223c2fab8d34901276f7562fd93ac5b02cadf8ec79fc08e379086fedfa3f30c6cb80dec756298bca34f15e12ee8b54175304;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h724ca2204a88d358935ee7bdfd52b39d1ec60e8586a259bd9e525c518e36860d4b179ad004d9e426c8b6277222dedecc03c11004262bd391ee09c234752efd33420b25fe7f32e56dcb8f007f5684592d38971e7ed2e8e94ac38d8ed223222644971948a4c3c8fa443c51a32d39f246bca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfee16f74a3364a5b7dba3dea9177e688b646dec66d7ae1220cf4370de172feca015065baccd2ec0e1547164ab7db3821eba29e81c8f703774afcd6c2fcb779157f8891cf1f1c8afcd462709a98c45c5875d1d20a6def054d4e514b65b7c28cc0bb56301f00b842c653bb6b65ea474400e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42bb2c8f8fc590f38582c1aabd59575b78e057559810bcaf4a49d0d8d70cc0a7fcef2edfeb760a9cdcebaa7c6134590079900263db8f4d6f27c2585a7cdfd0b26f54ac76e3baee90c2c98370e6774155302dcdb01be1f5a355a70d448dc2e70907cf28cb7687e145300ed11bccd94a4b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d085c7857b8fb4c0c9001ee9ae823ba42e1721fd79831e166930e7a19d975e6607ccb29e33ff29ecbb4ec2cbd16acd6fd75302fb7a50fcfb64b27595f045709def37b28a0917840767b6bcfb510dd2cdc72141d6b03eb460f2532896f5748f097939c58b257d23c53c1c55af2667d2eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd1c2dcb81aa2a8e08c4d6a01337fda444a610cca11331bff1b2b899d25c2d6cbc17e406688f3e0a95b7c83d198579b3bfc1929446b41ddc659c9e2bde1b0e1d4a2c65967c3986553811916c5bc3c6183e1ebf08c82a53dfa4d92ac071df2d123faeaaf04db219d9acd3e55386485182b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he45a1f31a8fe928dd3c786bc1389f3c78325ba2e17c4204d2d895d6eedfbab7fc8e4bcfe950851879a22ec3773cbfe1ffa9ccf389075bfd8205742371dbd234c8b95cb2688688df7b0fc30ce93197d59d1a377a5e4f3f0f91349b358f3963db08ba67a6549767f0db8b7f4b26a5e84074;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38fae1a8449e7a86485033db173acf752f342da27dd7e1898da6e0a8b9be96ce8045e46492a95ad8aac1ef2f85c0fe5ab21477000fbd0d4b84a51e92dc20fd6db7ecde8d2ae16d11ecf85df25b59e1365a371c2c80ffe6189a5579ef4413d045be0f7c66444b9681915bf082b7c3413f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b8425f949b4a5ded5a117e21f39083699336573558d4724e6a28ab7021030d11972626e27139cdc148fbf8aa0337127311b17ba98190501c95ead3a20323f82776f9bc8ac23cb4835a6d3ea3abff8464c72e871a4a847fee7384184e7adfbaa2e29f22f77588a2698f4c631850340ff2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d33c8555f0ef7f271bd86024df2b36ae81bca234ff4b4efb0835d372e24af5263ee349ba7d16fceb3b6a339a01e9fd28ab010e80f21d1de2156dfb1e30408e8a27b70115a068dc0481c4b152d99fc45b177d67ac73d6119deeeb8cf7e249abb6122f9d8b715f46f62f469f0f4495c63c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5da0dd98f72c38c40c879ea63acfd1f9c02b4acdd09fea6c16b261edc3f13e5f482477c18d7a79171d9e5d1f50baf2449b60bdc0a2dc122a5d44b48ebf43996141e35c8e21585818cd3d88ea28e4e8073d7cb8dce3b5c1fa2901c1741e9db1014ebaf234ee1b8c62f44a897071654693;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb1f44592fda76c374da6fb86b428f372c0bb5579c0210ab4f1213530db5ddf3da1704f806f62f1aa4b1c7a0dd122f4025c689fb821e1a0ecda21f4842688e4ec33d2ee7ced0449c86e7ed141f80232a6b73bebc45a00329676b32e85c7fc354f9838aa9b765f9ee012d2f261b11643f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8f7a8840f2f65dafcb5fbc8b49bae4ac4cfeced942d1f0ef476a0c54958e0e49525a040b1e3fce5f172eb53ccf984d539d757c36d86c87e7496067a67dad845c620efbbe1858753fb42b1ca9e2586735f5364a7d48606914cea2e8938e48e72ed70999530d0a891b8aab626fa00cc08;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddf0636a879e276f1491ae69317e1fd364a14228de8df22fba1d2a5fc8ca15df04a35194f720889b3062d2a5ee1886562e3dc33b783dc193f24fca8b51ade3fb302f3a274fde84c3b912fcb5eb1a21f17244f00cf4118fc70fe0787615154c2b92fd881ca0cd32359f43410a19131ba30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd65fedc19b9656d035302e0e5c981c2bc13a80b167bf8b39927166fb50bd689de4e0997a47edfc170dbe685bb25d93919d1911885bc781d2b3d411f70e7abf6576fa88512da2e326aa0103311cc6ed305df7f6a3b154ebd38c12a2862111fc536414c2ed0979ff5cbda7f57363e7b0624;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h458ee86078c1e7c9cb3919deb4c528a74f3a8b8e180fac2fb73e7f21e56d9bae0ed86ddda7b6abc81748cf42f046461564767269ad2df4b1d4e364e0aed1bc03ba422bb45b7f9de49bd77c52af2746949c4cb9a6016a1468e76dca91d750794c9fbcc5c4ffcb7812e47e63c45c306f505;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f90496b62bb3f307c1b5abc0ea70524dbbdd5a27f3bcd7aacc87d332ff736248062f6999d64167e539105b8c957eccbdd03301c78242340dd7973a1db672a8085b6b10986550ab4a24df0b8dcd81273ded9f9c03270bbe2545e194ff4eb6761c5b4854812c47ea661b3ee0528348d5ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haadb84e79f6ae491394cd7eb676e909b602993c7af44ad3c053b8b2a9cb0b9d652d178aa8a90bc6b3b2fdc8033292965fe5d4ca3f930574097ff1cab65c28f4d104ce55eeb04306067b0ea6a7922e654ea64568f7d69929efffa8ed4077fb18e2513973645973062de6e1d3e3b9a01594;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1178973ff8bb6156e1d570a80cbbfbeb6c868027c7ddab326aa88ec91918d20d296f814189ead262112cac17fac00973f191acccfb5f71852fe0434ceec780fd6ee6c534855d0258ece03194f5fc2d20c2618cf533b85f8379d0f7db64a6b0381074f5f8dfa9f02b6efaf51c24a0d8614;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0dfc441c0a28fbb007729ae66efc3ba64b63b4771bb204a93c5d16e66e7a919dcae3f0894a55a4aa409dff04e2a2da387f5105da2982fa6ec7768e8592d6e10fab5a1be99c48571b0b60c2fe77178b7512cc0316f819c7c9cdeae62d3fe7847c9527fc34fa2644ce6127a2a213883b09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h583567e2ac42cbc261b93114d94c7cef09765cb34db95f2ba911f2967f01f6d9b42f385474cee85ff64d39b521221f821c5b245297049f0cd1c27e0f2240e146328870246ecdf1a292f7a975d4ba7fa962bef18a127aa0bb5b45bf76171eb20c7025a1f95cfbbe06ced792b05d308ea7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56341ae9c72c10e90e5609db19ac2f1a20ad9cecc9f9c26c662d22f17880020e6b1583954d55d661d43ba3aaf778c8a4b6921d024db681664136da0e8104db8df3703d5e589bb104c0156cd7a25a2a634e65f6cd71b8b4096dd655bd401e1740a2354d19641a0f9ac80893dec506913bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ad0e1238e58eb14a2146e3fe6f321d231b9a3865fc7b66d003dbd4f0fa1a24d867e1b13ceca225169e561d862a5a70de36eeb2699c1bb9f2fc94eea66328cb595c95af6aa2b6ddfb56392f2efe13753f9c9a5eaa27c06ab89355ffae46381e7e81546ae1dc625d5c305a8ce4a7e1bbe1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc146eeaba1840b2944ef8252185a45ae3641b818b2fcc89de2071864e69fcd9fb0b919395802c4658aa1e1e53b25e3d7561d9d95139483eeb2b9ebf19eb14b8d1e0ac2694a4c68bc151374236e971972628f17fd8415b2c9cbe3306b96cfd9df70558fe5ff4283e4a4d709a365c137bcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81dd75215aad9e1336cf4be2bef87ae8c75626193e0868c7441b0926672111c40a92e268750d1bf3198fbcd8fd041646c2e79bb25261dd0002e608b45dbbee138d7df3b291dfbc238081f533af22563fd9b34fa9c91c4db725357cde03fe5989807d2a2cfe15c391108853cea4b716a3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ea89f98b9ad2733b25586ecf4adf51e441433a3907db0a407d3d5f1a179fe81949fd87bed297a943abf8ea29ae560f8c86207cc4e1e082fcf3354bf3a37397d35060429cead2e423f6eb2283078cdf1a17d36266f36f55fb96a3b99410c1a2974f14b4c72ae7ecc2525232e48bc6a726;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b97254ad2d8e3ca530bb6db8bd15f4bc51e3a99564e5c77793b506720922d8015b321354a83f24a0d45958cbb2a979668dd4a551942592630f92c9977a0408b0fdfacb72d4904025a145672f2f249e00172e044df8f8fd6ed32bc81373a584891373903bb2d51acc5e2bc2024242a105;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c85c70fed589ac8356cd847db125d36197208f8b84336e6bb3c39acf693a9d6d9d248d9e69afcb57c308ad6ebd0f4007c2e4dee08ccd8f564647283b5acc1d835994e5b32ca155f90db80cb3a6d594d84f5604225c9ec956a05c14faa3aa2d8cfcd355d109d9398211d9057568afbdae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h771a1e96a024c01410cd69902f75bbb0853752f0ada6ae05c9f7a937dfaf681d606a2b67037d42b7dbe7079c6ddf7176a6ffd85afe8984349a94aa21e3dbc1639536525b8b4bf2a9c1e3b84b2631f2e60cf691bdf4d0d9701ea9685a856003fde65c6e50438cc9891499728978cc43936;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a103e02e21a7cb3f701fd01088283756467d580dff711b1e2c35ecf24ba2099aad8c2a9285854f6d75425210f39d0a9579900a0403c16cc267323c598ea154eb1fd526f54537f029c01bc9a964aa179f9443f62594e72a67a97af19bad411fadd308ffcc920b777e9126027248a60139;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8166bf120f7a3bfab2538c434166b988404c5a06a392eb7222f5cb25bd8a6329ea1db89a1d8d9dfe17a45b6fd074efa7d5c621f55468026dcd85ee6538e5d0727417fffc8a656b9a51a67f0a263304a212cb84069fa9464d99b4d8fbf6e3272c3ce503a84bc33c6376a18ca08fc03aba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h739cb98c4124d92ca9701cbccfe73a414fa51e437c99f5ec372e22ae828cef3d3974515ccc0dda883011ab5cc37853226f68d25c52a8d44d1d8fc82ba7fe72955b15c9ccfbc83a8197f4f9cf59f75e27045d3e26e8bfa064a0ec8c63b8498a300d07b57088f02bd1739ba4d3ffac84eec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6662becb9521ca9e85fe3fbf2d78a8dae8495ff093ecafc2754615c06839cb29a7c655ba5f5fe52b0a149cb89e43954b31c815dacbe172c7353d5d1697ea94b3c6bf5f3f1da520cf2cc011df09a9722c04916e5319ed84b68ffe1c5432fda5679520a6878b850269b067dd727ea0a602;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h235c3263342660632ac2ae24d90ad65b86b470d0bc6b663074d773a1c314e8e32b97792d5f2f6a53a786891b108a654ece06dd3cfae7c15200d6b51800b6b7e4139e225d56ae1e995c9db43046580e3746713859600522b2be90ff45e03ed250080946bb71fa64ec48d605305226f219d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5425f41dc699a642ae17c0a5cc9169998945d6b4c876e096b21c1352b4c1c7802011efd897d78e68008a72333a7fa588130bb5de3a9fe63666242822334470abd590db927ece8c45eaaf657fe5a95597e58ab32459d919c8bbf6daca22d95c62b6c71aceeca99cfd3e3d6c0db96d6e3a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43c4d8fe54da20446c539d7a012e5f06922b818db4c59a528e6b9bc2e405d35b3b3927ff2c891695bd1a42c5f1f9f8318408a98e7e0ffc8944e09e2ce695c4a78e06a5a3176b796b010c392422820d520dae8fc6038cba96a25d905a89660437f9ccb05ebb20cdad667a6e02af946cceb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc25f72dedd803359adf984b09ab6e1cba5be5fc12dc04596291fa0d2e746b9ff57f2e67367999e8c796ff247b6a691d1d95b125ae34bcc643600ff53d1a8adc074435e40c9b86bd8fd8fc31c820141be805d701817043fc88d0d2d0ca93a2e8249bae46482aa7ec7dd55cae3f97878ebc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50bf693ddfda5e5b4a21cbc00693f0769b4558e4645b804182b23f11e289bd15db3e07cf3bc229679f78334fb76e98f82e550692afe70cf6f2e15275be4fd07c46309af2cfabe163c381803c6a33d3f0380acf64ecb9ceed48730a529d9d26d3c2c3ad1f6ffa153dc8a1e6e049a822616;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e4259ac6eb930c7bc1264be570728d31ae6ebcbb218dbb8989f8f22b451e3873e7fb21528eb4bbbcd8408d0f456cfb30f2eb2bfd1af0bc72501c42a914322b3858df49e833bb34108132da20e01b7967f26a24678b5f0cc7346879e61da525371593206ef40a627c433ea949f82a54d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h683f7475935a4384ce4ada0a0488ea5f168068a1f74f518a84d1e490232d5a4058fb74b5205da510436fcdda55be0ff3c16e209e5bd9d1cbf86894e1e5d8698860bd83c923f84e6ff1b71ea3d25532708f15fca1aa6cc0ad4b0fa0c3d6ea325997a3ab162af7ee694294585878ef5b5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c181093aea2e2e4ed8870306b9500a801bdb34eb51df8e250f5ba0f22fe60df60779ca6b29df1b7bb3be9c2badc7098d705f663e80a1bbfd53cd252ba5f8084bd9c32c6e51b2affbe10d8e9a36bf83659eb999745f07bf4f1eb7928cab1b1ef1058605c6f8146f79aecfac1790e7edf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d1ed2b946a9d54c48b960d092e795f54f60a02c11278d044183e6002b3515013115801aa6357459e252fa674ca27142ec1a28bce55a76b70a61931491df8278277c8a55f1f9e0727bbb78174e87d5097238b2ce05782746e01bdc665fc4e8b615f7f5fec1fc4e4ab7aa9f09d7b866544;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8bd1a3025cb046af554fcbe5d446383e721845c4e2a5eed0f468b946c47dcea1b9c33b9dfe702b87bed01bda67a22ccc249e6a104b508de9fe016b8e15976264937ff8a46425511e970b418e7fb003bd8a6d76f237a0bfb20af12f04217f8e8a008f0977eba743c52c815bfaa7b73833;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d5d9156e7d407ee97d4a7a4fac5c07c460074eebe7831dfd786bf5426b3dc442b60d3819a99f99a99fe0be54e39263dc96b137165a78eda3bfc54e1dfbb17870731dbce0545d7b6758850e43d057f1f965f950360ca5cc6f5422dc69f0c350253e3f69fddcc81dd4856e3522ac03de2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd386d77c160c79beecc46ed40caa019b7101ed15dd5b6ddabe41f7e83ceed7e1ce163a48635ceaee5ad39d6b00ded4e0f0ee5ea6260e940b2aba5e1d0461016995942893d4a1b8b936092448692afebcb859d6756fb50d481a1b7ae608eb726b72f2517166a28e1ec4160d4c197b5ec47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd28498fe1342608be4eb869d5e084d4221af64c9f66d33da036c22e872fd1ac108c8b85966e48e12ed48b079166d8ddd55d768f6db5b8b4ccbdc0aefd3d611c17df707151e3ce4a4cbab64eaf48ceca59ae838fa2b7ca563073b30b1365f96a60eb4fed8a681dd028403f7957c786b89e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c097f65d68864b2d681b887dbaec2f8b0d0111e3c6bd762adfac4b6ad3c73e8c37bbdef7ddf64df3afa890faaf8a072471209ae6c7d702a6f2cc848c3260567031f93b90552c7f80029c9bda4973f687ec6bcb2d7eb5807f51bdb91d6aa19d7651e187f51300b4d9beec5321b7e5939a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1fcc837d2c693dbcaa11d20e975d97e59adf78f44560a7141992827cb3f6067ec2643346f4f577dbe5a1fd957b531dd44b82ee52d65a043f94f1667ef91777a1dd3dee84e886a2c8b2932a300e63fec6f19483cb64aa7be647ecc082ac0039d7f69b633de449f21c04b47bc98e27a579;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebd7251a39efaec46f9ca4eff5b623f69817ed21362d093b36f6a1ca11f188b722eac461277c83752a0e0909b94abf98d2173bc93430cd9c069db20b8f1a25bf482d458a149dc271155388cc666995503ff15374840a627ff6b3b91de1e1184bc23f7fb2d45dae9b66e2a5e4201eeb415;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6da56343469aa1dd0190f2efbf6b55e0693fc40828462f45d7b78a613e91d94705928b5b65fac0aaf62f40438da8306b43e55bdc520ff0e65933267a805f8ce36a1c0ae048434a683adc67cbb1e1e6639bcbf3fb660ab292eead1b3d917a209e1d6c93da7fa894e72e6c09dcdf2eaab2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d19c0405e0180ba286a62a0d6cc360935e4c233ff8d86ff57073c0f721f0203d569996565b8938de39e92b2244faf5659085c762633651e90ab10a10725c448e4bbc74c6ac7d03ee677604037feabc55886f2139c6b5a11b9f47216b4bfaaf9016dfeeb0673b4379dba4b79e7cbefb82;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab07f1cb62e7c7731f5f5e31a431fb65b599c6f6bd28da9edcf475ccb705372b7785d6a577467bf94163e8528e5ae282a66098c79f68b3674b666067256c6792a2d02915f16ff176af140acc9f923ab278f113ef85a79eecb98fd5d5982cb5b3f0dcf814b57c3d252a7a851952d75931;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e5c2a1d2a1741942ed4af5ffd0d6a529fad215ece7badff92a2a0707fbeff0fb2b25706e5f82246d0548cbc5216ab147fb19be4baac6aa81a544b481e54cbb06741be52fd16d1131010d4271b75f47c302b884bf527de56ee07a1175ec7b5d790fa4f1e72fcc7183dd3724bb9e250baf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f45e4fa137b8de53904e199495929da444d716f683bdd88fde9d3dd9738b6919c5830bd193059788ded0130e974419d7d3c432f5ed84c3a4942350ef879a5b253dbbbce79944d6f50152be0cea1fa31792fd5fe8e8f5ef6467b04a9635653cedc9fc43898f8aaf0d8a30710b1b55dab4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2591bf2bf526019929ae60a4b1d6b5d8cd743ac3e3dff8665c7f011e90f9286ae0b165ced66b98970f3fabc6aa97d589a2dee2d1d258205f5fc9782b139bec838c34d5e14c04f4159f767fc245b917aeab1141cfcb6bdde69d83aaaed5822eb4cb653033bc49f622379ce01ebbcba6855;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa72f8a22eefa4c77ee4beff3d25e35136d2458e40bd54059f2a7a99225b0a5da2013882a02a8f72717848d346c7953b70f2e772736c70f96bb7e48279ced26daf23d17b94550851e7e6a3eaa414aef78b3f93a1fa05be3b98316858cd96dc90b84e75c48ca6e9e2976fd80c5e7ebf08a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h836ba3322ae65c7329d8f726c18b543e29cf28efd2c2bea7c2cb0eec01f01f1ebb09f76f3d552cd8c7e6ee04d8bb834ed8af59ad4aa832fc45f5bf4d97a74edf269fe61d5e2f5b5086d6ac89b946642c4242c0fff27b5a8cb66ae9ef904e763191b14ae463507b43cfc4f353686451378;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2226733616fa6329e535f2bbb361d8a99229730a886ad2d72c9f081030105bc4476b16940432201ed1e331ee997040a5c824ad23d8787b647188e525233bad9b14ae81d5ae5b88adc841fa114f0fa151769cd464e1b98c06a16764d76e0c6f232615848672c86a51cf31e80a4419c0432;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5666ddfb2d273b0b6c1ed90b4322b69415463c04ca4fa5162eea95312c7b721c085d442fb2c62d9d7e94ecaef4c6f4acfb97d7b06fb2896ccf4beb4c201a08771fb02a80c75117de391ef4a9b54aa60f2e2dfdaa125aafc541d1cd658012219bbd2799c68402e61ff03fff96981e5508f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h860239d202811dfef56f1d1ab42e86f5ebe1c1565c0637e40874e7ae41214e598cc238569a565de4f9f2755c9ede66364a683e371884e62268569943ed4f8700df09c363b87568d840fa058be852f7a33f193f4f0fb143cd8db4dd5ac6c7c2c40ae918877f0b0579d61938ebc63ae19b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11bda0db8087e01983bf481a7b5dd770b257a35dd6312965192d6b9d223a14019512418bec72f9680da58bc75f7ef2440d7a293a0e26f520a30350c24d41f712312de7fa7e81292faf5ac9349ba5b505bad7d8615e37af1808eb0c201db4ccccee63a30baf6c9225476412d2c29f6de6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93c9144e1bc8ea63fa0a2483a504e35b78addd94faaa1096ccd4046a5e1b3171f31229643e32fa75a3814de98f8b25c8ce3f94ce49348e7db9a764043ac2d27d8ea3b2f88a35e0ab69ec34f0f48a0e1d20e28e26aa6f725859811056c728e4bd6fffd45e995c94edb6f169cef16bee6fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7c1e81c72d95ffb86f279cffb51837c4978f0b75120eaae598a5ec68df9b58a3e27585af7f5dc8a1937580c86e8431b786c9f73e6e672793de64417f8a84c6c632a671e359b11c36227bccf801a28fed2cdbbd562194d35fe928bcd0961f0f36058f081680cbfcf9b04bc6af1f60018c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h268450208cf15dbd6d24e04e81dc63b44a9fed6371ca8b191cb635d6b4de159bbb7eccb2e941f9b91342211ee36e88a1f6a4aaf0dec45904f3f3601a6653e828a4088ac13f5bb555084244e7a06e9eaf100dcf3bb12b995642102cd88db83b9dba6630565baf010988b75dc699c3c6efe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45aa009483562b7323464fe4587df82edfe722aec6a74a8a0c552a2c6720f748319448e18349c9c6d5e014e699638d12950046721d4683bc352b4bbcef03ea033f494233d95911005638b1575fc8cea797be1dbc6cd710c0a6d77a5296526b04213b177320cf3aee2c40c4e75e2ec043e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1c5c0db113ff28388dbf7318678ad922d265d3eb9f92f72c3fa16e0f544e2e149ed48010927a68c73516aaba57d4172b19a9903a4eabe8552ccb8ba46a09b90898bdc19faf8da475ae38cf8475d124c207f778a202b7f299ec821ba0677218376ca5c0eb69f5ce95d7e696e932dd2ec0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ab1da6da60d2d6491f812e06b6635ae534fa871625a2abbbc70864520bae1abee1145e8c2b6ca6d017ba8f23492af57398dc0837c060d6ccb115476f5f868b24973eb21c5ffa786a9b7576c9462e569e0010395888ce473591373656c0cc48a6ed80f85d312734586bb66b245f3a8e44;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6427c4af30bcf7132a03f0eff9efe28addfe836286982a1126feab72fe61a1b7bd171b155f9839bdd975911fd9a232c2eacca6f8c7e31de4bd9a3101de40befb0a3ad50e9c9c2fd7337c43e5dd48f7fec13b94348e7a7893d4f88d7e6f6c806229d753eda72b22d43d7ef509c533b37db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3f800aa678389d48afbc684fd6bfc0dbe7ad3884e083995cad1052511290eb1a9dcf79ccd56040277cd515a43162ce43c2cee6b844efcc189e6937a8f2efbb0574a129ff7911f8bdf64204cfad0e449073ea676cd31961b97e6ae5168cb4fc0c2e56fee576017e3c94727039af2f43cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38159fa894d3482ed3e962cd7983b10f9e62c2d79283160abebb78e728252593c5d1653af71590da9d627afa7f6e6f0ec4b8a2ae45502258c43a2cc5c0a2c65ce67a714add46f9c73272dd66899a080bf8afc21bcdc69f91293dfec60ab75d0be193dcfcc42361b7c0bee5b8af91f7b81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56ad8a5aec39157f336173223a0fd1031c1113a6d195f9214b2298f36e7d4368898918b083c13c3f32850a19eae1056f077113399929b9f0ea5958678c1ede205a439783395e6ed840e55da18cf19903e81140d4bb442167fda70aa84afc30122e385ae420b5c282fc0a6f8d32b8a56a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee698c853d1f49d9dfe52231d9426fca6e8bdacdefd5dc99593ce6fa6bdeeeb951512a518cf97de93ea71f9e9477f2203a8aba31980468ee35b27f56484e09f876773a14f45d7920016f957c250d717b1caa45737ba5ac386007a0f9aeff23e6911d725f843baee482e446742adc0cb15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b536bd5d163b0fd42ec0d9b0cb7f3b1c8d5ddc3d4e19e2b85f89a1e3808e4f3af0b82cff11160bb1ca516f1a3dd44a1ddd372cb0f939a76a370fb11183a958318c91ea245d66e5f576e1e8372c1709c965b44a7c118c64d92c998d235d87b01c1cef5552dc944f7813ab8708793608ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2034b7fdd0c075118ec011be2f4f5be0fa04a3f534b45d377cf9449baec79620aa018e381f332a778659245a9677caaac6655e2d248d192ec6a77fa07d6c6b1533c500695c5f507f9c63631ca6362210b2cc5d63af8c4c6ceec982c2db31fb6861470b525e3a1deebcfef650adbbc894b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb934b31e4c641e149a1e15750006cf5c28ebba69878da14dd54b75934b86b8774b33bd38d5c79805f5998c44ad9617f531731777167b5782eeaec30682886b030ffb0fcbedba4f2c457ef60e013195a13d3eecb817197a77bafcb591a69b0f00db9f7f752d3b4ffad94d24b51d8aeb0ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5dd6832523e8bcb8d4b846b8f3832442612d3767b9b0c4533817ed74f0dbd3c0b289c5274140a503342be3483e601e82b21bca61df3d5bd7fcbc04bbf8b281a6f95a2fb2848441ff331596258a6bb74ea26046319da45308c7f7bcc224b86d6d37893dec9010b3f55dad78473d9f217b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18a365868bd9081e18f10b5075b5352f59b1126b47551f2603ffe702e3c845dab2363f77b0c2ea27f0ac91dcf725aa93882f628d3422610543dba8e0b4ac5c65bb8c7bc6b6567b91f9d6db132b2a5317f72965521f441b94dc9a03c7741015bd4e355f85f5393cea077d8e35b0815545b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15ef71941049d69d62f97b973b98ff9bf0bdf227f97455480d89833c6c7c64bfa98a57027aad3bc0c4c92a40079c88c9ac0217a70a439043c796f80e751a327ad0d47748caf3217877f3ebbc6ab728d607092bd2afba0e54ea1c16ea79ca659fc6c075939075b3a1c371d7c1265e3e77c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd38d03d26d2fae6f24fb300a53d9c00d3748457286dec7fc0e20f8a9438fb2791178151842ad576f324be3ac9869a28960308a0718ed43f3194e8b108ba139a01cd2c4522a83b5ada01daeec0240d695fafe7e118e50eac999cd5c509f9f6cd2c26f1121df30978a17b17804611687a4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44e57a437a85736444e6edae8dea78342c233135212b0638b0129d54a1406d8406a149658861e4e7158eb34aec77d15881abf9a4b3b410e7ab398f99959d4ceea9960e2b60ffca94f4cb839955530db4e699090c690daff741d65791b36bde611184ec104abd81dac66f9d55febce0447;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d094ed473654198c42a196dde71f6ac2e53121e8c332f66cbbccfff018e225ff17a23a4625e41bb6eead3701b2ae1472e4d06e6ffdd8f471238f7b43f52382cb6525250d5eee018f30654a3fa0a085a652d3d5ff876fb3db0ab50d4336842ec29731bf9307045da5196234323ef40fb6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8870c19aff72662d838cc7938ecbbc4b114342ae6d27123bbcf6441b2f90f1e06985477bbe72c34229a2adfc4fed58609d93f68206e0068e2778179038b603494b2eb38d19f66ce0a95fbce801d30207c6cecac2a5f6d209a2f347f6ed68e0d6bb1e0f9c89a5d1df879121a6a5355f9bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f58e86da9fcdef2744cb8657b789a9b470e9d8bbc6fdc40174cab66acc6978af46766a3d0fe0805555693266f0af9e6dfee51b3ccd1efb4157e537ec3bec6d4b551122d58de4b791d199b699154ce9299eb170db5d5452137eede2ec454837add2b19d5f3d3173b5951b1373979a4795;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40de810925cf182a91928f834dc7726257b02dbe042d8dc33c11d13c0e146aca40672ccb26d611cf87b510211d7444397963434d590f9bad440033bdb24e42272f892b7637fca6dadf9977db1fe32ca80677d19458ab5f3dd85cf8d0b04e5359433e98eb26662e2c96ea333264c2812ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h616cc5255358ae94e3fe6af136d4aecb3a723c5e95154ffdef53964d02de4fe7b1c16bc872edeac9b2559d7696fd37fdc35185e90ad10bc175e2792b4ed98eb606299e376e96270dc7707a7ee09c3cea2db6ffb155bd60bb1bfa6f53be017ebb4ae88ed766910fe6c1a7be00ee394ab89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he46b4e8b82217564921098f186c8e1c9ae1b51d29f5b86a8db05824c3590fe6b9f05d73a9659be1f7219d621e7191274ad9178f9cae10fdddfaad6eb76c00227f273386336fb704b101ae6edfad51d7b78f0ac368a36d243fb9f407d5b0b32ad657999e987a6882fa0bb73f73366c09ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb28a32bc0ff5d63efbf85bbcff6a9f677bebfc4c7934f6cc4f37765af5d86261d216f295e4a72e74452aec0e6f67b8d4acd09300cb2261ee64d64c1d402a1bfdd0bb974b90dba234c561d28dcf25eb1bd5209acbea3454bb33074ddf9c91402c37a10adf56bc0a1957128373eb450d2ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61398d39bb1e5b119dfd7e44ce6f034cf6e8103964d49fa820f73ea647e6f046335b95983cc33de2f974584c6310691b8911dd10b4a86e06bc147efa955120825ce1b32725d0f320bf264ee3ea41be65137af33b664abcd6f2d060093681c109a0fc0ec0a20040255534b4743ce4b3ad5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a1627f65cce3bb8d8725c9e23d26a8699ed9d680b6083a63b7883f958c0559b150df64d46f6ec274bd3a7a87e8a4f74860eb541c927f2fa3c2e7f685fb76eb40e36c23ccf6b5e58d537dc69ae99bbb3ac6f769e5328eddb51c7a73ae4f564a2130a1c825d9dbfd6c7889508931b457be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aed602bc782872654d8b9cfaf0ca9fae347db4463e71dee9aafb767e1e40cb362df3a61f8710c40048ec098a700a305321b87cca80f0d9621d6afddad6df285a58b3ad6b2cdbbd54d8184ba4264ec632ad8b0288d7d3af8d0810f9a4b600ad8aa9c1ca177829ccfd29ea29c2ffaf4c63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cb30d9afdfc877ee9d452eab4a2ec89ffcaf1bf800a81685fbdcf2aa53059ca64c80268abc32785cd4a885d2d6798e973e60ea18ea4d3b531e05b48c78823f1fa5deb79719f555df0e5e5162bf063206fcdc454bda6986d3e98965ace19c1916b2e4daa367123deced916f626330d2ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e67fe41c04bc63986b1ea47ac2667e7cb01042a2f504b5a47cafbd83c1790807f81a01e4547c214de3bdd7e7cf99eb60c12f20247b29e4932951e5ed79e25e177e30ac3986e7ffc6761ff2c626ec73110c9c805f369504108b0892e0814684a1c617333c558b85ea90c52d11b62a7935;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65cd9c75f44646a2f693b61868d9c745b5b40a37cfc2ae1f524e1281dc1930d8a1e270f92851b197155738d24bda9ac90ea2b6c9a80053331ec37b96f62afbd6c0091bb3befe7c85611f77470e6b9d841f15b2559f20b8ff05ad20c166c1eea0b964a943642aa7bbb49a9dd6c7638e3b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8745d4439452d0742bce5e541053e4f59c195af5008daedf05a9bf6bb389234bf7390ce487a0235ce29bcfe674bdcb92fb9266e8223e3a65378846a294fe01021c4690b3c697ca75b05f36fe0ddeefdb0909b0dd3c83c434b704779232bff1fd791b74ca3474ca6720ea26c6ff6417c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h562be958de98c12a733c3eb5a91a6f3b758e950a385a9a5998a5c7b64096229061b3291f1190f20fd52ea6f60d237c0a095655afb2b3b198b1357557124a7eba2550dd55c634395a510eff302d23e59d269720e66392d59e45ee0ab52fe8750156e5fc98f108869c89c8ff837e7f7ef11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcdafb04b629a6c9aad0113ddd624bdd3333263c857b6b43c98ab6ec2779cb5ed0cfd77e8c7b832d15cd5bef8663da0a0e2d3acb49cd2e2f014f3b2e0d7e234cfad937aee65410f23115421a7c97c683fd06af15e3cdf17209fdd92eddd0534c420b010cd81cf189a2abfd8011e6946a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9d3d3d7cd6022ce344df7377569aba2db12a4b40f1e5ccac79888055d0ad432c0bb21cf0c1189b2132a5589c932b0891fbe639e15b3a071424da9fa8fde6d1f36a1d525c067acebf22dd75c122538076045a561ac945b4d9d443df744589149d4a1ad36b4ac129531697cfef94962293;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78735c44cc274c03a85c57ca55a5a0907bc33770d0c722bf0c7fcf0f43bb057884b5bf2f50a1ff9fa4589ec850b8fdcb713dce9986cef904ed0616f0a9af58130aa7d43b834225fb3c8482366b860a09a64143ed59099ca585d8932eb88354de9ed1cda1c919d642d783bf6983569568;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h745d4b8e7d361872ed9c2875a87cc64b6a83a83f84e25ffee1f75404d92392b7a57c836a51cf83c269290be954694fc8e4a1f73e7d4424820f1de0157cf6685872ec8d2df8d210db19ef6ab77439f8b9939930d0b122f35e9bf76455fd7a592fb73b9b5318d0a804d470db449b421368a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16dbf20cb50f5bda8c01aa2a6be93ca6434fa99608813fef69856d6448126aba1abbe864b2e7a888dca169a0ed5f7bfa78930859a0518c114b1deb92573aafd09e9f9a72ea345100d1da8a05f9112b980c30957e764abd861e0d9a8b742c2d21541430836ce938a240d35c0be6fb2faf9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda6ba6f03301984cf581bf2b187ce61781417c8e940727275e54bf96b94879b5c2e0a1c8d11f2a7d9dd0e60ec26098848ccc1c1f92cdbc795513e3ced42b97f23b373efb0ab416ade17d7a7eaa70000f0fcf1a69b9c3b209e4242f17cb5647417cc7ff7352cb22bf210fc04645fc230f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7afa5e0f1ea01b19df9f8aff431ae9172f13a2116cb2c362fb6f1f114a77d47a3da0c8c3cbed9faf45091a81e7d74ef112b66aa99d9d83616cb4a8c84b143147cdc0ada5dd12bb2f4075c7f521c0fb57a8241d8f00e573a48813b316969878f8e92f78addd37900ed32e4fae0abefa5d4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f941e7e454185d030d49d027993ba9e8abaaee34ff9e2a1393509201b47b8d7c8484cbc099920ea72f56c5b769d0d5d9beb20504303ef9783f76ed1b3ac70ee9e7cdf2642ca111ade2ccc868bbb16eeb7015bbcf1572336703cef3f6af548911ab1e7060815d7bc2c9dd4c38f9a5a303;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf97236b64cdef682d6eb9cea7e908bfcbe30c2e7b07130f506ce654473235e2af7586b3e5ef516f087bfe03745f1b63a3ac2fb57d87c7400a420fc8b9e13c4b9c7702b2782b1136475f911c90f601da97ef3a049454a9f843953b5dbd8d1b77e4b9f7d82f2605f280ef8efcb7ac9eb9be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d71fe5405f2e09a7b9b1911191e3604f1e039baf2957729807343230ec7f66de1253e37ac8952ccac11ae2626965b93f0b2ccddf46ea14daa9f0e80baae831030d8ba44518f50d98c68196e0026c09796d61538b158e2358ad985b21d464e77c7cdbedc57357e9e19ca1765fbff40906;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0d6019abe159b834813fb9769647bfe5bd9e2732a5bf99507b4f4b384d5b09ea70658dc07e993b72c104d76046bc117121186c3cc6f617f5da522b8556632a9c9844b7f8fd1976a03c8b72bee131078eb435cf20a8395704114b4d3bb6892a44f01e0414f905b67ecc1867bf09cb9e1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6766789bf655d6bd799a043bfdb90ae4f7961540f697a479ef651d870a7a78ab3dc0c5592d892a6e14039bcdf47228a01112ddec3b94d242048024f9027371d3c9801e4cff88dd38d3faf4b0b05ebedd30afc4cc57e03d927f62b28dd26862dfbdda59cff0ddc7fa068f11b0b6ced3880;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29a95207161aa8719e87514220a2a47d1a5331a86202f2bd16f4ef77176410288ba4935060a3544956f163807a05081e3f61e9188f9472e23b0a629cf8177a69dfadbf7964a6de866e86dbd31112107e68d9bd81924125b6f6544a3d759c7163c93eb982d9906d0065a93dcc904209def;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h794283ad0cb7434fef7ba0d6184172b3b0a69ac9618d0ac9387d113b33a477a9fd91de422414e624a4fd1843ce759879e4732a8966c71dc588c98e61bee7c9593b6ce9ed501d903b31b0d4f68558f5c9c588bb2f21828efe831e73cd3dc52dfeadfab92933e0dc570c6c746ed6cd54e93;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52a948b99c89146b45e7765bacaa9434ba969f5f93d442597614b7c0027bb59790a94accb759c86053e6670964eaff099500d41d3aafec0785055fce08fa65c1a0142c0b217ae3005d1a07272109dbd64c1c45a9680a5740b7b5b03f64c91bcb0ef67976b0e5510dc6de36c407a222af1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he557f4c42c1b77b8cef1744e1df2c8f10a2b294589830cdb804e0e8e7ce2c603b2bac3d9cb529dc3d874f92fe4ced472692f5b052da2a0b0b410905d739e1f777a6069216b62b621a21caddb4c72c5046a18d433192e003fbf64d00465c3a9fa0fdbccdc04994e4bf3ea541de64385b18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61db904d52fa1b011dba1286b2a92d4c6e9e3e4f7fe0219b6d776864e54d9bcff3c0a53c333423d8cf4aeb2d12f75a5ec666abed65684642308335be364c92098187277144b475b6055ea07d71569f876583bb365e61a96180c4d68a8ddabfcef930c95091a70221c8330edc913b4dc66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9c227a7617e09f807e4b8dfc16a64a6ac66727fa100b5d979ebb7a2b6e9932cb7e5b4ebce3632e95b71c837c9a76cf2a8b51f729ea2bd313ef72e9d7b45fe654747ecced6349a559ce57f8282412dd5a518ea2967235b8b138cc5bf34fb7ab4ad6bfe491cb31b51456ecf4613bc5eede;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ebcb238db8dd8a018d2b1a0991b7ecc032c4a78e9ab55c3c059e42068d05666a6402362cd8c4d1cd49911ef7891bfda75778530a64fb43ac11f89c22d12766f89204001aa0b0436a2575a01a0964ec3f4d03899ac845a6933f6d91462c1bee072df2b971edddd515c20e8094d19591e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc35d8db0df9b354deb03e3c2a5a1ecb158cba0f1ef843bd659ccb3090b910111adfaec963c557d9e0ba60325d9ecf928c82f230aa7c41f18aab03c79e6569da297fe06e6812b8c3a05cb222370567c1839d48a3ee70b454febad17f61e1ec1cf07c7ac8e1793299094397ad91879b1045;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95ac0306eb5f9fd3716caa4c117aff17290e0eb72ad3a0a80107675e599eecb92750c0136da6571242b7b173cf3ac65975ca8f4c6288309d39da37e5ca5e09309e1b361844c568d978d866523545671709e432662c0fbd79e79fe055d2c08f53e387aa5364304534feb2f74b53ff91b0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54e229e4d3e6bc9de02478e51919c08da761384c54e6ab919066f0acb612dec5c128006680ef08d41ee2c2d4d3bffdfbf1a5baf6d990ba077f0157d62f31aa6fd4887764d5332fda9cc0ed22a4aae978db3e84d918f3bad43d296085f48c8f3dd939004c5f4cdbfe379b1b88f076fdacb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ae9e9ca4231c2f83a23e7ec218a760f895314b5ff63a0494c3175768e6e702d044a6c5069518264c4a92a9182136f6301e201eca41a03957a5e53960d40532ee84b74892eb438fd8211c17dcc6dcc67eef84691a1653cf749b161372aeb93c0a69dc7507a4466da64f369820dbd9749d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c7e4cb16e44762cf201837c1776add643e3164e3cd24a88e359123bfdf7313a7053a8a01bc1fc8780a85c4f3c9258890f9160d2595ce150413488711319f7ffed6f321577029ff67dd3cb18c9826766ca203e0f856bb7eb80cb6574ec7da2962f53a08ac2f1a5613c5fda2224e609a04;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf269345978697c4811999ac2359d0e6f6cffda0517322755f0cf6add64e75134e54cb6ac22f46bdc4ce6c708fb445cb9ab31157ad1d79c656678df256a0c482ab17a3693719e1f4516ef44f978f8df04f000c3375032d63b78d20886fb2e743a78e9baec8f87e42e1dc6baa4b3f238062;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e22a8d6d0c5b11a71d2f59dccf837460d75eaae98dc9044da82651ade9bbc780725c75a31e400f27d6452c7091d679a98b4aaa1ce89addc8e5473aa437f10abb70b6baab078cf35d8ef71c536455bc9e637ed156752d88bf1d71b72181d381b1a68c0ab832b323dc43131ce5c0fe613f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h493b79a1cd612784690f8f7b803704f59a9d7d264c189646590d0ba7d52fd592d22caed53bb66558128e3a7b958a691c0041200652b946362d0c790c333d0780d264dab5793377e4e3e2aa77f56a501e02536d966e1bc72d784f79da741c70ad8e9deb25e782cae5a3a86dedf6b5be21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5713663a80d084ca0f87862b246150ecbde0e60cccb952f5e3b6084d80fde90658f6b5f7fb915373e1d85e402646b3acb80dfe6c6a2dd178484b9deb40e6ccfad86c309baebd1f2915d2b821342acf2e40c8bc14cfe4c01b0c8a4ca224ac1f8eba42ed88e44d1272876bd9082852cfb9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfc3395751d502b4b5375720de1654eb66f0935561d755ed7afeb7ef9d7f345f3bc0e915ae952bc6f81836d36f7ea9e723a377ecf04ae9ec302b5ec5f1dec139205727e0e12088bf096b8eeefd4c111d4e4582f767f369043dbb15ba38ca12846f5b117da961f09d334bfd90ce6034a65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61ffe3e8f349d6394ab0bc1c4c4c30960a87fc39333c78ec96fdf282bec6c17a779d845efbafd5826a2cfba68f51cd9874bd6c6d549ad6407ea08b8bc03ff7e096175ef3f12023d7ecf2eacb75e62569aa307f531e7030df9c68cf560a2c25bc26e8a21dfa07a88d73a5fbd4d8129dcb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h608e4f95e4b147ed108cae996963becfaf5290222ede7c4316376311507f782471371a60fcc091534d8c30884222f9890563b6cb875aa56ef87615175d710dead29b678dcf4fbffd01caf3f2c85229faf9dc17061d29b9616ae8fb59d76f724927f8ecd4219dd36041ad390644442d7ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb349e86a9ef1b5641172ea6d6c8f955d99577e5423f11673712f28f77742300fe1c07b893554c15c9a8ea9aaa2657aaa706d5f3a4870680742b798249997ec20bb6f6c8f0a9d988990a9966e0406d7112e7d2463d821edcb785f199d500468f939d7b0d18b013ccd9888f087bb06af37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b35faa2dc27cc6fca58cd116d69d098fb169db84fe9b3a431d18d37cf18bf5c2f360c66e27258a939f7cd2c4940448913b6f2ebdf68c727020c80a35f2aa52bc60697d1e0e65b78be5ee5e0fbcfc1d846e287ac97d966e3e59236e2c05ea9c01309aa956d6073c3dfab12ee19ef127e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2f3b0ce95baa4eb6682da04a206b8840bd61ea008073967b67035632f669aa4c2b6251dabd6ac036c3ac6d09e988e9036c913dfbb21fc61ba56ae88281a383364165f17389369d204f492b12d3634be3f2a8a5074a409754aa7695529a957b7abd0d4aa27b86385ff802f3f08174c47a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a4e334a68864b7d2eecd25b9b8bc3b8476a04b02eb1f78bd87cee7f9701c7fc72dfc1c67e8d2d0382a182c2f20d86dbc12e35fd90c781f4b6f487583e8db283ee3afb9d1d197479c3bb199e608c0df90b1ba883abec91a6477cfaabbdd33fcb93943ff72096ee090bc6f2b18aab55008;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd22fd1e76afa6e61642ddc19b37e896bb0474b2ca31cec7758828df0334d18aca0ef6445970893ae6b0f1c1c727c994ec10b789032a6db6c45883f1e829d38472f73af1251356d4d3b4713736a4876b6db648c112f98525ff66ab719f2dd1b1ffd8dfa8362a55f7e89d61faa86d6c99f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83719763db6de90e54f35aa5567cd9af2b7098d95d98a657d67cd19834d90fa1284c1699c12c53805f2090f1690dd4fccc9b981349b964408ebef55cbaa62709b9374b9e0cdc3d12c99da202cea3a8654f15e1e541b8f22b60e9e6fb470c91052975fc006c3f790455990a8b1378cd26d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a0b724f9828537b1d816e6db9a9519152896c4572a662fb41034ccffbce53e87f14354de94fbce6c45e48a4fc20478994549a52459d2d48cb87cae10d06ff365994c300a3f4c2d1c4643942db1cc12545fdb2c638d670793e4a6a2ccc4402c3c2d47d853e701e2614b2dcd80cff80c98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd910b88c171a6e7b6e5a48eae2fed8a317ec802a44eb80a13dd404c4095f18b7539ebd00c6c4b96f51414686657c9dd4dc98e53dbd78d95c78cd62882f0fe2f50c94d19e3b5b899fd0c0a82382e66a8cca0f990526a1091e34ef19a1350abca1554fa3ede953c1125abf470ebbbdf9529;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2579b0a850671864347e9dfdc6253ed91b17429118bcbe2c788eb71aed1b2f9b73f492f999741f75ef473ccfb9b5a36eae25002d6b2c1b6af4c6cccefd8a0c000e81a07c749984dc28f7a7a847e801fb88f1bb38f1cd936e09c731479b2df3259b2b3178ca9289fb9324df36f28c2d2fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d44e3915e0dcd3c1756739e901a64d4a1c78283480c92d874e95a3390e8cf189a96815ee25e3fd98f69e6be2ef8c93fb7196c079730672f763a30cede48e0dfd0092121f63f9d8c974b775eb6cb9cf9333a72fcf4d5fff0faa3e0fc53eaa8243aaca2fa5cc308164586c6cbb1fcb59e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1896774cbce48f786e9cdc5dc9ba128166a09ed497630be6bac00985866e5ff534c43cd96ff9bacd36882d280e758efc705dd7c56f9f3ed9afdf2161d1edd02ca4619d294a93bb0d3f39223d0a2bd2b47756a838b399b6896bdd967ef016ffb62c790d0f11649c6ef3d621c68125d399d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4eb0f02bcf5326993bf99ef25a5bf2a3521628942bbd35f9f47552a2b099de09783e88d569310c946b0ca23f5bfd71f776ddb0a82ff220da3a8a3a322c1e7324cbd2dc938cff3d0d3b655b501e025fa3a4ab0fceb67d2a73b64a5fc2e2a0268eac92dbe100143b20590e52bf626cbda25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82712682d27a33de64ec078a45a83ee55fc3f0ac3fab1d0f9ed6a7ebfd4d66e355cfdc8fbea988e55a204421ce63772ba93fd625ff2d7d97a43924c2e48f018d6bb50fa41d99a03a071a605b1fc0c68fa62465032c5c95bbd63c01e8041349bf1a5c9387b6ba71386710ad6e12a642648;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8589cd70ed55fa00e9653434c1c948617cae152fb034fd355047c5902621f2d68581041a96653646ca12998aecdea7463882cd2d5e0b0a4992ff72feec4bc08a8c108134e4cbcba20a6241546d38329bc49005b468d5edb0524e32920cc448e4ee16d0881c6ce0fd34a0a1add4628ebe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h551eef562ab7dd9c8c893031b67226c66b1e3d13cc8e6959fd03ee566d65ec30e4706e9167a1ad98ac9c9af84a523b7d94bc514d722f380804d16a85a04e7a78b9b8a5ff90e0a1378384d06341b0c99a59e787238ee1563b42faa19a9d922d166f19c0b1b155a8017e316e8c5cff55332;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f43000accf0ce875774d07ba8502a14e340e86c1e89839877aab81db1bd7edbda1df0771141bc284869997f0a7032e237787a2796c31bc5a96fd6f21be6aee0139bbc3809253bb71f8150398981df604127c882de398bc8296bd85af05163124c53a6070a445e092b5ac167d7d9b33b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673a90b55cb47505203a4f6222f3c60c0051b3f7b690c3685969e71da99f5b134465419fdf832d33c8addfd37cafb0ae1eeffacce2b636fc55a809a6be70e21f5afdca8056521c5d1f3be7ca02009a68c9de843919bad7e7cdc075a65773389b634f78a7f46685118b5ea1a6ea8466d61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40b60bea43155c8b548f338de4cc872b2fea808778f2787ef9ed782dee4015fefe6ecdee327cfe1b22abb763da65bf45deac94ca1e00daa33d9ac16f234b10bf5b9b72c77de2ed98fce3f2e613f25d30d3e7b697227c6fcb1667141273fbab535dc6ba051380d5211ce0316c830ada7d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11595638ec44f105994f58cde0a4f5f3f0d208b5e8445ceb6689ce56f10c0503bea60cdacc81fc944bd2fc3562757d1b73b799d1c17145177e00159171b5f241f97bcdffc32b975334ed59a57122344b10bef4f2a1307c723e6d027895917a2e69a3c3902fcccc938af11230713d8f67f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdad97d7c5832ea24169d33fa9fa3de9b6755d8989008e8ace2432381ce3fcf58bb37f1af9440fcd1d45358dc8218b1af613734025adc32ebbcef4df81dbab3e6821237b3f23400b9d65ca2e330bae8fad393b478f027452aef847329dd12d04ea2397501b63aaed4d397af6789a49884;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde2bf7dcecc9a2816f738aa067c97438fa3539cf94812cc3e0f4600ed3106b4cd75455ca4222dc4dfe35c473e16a6ea01432b64e73168656f20d6c4a1623fb0d94caf0f0f1a00f2ebeb721305b59c45684820851e16d24e34ae00630009811ad904e1503463df5dfde85665d81deee3b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2167bcac740c620c401e51bfc6cde02ce4231b23015a3dec702e3f0b6cbd4a1a34126731f2af98c672b5c91d248b12e031683ccd27a582cd0d40beb681be88a86bbb14d02d3f838446cbf2c0830d8e362e642e94bb356e93fe6f7a4c26b6f80b4d836e74902a867b6a7363b8318b19933;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20254cd6d4eca2b4df509ac525aac1ec01de63e1acfed20487bed5155abbd314f159c8e9aa91877c5e34814cd724e4ed7cb4bf22c76609c5c83475d832705d5892d60ce61ef64a68b92cdf1cb96a3e2684ae29e59ac6ad1600d7cfdcb62bcaa5bffe70e4465a033f2a61e988facf3cfcd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d669675ed22f3e1c0534272ea8e7867482c56997589986e7046e9ed3a80d5ad0061ac00aa92e590328556eb0bad61720f2a3ca9692801dfd5ea8eafad25f4f879eed274299ceee389214f8e42bda757a57fad8bd7c7f350243188f574d2ba9377d5401e1e222914f23b178e93592eb98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4d1a502c22a7634fa4b508eceb073e0688ee7d35c3af21bca39e253c6062155c9d34b090d8ad96e3e3b93f8df6943f9a5708f911fd7cca43fd16023d497f5fbdd033d3c1aee548dae907bbdebdc39f23637efa6269f6d558cfec525719a5651432e15ac0b86935e847146ae6bc88c4e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c41efb6b51e31df7e2723a49b10f15c5e3be54b9e7f5e6d45cd1001da371714a2d1cc174db0087271ea8dfc29d34362f37fb736206423fe8239cdb62e0623d64da003c2e294056954a9d02888cde7f5bf3cd4a11b289956e3acd5f073eb6d37251bab6037739781533f3bd84b35aef4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99cd454a5d1aa888d59c1142ff09bcf32ce2670a172a73d738b86a7cef34e0ca0c08c97a89715d40f6fbd1871e518cdbbd17748721933a7856f9d3b7a151ec38a0b5fbaabf63fb064705c43358acce207a3bcadedc93ff6e3bbfc6813d8aeff1fb92a5b4263aaa4c185733cf14c51e4f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9966f2665681ff0b1f302d89498225b7d667b574637e95eb33c5dead6219941275fb6ad337b10c4bbd0d0e54cee985a4ae6643af96da20cf09a2ba78283510c111bc717004692d18d00940d1e9371aab71c9280ab116f7dc742680a3013b1fc3fa5a34b2ec400a63ea42a6e821e2c7d6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee3c9da77368a8f283a26df41756ebf113970d9278a491e3934f8fb4d53446ac6d30837bf57c3af1b7ef186fda98d3d8bbd9efd32aa3c4a4d85e2cf8f1615530f156e42a5f397fcabd466cc01b4ff88700dceaf984f5a77fc4a4362e9bf7cc040d9acf2d2699be3c6a9995c19593080f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5be368adb9645c3c435a7dcdb04c9818a98f64e2cf2ac930498ba16ecd64c250c61b89b8c04778236af17c0b9a73d68355954e8085123a5ad6204a95dc686981fd976a7150b7af049084457db399618ba08c57e96274a0e860d7bcc3587d2e9e19adf465c7eae7b924b614660d333db9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bab5add04a2af61192e48ba56c3268ff6ad9a0314447f7a1ae5ab172508f64ddd6f36623729070b54877312f144ca02f6111447f4d2dc27570567aa78244253b844ca492e297c04b6e2a0fa9f17b451fce39675407b5edf545a15ee332bfbb5de4667b3b1e6968373a0da8ccb284a59a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49ba093fc368a8bde355e18b8f21659f27d19592f7ade343228e34477851d6f20eb733edfff65ae603405b7147980c08ac73b4055eae7317ff784618006cac997300badb1f155f431776663a8b108a59e6ea91f367f7e09ae5e981085cfad0e4e8ba9baea106f5671fdcd607146f6fcd7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha96bb33002dd233477d61ebc213a6b85e9793015e3b0254cfbf293732e45eb3ce7a066549b1c5e8768240659dac89a0fd06973e180d0880d93ab35e1115bcd92bbdc929b742d91eeebd260fb6ebefc488ed0ff3d0725a38ea008167cf6660b9e13eb1b1e4f13d26ef0dede8ac5f8b3d91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h117e275a0a93012b89ad460faeb4e770f1ecfa24913e212c16c6affa7735668080a087bb7ca0a290f6c17748315fdd7f2ea090d65c780c8d98c35cb2ab949ff0660acda9ad5a84d2d51958384c5a821848f1640d7a5e7040999cdd8b85f6a7899e2438a5bf886aa034dcc9f72f7208085;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd53ccf2b6be408d0e29b7612c882d4b25f30cedf0f939f75bc1031df00cef827fe72ba87433341c6ec9f01c8bf026266beeca44d846d4208bfd4b93e2adea0e477fe3fa18d52fabf073d9985c33d0c1deacfbec59b8e4b58a0a3bf326c314acad2e7d25e50f876027a00163e1423f9057;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f8d0261335c5f05f932a375d02e72465ed0f689cba878a8ddc79eba4e8ed8a4e93400999a7ac4fa3a188141e1c56c0ab2ceb6da92f7a33d2b23fe8d067f5c61970d4dbae1b47180671f52c034770d63cc68016742579626e118f0d4fc728acf95218b3acd2cc61d32759da2bc2632d91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f79dcc9b5d7af3c0caae3982fbd2becb83ee965fad33bc293eb88b6ab36b74dda0b2c03bd75dfadd22651431ed77d06cc21872270a4432aafa7a573ca84a83107df1eedc093dd52225162eae929eea82e06d76d0cb957ceff753632ddfd29b5fbcf8d91bb7e0b4b46c554e0bdab74fa4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3069bbc655dd8815341c0ff4a8b162a52b6d2ead1399a591628499ed6ad47ae9691daffda94800e58bed501a99b4264d0a95293e2ef7976a4a8c0ae15d5f83115931d7d109ac54cc67087f45fa498a449fafa401308d3f4745415abd4d0908e27392f9409b20c356673ebd104aefad3df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d52a677162e3750ce54009c95e0bbe0cf97a2b941586e685366dac8afa484104416ac56a935854567cc473e8743af08869dfa2b7ddb1c4dc8c8205cad3cedb65def00f1eb0acc46a3f42c8753a20a2d11068788bbd40f904be076bd1575db65d86927c7e0e7fa56c2354dcc2200b94c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfa522089e4562e98105a4b907a0bfb708571dd05b74003712b98daafda9c6f461e99f57e67bddc7e66d6178037a3b6257a5abac79a488a7764fb092c1020ebf316b917a7909ede8c25418ffb429cfa6ea674eb6d3755a98d7192385e563349a797b0f612bb17d1a920f87e63b93fc3e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd52c41bfd32126747e7e33538d6b086b181202908e5fe85592bccec6cd02f213d3e0595c8279943918c36ceecc59fc37651798bcfc81dace9c62d27f66a100bce5a01501f920091d6ccda062e75e7c9026f1896220f8ad1a6b3208246afed9ea99ff50c317825d68834d4308742739bce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6d1a67f248aa33eb8b28a919c21ca2cf2bf19db5afade7fc099909341a4e6ad331565c828606feedae51b6a69c8f646b3fefa5af451e577a13414c40899351b0dacbe6481aef0be2ed89ca92bd4bc2e360c02d7f0ab0a565b2b66223ae81d0dbb7c5fdb207ce4e587f428eae0ff2ffb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54b676b5aecebcfaa9468276be63f3ee3369a01b1af8139071f191767751869c5d611a8766f30faeed7a809da8ba6e54de0fcdcc9a6f137dcd6801a6e04065f0180f66af6dc27864e91b7167176a9c6baecf4cf0cc9da6438928d27178ae0f1dbd8c3dedadb3b8cfcad8285d81ba5abda;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec6d5f8d590a1369acce2a3a92a862559a9363e7edbc36a481fbe88cec2047eaa07ba904f9fe4d3f3eb8671b80edbbf169a5b67e86cb007f4c55f9ceb77efa974d9fe84db31e17064576da34845cc4320fb5cbf4ff17a8c35bd9fbfe5f3f38a738ff5bc09a423b6625d03c4b3c2273b85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74b4f69b5571a8925326f2fa5c73271a70d4057a37a1a27a8c88862422655469f9a1e20942b2c66eef58572e59c130816ab2820007ab6d5547131900db213f3ab6fc7e747c76ccb2f4924a2c0e21190ff4ca151fa343e109cdb1cab7cd7364144ef51b2c1d34bf4f64d3b937e46a875db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a431f98e94ff3b5f029f62929ffe980caaeb3adaa5aabf314885e5469115b1e71509ce95b595159bfe6ea2bb2cfb78e5ce9c5ad47d8642da65076f1ef0376d1bae18903949a6313c5a16c0a5c811505f7773b3da5fdd9d789c04c56e703c9e72e6697bcab5ee8459f38145770df406bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffe3a0b9b1f77a5096f6df1a0f2fb721be8d08eff3030a1b7000bb0471527b82d6b4cbb413030301498a95ed9a1f992b026f93932dbe6d8c8e42e4c58cfec499814750e78f16f0fa82fba528b8eb3439f88a17c2c8fe469b5189b47018fcf9bb813e2b7d5a2b786f2c082ed12c699326a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5538c56c4e82dcd822a41b47b39b80881b98585180c5d9e2ad0bcb5b6f215f44c7f8bf72b407a8e2123ff06f462b24a9c7f5bd85c0fbab1fa35be815e719b57c8fc061d3543082af94b728a6efe227bd2cf4c61140354fa626386f88a8f1e5c3f2f2a13194cd5a4c2d94e257b10fe005c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h660fdbe3b3e2bb070c4423bd0c366427c4e6cfbe0b94fc9266e35934cf6d6ac3dbe8445c47b09898cdfbbe0eb47038bcb47a9773880a690ad6b04628c5b74a4e1cd7cae851b7855479e27bdf668ec19faed82a8b3cac92a41a660afe36b6efd922efdc02325bc5eb4d502b8647ef24d0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfefd9fcc4006b8c06b7dd25d26f13b35f489717a0f7038445003dac9eea49ae7fa14cfd15c95e9a832d34628d3f64f7d5004b033fae76c6ccb9ff7869d0b117b79d2cffd7aa672108b21d167495ee4adaebbd37340c48f315b09a59bfeb4bb2285e6aeb5c4cc4df3b7c42a11599728369;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf36d07322f0a1155a799b6d1b2530d43787db0c97d4eaf44c0b10effbed68c09b7dab00adeed4070571ceeadb24b045b1e93bb57f90b60d197b5936e8d13c6c842d1efcbeb6d8bfca1b3bdd85e7ffc23b46cb0a24c574cc95b40ba5e0bd5cdd09dedeb9381b9f54fe105a4a41669d16cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h430b7262d73c6ec53ed6037ef95b06e88e6823e9bb656d3bc11acf781af709fd6c50b0a69611bff0d526f9bf9093a6dda60a38ab06f222a70803706aec2e1ea15087240d27e40de4a96ed6d9495d0d95f76dabbf9162ae7a9de5234cd088d483c750214cbb963d1f67ab68506590745f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d551933d47a494d7952a45db9055e0414c3c2e6a683607b890bea6fe2e059ae4081736bc308cdd1b8915d4882a8e58ae6f2a57c1831e5aa1cc82ea1edf6459d73fb14a44ec25366c12661551547b4b279bcdba05b69aec246c9d4da1aebac99f1872b8eb6fd88a884a73c21c121edf9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c2f407e0c07d8e5ed11822499d4ea3d41a934a13c5c1f38da56d99593f069c3637e7914943a92dd5485698bf422fdf3a4b416ac20ec4e3ab5f06d85ddb3f051dad81346438c105e98bd778b169e7cf4a8339ad76a71744db4800dc0fa3b060536ecd4854789fe984204ac928c23d1ba0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf2e3fdde94ebd48c74c2abcc3b66727dcb17a6fa8b069fa3dd0dfbdb9336d6555c1e97bed0465e106680f41d487d1902f3cfc94f6ea3645f5cfd3e92b2af5d42e0fee2a9b868216561cbc1a818872558ced2c0851f8c2a801d3a1763f0c951187d972b934e616a387c39c35245f5ba54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80c4c5d92b1975a9153353ad3c62aa260620f980fa764ca2cfec7d3f8f1d2473403a497ab3243d4718394161d91b956fda163e10bc3e2205aa39d38e845886a3d5372001b7c5796584211043b04ad1843a70155fe5013825df394afc108e8c0d56b9ea684a22f927f9777772ccc4918aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4cc6871b21e0a5d1c043498efe4c47e3a05165f0abf629c4ea646472e1281c1eb639ac7596f3d2344b9ed10f0cbebcb5a5c77f56f7a6e27aee740bf9b1383aab7662555a9e374240f70e3fe438927d19c5e12492daa20a4dbe9aed6fca7da63ef881ce7fb59671981179a1e23fa01c5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d88a05d257a4b35b9286ea7262b02acc1aa7393173923f30ea3a6fbec9056c4180b92badb40ce4afd69cd273e01068d827a47aae75698e4e6b8ff55e328ee6f4f46d8d2d1ccf916e695d5c5b9bb2afbbd36af12c981f28aa66ba57573e65c23161f400dc360cf45a1c719e04ab0a9d32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha453e4f5556b0e0e7f8459400f801ad3bcc9e05e8c65f8aef552f6e24155f1ee9e297194209adbc464d4bb6d97d03a748b99645bb43265cd91703da8fb60e051fcf01834567ee7bd40a2eff7bea796d08891ba270e3b125061a9307d2ada9bf5150e8439bc372cf10a5fbc8945fc5d3fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb00ff59b3cddf11909a6b8d3f67615bd7809f3c5f6c372a9695799f4cebc2a9503b5037ae223f64f7026da776b394ef94e104c061e22b58b54b64a91deb4187a5dfd504a4f398450fd7a42807eacd0d5540e40f1493e7f0d6135768637c51df0e23e327f0adfb6a3cd17e8a9f0e1dfb5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha114ff24990bae3aee1991cbe8c922bc17c949282e85cf5c1a114f5aac310ec70e64f085ff09844eadd50262fe86ba1cda5e235536108736231f179d586949ae5ef5bc97e8b7e4043f38534ef080a687f550f6f728cd24b11dafa29d16f08106847d96baa75db1d5852edbae4b653e982;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3414216c02e77d4320c41ccf7bfad240e4c14a6593d14b45c0275b22305b521d6b18d9cb5e6ce90ae0d573197dbcd9768542a618336b511ed0d4284585653bc721f9399d270b227bf781425152fe582003cbd753c711a0ef8e1c48b39d0c78250771e760c925af44efcf0f9b8d4887ef1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he23bba4049c88e7098e4175c02795bd3f80fce71761cd5eda13c5eaa680b23345df0f91cb85ca0fbc6614f218ace731aff8b72ba35f1fc4047383c5899a06e0833ddb9b9d18085b4a7f92af5cd20ff8787d9ddc16e842dc200090c739870177976809983979fb120a43f926300e73130f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbdffb038e4077c79abcf09aa488da9fecc64df4429a83157fd14da9ab39df80b11043d8496a49ffff80f67fd6432c97dbf382fc8977963480d1a84dd8297696986d64b14c59c94c252d464f54bbcb79d9231aa5b9d76e4f8b2d71570c482d47d80ce01b1422e242353bcc4a932a84cc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3fe10f8f62cf2308e8711ce2609bca8144f9d69408af4349f3ae09cd7e18fa6d647bedef90f87cd29f80391fa380b5e31fc036cdcf415cf2f5c3209a7b7630724fe28604bb1645e3a1cb98973fec2e6aeebd4f44a3b22492bc40b9d12c6b67fc4132b96fbf58831c7852add9cc04ca0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eca836896fe54ed8b583450ad47dd71dc776a0d32e4b83b585b1f91a76596061726d48a6958b7af7ea34a0a478ea7a5e17a389520d7c53ec08ec09788b8287b3e51322310d1dc0d7d7b1dacd45a386fd78aa9768171e01c2024e9c8b50be73ace8570f8bbe2f680fd0b0abb84d57120f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fa260bcca50411e4171905cd8e3cd4ec304d947605b50bd01acc367946f8fe5618beb371d0afc7fb2dbc9c68d673e82bcbfe45b8bba30325fd397ea38143854e613fa740b67b5511cd8d0f1b98d6ab86773cd9f573dbb57544232db19c4c803e9b1c34facf6d85754c9b3ad536e63c22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed57eb0b71699f9f1be05126c167bc96c2878edc7acd57dd589d9bc56c1bff72c4ede3c0d86602b76289829b7f8949b665e9687cedb3c9b637cb140f228ebec31368cfcb954c2808fccb767ca0672709d07eb8e526ddd844d34c7e94c2e42381b96d03a31de4a52bf06933fbc9380894e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19081ebde623989bb12bd0140e6782367be076954da40bcdf14ede71ec018f64eeecda498e299526e3d835dc9cfcb31104ad23a26f7800939e53a92483558da7cdb3d6ddb3983909c05db1afce177cc8e8df5e63c943a60c20ecd8382beacd9ade3d33dd05233cecbb77934f27eb03e28;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c7bba763c516d8659c87e0128c26320770ac6775a542355eb2126d2081bb67deffa70b239bd9a75a6c1d6776532f91e838c50acaae8a1ca95cc62fa2e66a505974dc1fac1375579b1a485b4b4b9f59ad93ca00507c63646023bc45760b2ff78097335e2984c6a2473967ae977f0f6315;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c44ff75ce731ff0c3e64bcdacd0b953970e5e602fd383b40241395d83ac7c96bbbcb37e9b199977e36013cb3624da972033fa64b0b9d005cbcc1ea1bd1d34ba0699029954ebf7aa48fc82fedea5cfb644319d76e2d272bcbb0cd8d827f8f9025eaf09571229e6eb28c958edab977b35d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6a45c9782056aa6805c80f8c4598bca251117156d623ed50d5a75423965e6e8908a29a2a7da0b27222aae2c3cceaa503a8d974f023ea8747027ec447aaf438b28ad9140629db059556335538cb6fc393c6aa790218c9334c7d9bc409da90a18dec23a3e9ec696a75dd5f7c1c17a545be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2c44df6e81cfdc09d9b206a414d5dfc208432ce7eab13630ac0b718ae69332560540263612e50141208ca6abdfe8b5a8a5efc880dc19c12f5c3a0eb0f7ba319e83a199ac16d61c969966368a76a2f4b132f4240b203d841f9e486b8e845013199651d99d8bd4331988b42efd230340c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b13e0752194d00b5ce0775eeb7e3e154bb4f32b1614feaedd26e9855cb8bc32c1020ca6782e32f47875ec2d052a0aa25215c0178f5a000a3964d890ef571c7e3a3b2afa980fc0ac7fec58b7d49c02af8e68a8573c4e285eed0c266af420ccabd72bc0216791415ed9221562709fe1544;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2af8f839ac33176353031ddc6424b0f1a8fb435fa9b16d0a70e3820c3ffe2d0020efa13da5a250bbd4642747674bf00574abd984f3ad1cce6dfcee5c563d2e6d1dfbe4efe80255350153d5732541b0b84a745e09cfc5a1c01919bf8f297888dda6cbd1e7bd6998f24eb9b4a86fbe508f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he60a47d2039da180c2781429723f6eab1f829e0b163f2495da653bd826d242fb15b9f3ad8b5a2e973d197c90ddedad3f9d2d306a930aa5ea1a2b1305ecdf332766b2c9dc80fb0288b6d1007b819ca4e25caa8b90190be28b9c529a5ea8feca9b160ffbb835147c9719447cd3cdc2b3b41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6bfddd22bbc90a4d9d5833de40f6d1f13f79adc4e80afd8770ee0680200a593afaff7cf6522d1ebe757ce14cc30f6b546ded281baa9420eb58341ef9ac7d233bbeab30e11c809dd1dc0d612e2cca9c202cf56f77b1be2f67084fa29bac8aad6f00d9c2d82b49f96e2e1a54f34cd960742;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59188d5b81362d6b653f6b81d3f193a01731530ddf66ee18db7202234d7bcb8cc72086965b329d0c6bdc2c44a5d94a152a9a5726e982ca01cd3835ea617211540b3b14f48462c9daf647814b6285ced0ff2bbab522632be1e0f0960768e3ffe1ebfbc2986e8c419ab33618bd3f37b2e7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1551e0a1ad55528493466060506de9c70de52fd84c4f6b68f074eae404cd74b75ae2459e0d37b0fe60269423fd50b10fc538cc37eca9a70b56b72346c6b902b0493a79c4dcd16130b6e461cee5bcebefa88acdb13292c76606353a5416f61921081bd5422ad41b691ac5bca3934537880;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h344b3c36b92b99207d433214fba85b64e51bdcd24f86ff1c1be8b553f38f4a238dc782f2949a049c1fdcc33297ed5e3401075e2f76f4f6c70aaca387766231049ca96549cd08567a0a97ff6246cfb4945585eb5d500ab01b409457ef1afa515ffc519f93f596ceef2a9e8276de83b2d9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd149cb6306bb408491796c6fdeabe61edf3e79f828d0d8f5b3363c8abd6020f94d7063ad8feace8f4032f57a001575ef5d09f3c9fce77eb2000c916e24636cda7460c81d28de538fb8952d22159d3c24a04df23030b8d8b626f986aef9f28563a2881ece8ea1aa722c2b9cde37624ef6;
        #1
        $finish();
    end
endmodule
