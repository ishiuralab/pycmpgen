module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [21:0] src23;
    reg [20:0] src24;
    reg [19:0] src25;
    reg [18:0] src26;
    reg [17:0] src27;
    reg [16:0] src28;
    reg [15:0] src29;
    reg [14:0] src30;
    reg [13:0] src31;
    reg [12:0] src32;
    reg [11:0] src33;
    reg [10:0] src34;
    reg [9:0] src35;
    reg [8:0] src36;
    reg [7:0] src37;
    reg [6:0] src38;
    reg [5:0] src39;
    reg [4:0] src40;
    reg [3:0] src41;
    reg [2:0] src42;
    reg [1:0] src43;
    reg [0:0] src44;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [45:0] srcsum;
    wire [45:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3])<<41) + ((src42[0] + src42[1] + src42[2])<<42) + ((src43[0] + src43[1])<<43) + ((src44[0])<<44);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e0091b29deb42dcf7c58d40362fe492fa9c311676472c8d692aa951e792b52424cb6e1622b259114846e608ca77cc451317dfcf4d6e27a6d7b050676b9143ee04f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f61b7120cce33456ec2114808c20ebcf74c65abc6908ff23fd0845c26befd1d9847536ac3a589f51e8233d79a844b3bc7fdeb94a24b80784d40699ef2fbd4e919c4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9b2160ce71d3b3d7c3d44debb6d2655ac9c44cdbd8e5db0466faa0703bcc45c9ebffcd7378ea9675d0dabe7dde0af316358467f0b2f1b7e5d4e6bc9ffcd2453f686;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8f8f80848a8f0aea2b2afb1b72cd6fdc7fb974b241f2ba94a0fc59b0e8e878592e5ff4a5c28239f225a9583463ff4e4945c9729c6874cad5b4d8c099117a926ea03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1202a02bd9d4d2daea1d508ac125176ca7012fce198ff5c58c67d17bd8ee5cccd3643b893c7cb59941d8772bea92c8a86afbe3c1a660e122c2ff8d8bcab63cdff7a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e5645353b1d0f53241f5a5bcd89a881446ccb362a3441442f81b86be43d58fcf86ab5bb03e379d5486780e6503e3676630fe1a1accf5efab76bc84abff79b18dd4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1354657fd2702519809344dad724eb0069be7fb36b5527c3ec8b48a7829846a0eb5b467ad23f5f12d2a2ad236992fae5c44646e62e4ca09ca74cd938853169693fe05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c1fe811fb9d3d89b21725aa694ddbf186c28ed13794a00077a377040ac3ffa587c9bd067c5c920fcd14b52b190c82cd5525180033f676a96d0c6edf2ff3a860b8b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc74526a3ec65280d4b796bb89c78e10d6d1d921539d3a505e756c25965c9a9db7d78257faaccbb76d9863788c7bc3023851817b5aa0763acac0691a1470fcd069ad3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b809f3b14524324e28eb16322892cd036720c11fe0863c5c497647327d762ef3f968bc3ce7f0a197e24cab8bbbf65b14ed6f3408d84c1dd62aff5969e145ccab490;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c95df1712f43b5d3741bb17929fd5ae3849b5796ee2b046972a205c532996502d575c36ec306b4d8029ea34312672c342695e24c55be63aefa1b1aac50603b321e9a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3b61faecd5009b2cf004445347270e8722aacf76acac036c2b07c46abf1e8a1694b872c1a5a90ca9f58ac2f90e893dc55717931ec548142538bb0ec5a6b90418426;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c837c2f21660bafcd537adef50eae2de9c04130cbbd226fac991e0b08051b5e584a74cb4333ecf46124e5c62e2581b8fad419afe1f493a85593a55a63a85e4db7677;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7d20f29d29e243bb8a26085eaa008c99b597e92b6b393c9db2d88b7eb80e49c3608d4143593141fb60d266f9753d6aac14eb76b6cbdde78c5abccbc090bf5b661eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8938dc985214dfe1d637e6fca246369c4f70eec291bbf0b4cd6d93f7d2f567024894e5c99859b1268726038c68b783b23f0100fe6b230dc35ca81605dc06bfbe595a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7046a15aa04e5ea1d81482424f0e46f30d56b1d8e6c1dee5b6b7c27fe2860c6f58ba51935e8b0a21c790537195e136382fb53ea6da3f10f95315463f8335e3adff7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1852378216c57ee3751179464207121ce6d9d0a27ea77196251d6191da2e5c37b1bcd26d61841f363f259a43badb28dc99e60f270560bd3f929323fbe146abb04fcd7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1375177a66dec6f3e16ed7f70d8bc0957fc945f19c3f64a7b6f95dabf3c86db83bbd816cfb16f7a43af32c72147097e353e85b6bd9a935429e6925daae5f4d78a395c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h278d83405792be1c0ac29ac0ee132baf3edb92f402e9df777766a39d235a1247ece84192f485fc094dcc6a4566bfd3ca4be4f270251e9cb9e5e049e0b5e309d23e1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1803218666f455560802ec08f1be3c473362ae67c9b50afc10b4515d62906873812d0572e59ceed45afbf468ad56b840453f72cb5d2041f34c112c6c5031955e43d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15375dceb434f684d0f875137eaf634a65b267035dd5dfd65f088e9d203f37c45c34ed0c2dfd0b86943e8dfa755259029b41f1cd241f783d241dba007f8fc22c6e33d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a53d7838e598053bad36b34aed5019c0038f48b0a40cc5e8d8d9f73a8117c5477ac6cf44b8fa2d972abbd6867be8e19d2df2e7a6c37ceb37845c76750bb81267c1d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9551efce8a2b876c321adb27a0b96184306c7e64e8f327b9e546a39cab057fc93acc62d3ebe6f6ab5c1219af76f1388568bf9014cf00dfeffe1d3067b6686b1b3419;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143845a78ef7aeb09202c54c9f4825936e3175de01ee7dc7999e1fdd83a785a9a27ed506006e81c9d1211f726c900b24e974f0e16fd825cd81f326e3f898f48ec37a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bea9733ab73fa827d7f9f6256e612962ad5e4cf792fe8f4341d19b6efd76ac567273c90c0323f9745b952c8fc3031453140b0275aafd69aff353a9b62a186e2baa5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114af1996d293d2a56ee28e3083f7607034b9c1aad898ede63cc0273c413aa1a465c768a0b1281e97ccf4dd27cc8340d89ebabd3b8a3dc61b7bc16917158e4886aa8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1219a96227ea05594345562ce8aead039269bc88060a89a2b92093469b187e8ace8b53d9a09b62d719a62a41c10d2c8a5f733e2d656f1d7affc11ff36927ac9b3707a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he43f82f90b2d8f572769aa085c0ed989a3215d1a4cdb9fa13f182e1aeee3a980b772ff115cbb2c1d1fa473ba08ef32fda49d8b348c77256bb2bfe620320fd3b94da1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8811617dcae716a76dcb04129883deb4903522e6264c0b2934dd9232baac4538ed76e7f9288dc9a503692710a52617a9b981c969d1458d11259299cabef7a534915;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb3331ceaf8b83817abeddd4d2c1e5484ff6d2670eaa19b09fe43907b4a5cc5d0db09d9d579b00239c138b5e8beca6ceaffe157357c558dbbb04b162463167fce21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd886a961782abd4f8449a555ddc646af57392705069fb370037c562eda3f5dc4b6b9e34c82052535a0e8716cb2a964c3040bd9dbca343d899ed3d959d548728fd68;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcfd7e35997c77725c19d0b02879cf535ea8a544eb828f543dbf33b74f40cbc35e6b516d7f5bc86576ba06b51eea6ad43b957bbbc7fe8320a8779eab5ca83d79e648;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173b79bcafbd54009f03b103d4dd47969d09bacc051723c11a861243f01b076a4a354a4e35483d0d19b82c1edb360111ad50296dd11149fddbbed56aa58a566803c48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec784c6f27502dfaabcb767113ea50fe3b3e8f117edf4063dc1e9cf6d0211d962d4dec85bf5b37b73fd56d57a26cbb6df6311546bc0f917c592576350359cb384083;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8c9414a86f20589d460850a8d27af2b088e1deac029125063578f1b8f1ffa8be596be3e498ba21602ecf5ae28baa8d8bceec7ef825263e4534c401e7db4966ddf04;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h598ce0f667bb0049c7c420ecad47298a5e97b991b33ea794df74220ce69cd8617ea3dba9757f93148ce5e7c6cb041ddcac7b418fd51ebb9ae85418d60a60c1055edb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc96718d25c5ab16ff566ae77417b94ea8b4e811d6ff898ae04dd3aba83b58e6a47047540290a36b94c3f17b2f426f6044ab076ce9eccfc54369a4313f5b90d6e4b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba526ad9f247e6a9b7029c40be08378b1f354ad5a694323f4323be371ccffb822cc9d4311381f34e088e08e7684269c09779977e790afc8a746c6162bb920b4b577b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42164c84f31554e25b937badc0bfe6c21c65fa508c035a120ac177c7e94fde34d824b61fe7ba1fe93744998a48a0e63617be78604ffe746e8cd2b1fede08010880b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a7ab13ace105de90a6fed8eccd321be2c2154507a40db36445e11d9f7954393fb3bc9e5b4512e579d2b6acb6c126842fb27b38b75dfba1254461a9e630d910aaa9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b3a0ddad32dd0d490e3b4aefa3975bc78a0dc192fe76eafe04ed83199feabe021d5b77141cc0f3b86fd82d67d9732363e5fee3aba45cbba6ada6764aff323884637;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h33e7a70f25da080385df2070d396ae3c04c1b6fdda4f24b127809294bbe077e5daa5a62193036bbcd5361b0469ad2db968f943bdee7f223bcce52a44c4965591dc32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1036d0f432c0e9a18efffbb92a942549dab52f665af590e28b606bb6e5fd67e17e03742e2441e1119d1ebed1be7b9dbf63013a013573d76fabf40ef7f3d19357ef557;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb584999c0aa1a8a526bac8898bc103187d6461db3502d759be36d69deb07d0baa8abd5f18b84dbadb6849036c5099d4d84200c203ae81d5626ac1aa34086ddfc4a6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1422991e89706dc0bd2b5a435e91a8d024a0be7b9a4064cf773ef0c01885c4d59e32369cd2301a72ea5d9a83bca9a9be697114ab061510aac63d2205e8fc246563e11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3f4381d28dc77ab67d9ba4ef19c90b2a0526cc1d26389c2efbd0689d411a9a77a2a4aea060114711a9adc05842b6d8e6557833500cf4718d9d9d95c328672504fc5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30c23adc8866be35ffcfc9f2a2b4e8b24b082cac209d68902960b300b27ab7d7c510ad22e1fba14e380d0561b798b7cea2ac12eb88a5a9efb5f229fbbe68dd0d5456;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151a146e4352bf2a85a2c987cbf0bac5a9e3486003a732861ccae93462e8c961afd69d7ce0c342c5589bc68680a41e2d4fb6e564254d23dac63ae4433bf0576f12848;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7da538d821f3cc3d88321785d0cc6789c50ece75051c6337f0297838c14ea2e8464ce97faabd219d913641f359ca0d417fec60f67553117b5d6c8898e6c1edd8f74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c4afaed840b1c8fc3f8319584bcdd79c0a6b287478988ac890ab414e66a26850dae5d4a713e4a3cdc18be161d51cd0fd640b6b07b7578001858a5346226fe236644;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hedd4706296f8721de5dd80257b46400b267a263134379985765b78defddb7d10cb90644c17538eea0bbe4dbaea479dd420ff8816912a80d6231e1d14645254dbf6da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7ad6870fbca443fbd37e8e798105520aa4655085b0d7b801937eb1238fa2f9a607212de7aff6e5f1a71c64d24eead5573b0bb1bb440b6415787713b6185bb60a7b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1905f9ec5cdde75655c769342b56e4b11adf79fff399a72de7f8b40b2b3a98140b7ca188ef1f375241a70a9a28fd22098d7d543f386c74ec15d68957f2f535ef13b23;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49eec47cbb6e41704279626a48f431526686cb9a0ccae1a69b5c9c087b2872afeab1ed4070adc68732415f486661865155f2605c15edf7534110ae484e6cddb5732b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d903241af7b1d052211e3aaf0d0a91da836e276777165b5965403761c3edbc5503ab406a5c6efb804fef73827defbf7b77ce0c49fd6c922c2e1d48d246bcba97a96b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee1a51bbe25b4042a0cc20b479d94181820ced6d4a44e6685a831b09e9fbe2b1880bcc22caa2e6c713f37d5500eb6e6a05716247217edda751289cdf88d1a4f017e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e53cf820d1cd448d9fb3b4e68c02bcc9dfad8ee01369b58b4c101b865054053632034d1961e70ff89934399faf264134684e34eaa0983bfe12166e5ae7bf35f947d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe89ec5905e26ebe7d5da41f65c8ac4b23cb4e9a03b9bd616291e4ff3de32dfeadca1fbaa58455727f667a4688845918193540bfe48e8e6f69eb130024378a800aff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc986677bb2140037674827bda35e649e5cf22d7144ced1edcee2eb04d3b5e5624aae894030ec607ff69326028b489b198bb23ceacd496fdd1c878ac054de1849538c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11dd1396800a6b26adff04c1e7d222fa4a647978d0f592a27225f983a8713bdeb795e00f0f52a7080d2c5384544407f2345a888319e0dadf4b981cc218847fd8f399f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea6b16b508470ca8e96e485eb69c1baf06dea4fe8ab73f2b3da6ffdfb7c21052b82d8a5ca474ebfca8aa7a9948330b139c3b20a65a3319cb50e3b4e27f27bf73fe5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2be60838f29e9d0c03c3d161404fb1501bca07db919db9022e93aa6e1927b4b2497243576cc794fc1515bbd34d075e313e013c0133284e3b42c35f2a797a2748171;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bdcb893a49f81f9b3df70829b2c0e53ff83ef07bbd6f1798d3a5ccb187139ced8fba32778883f0fa535de698cabf6538b819f845136f3d7d266fc0a24ca979a93cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha05c13f74f04fb8bd3f54168ff708fca5326bb626c6cb04effc70030b9923a8d09b74a2b99ea5c073fa9c65613c3aca6a867c152055b85fe53cf81b921d349355416;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa4f44f80477d924d7cf1f151a7d4b32221d0b1c41e375a240181e4c8223d6e41f49c82f22ea139bd9a3ba43a48ccfa38bdb94e8ea327854c124c06c488c74166bd9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136130ab2ce4d386979962679cb9addd3d46910a32150950bec173694d2267005525634d4e73f3c506410dd26f3e789c71b48dddeeb131b40adc7e417fae38bb00415;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e3739480479d32f03a16e267a568dbb465c12fdd31f041ae0e46c92b3d03a216d598c0844fdec4aa12acdbedf5752dfa28c9895f544679019c32b2ebfe8d31fceb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a0d45bbfc30a06d843b714dfa9f48eb68558caf2fefacbb79625ddd0c68a4b9f041a1d8d35291b88ea0250ca7b5e1588da3dc73ce10317421f4d24c5d172abb7902;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f5047b54e03cc80d3e9c9faff3b053bade02341b9091321325e0dcbf5ca58a4c7ba4984da4e8df69c6839312c7b15dbf2a8452d3a33b19944b9e4c6dc266a7272dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11dc0dc7033fc90aef945a5f234a94b60d0647c2d7386f161c291e0af5370b9201886cacd5955439e6d3d287c630a1db25bfff8e535d3b85c1e01cecff8794c470205;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he788a2e7a1b44453880743413d26a884d4c57710530ec25eb179b771131ce9d5e2d2029d74c6c283bfb96e21357ae785918c1e475957adcb006ef42715375f5ba850;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1041d0e55cad3b36e1ff31f6f4e0307dec73c61180896813a147119693bdac9e1f55f45610febf9673ba6ebcd2fa692ae7b26d760ec1687d4da58ea4d598e4053a985;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4bb17bf0ab9d8493b79fdec55fbeb2f8a1a4dc2dd6910ccd13bb57d560ea861900bdf17c655a0ca4f5aebc2258c20d19c66fa1dea1c7fe17fb8802e4f48e5535378;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc907cb4bfae4e4cdb253f51881652c7b1b20f5ff07f4164ac29172acdd6a6c29562b3e03e36c833cb3904f9336caa42903bc81ef900ed248dae72fa5de5abb09f1ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133fa485aae6a1f8a9bc94348b66079dcc87121d4aff846b5edc8e1eb2dceeac1c4e40e1ac7dc29a943a3917f1ebdd482ac0d0bc3eea04f60004f5708e28a730abc1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb212ef48e85f55e684b8c5a9efadf1a7abeacaa1ff7ff3ee58c4e9ebcb6599ae4878bb4d8c39f6c9ec036064f30ba037df9951ef02d56cb829b8b04a6be29c765952;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18947301327df86a36202c0e55bbccc1aba52116e86d44c4ba2765cc478a0ef0da8e59e60fbdd66a83f51158a1811dbc2ca7f29e58a7d4dcbf9fec78e1d64f49ad31b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162f749e957967020989e57a5e43ceb1e67f75a4d772ac056e4780f20a08add2b1507df1d1d9f1090956abcd574332ecef0b8f04d77b89d4704c322b391c8fa25218e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1892d1c59a54b7d59228685297171e333f84a9ffc162d4f4df5220f4f117164ce2d28e01a8c2137f2ca8ab764acc4c059ce1313bf04a1ab0190ded7a17304ea852003;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5f1438c22c08d60b0ed515bfdc3e7e8d46a04b24feb47961b65a1f56048206a119ed709a46b2f0e4a7d9a2f757c744100eeeadadb7700491e5a5c4f3eea24b09c58;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1d6667f04c19ab06b0382861184dba50686e0caa9983403cd888c287646c6a861eee6bd0b4104e585a5561b30c60ce18db35ab06d8d84ecc93aa40e86e09641608d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ab8084b1d91e62d76bd8db7da6383f857e08cd82c6eea5e0d72f3211c83db1970fe443644d341c74c0b18b861068836d8e2741bdb35b353482a45d7e9202078cb92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ab38009c6314decdadba2f588806c0e16746bf543fb9bed3748a5080d96e56820c99b820d53f3a453d9783edf705897b095bd294af6a2c93988c79b1da2c838503f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f15d6f73b6ddacd730bbb044be8175966f248a6b44f2fe3666c3a49bb7b5bfdd14ce3cfb4157054c495f226766a28b0a4098a94e340dcf47366f9b1669e491fb468;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadb506a0ac1d8cb33dd14b5b7fed690b6181d7326418d8bd8910a463bfec9b83a436e785b3bc0784937227abbc49d6549ccda999ea4faa5a1031e1821177f23d77c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd361ef23672c0a43de344b3cb4d4dd5565d118338c51ef79142c13d6cfb7bed264d2ed6a67ad68ee0fbc9da8761e937f2ed871e7976d40a11701cbfbc06804216492;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cad463b7ceaa52798acb19335650b8a7c3943e3419ef3544d857aa24090a030210cc07631b377ea912742b9e1f7703ef625f08072b23029805e6dc664111995e1ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4e7b6a68eb588b8140556345820ac88f17e7cfa9b76ce63320738fd374617a382866c5f26ca311e5471ba0f977c294cf16fbc29cad474fb712b38ce6bd2e989ec6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5b7d87f25f4769595863a02ad0d58795d1cf6f4726e91ee6707899522998b9e646aa2de860957a7bf56c5e860e803297852efde4a48f3a939179a9bbdccfdbe332a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h331e6fa074f2c9f672cd15756cabd3c96f67f44f91d30a2ce55b78a964919f798f51b6d990abf43bf91d28efbde6deaf9738edb669b2c6ab06edd74bfc8d2fd40555;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ac2a41e5682fecfe9ee7e5dd42879654021ff8c02f9194a79bbfc62a4543927e6723aedb5fd6d1954161ad94676b40c201765b9eb17256d913ce3cb79664441218f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8cf0fc8ecf77d4d948ed949ba554c7ba99fed15f941a11bcef7ebcb3c5504b37c635f67f3b5bac9e6a67c6dc0bc67cce91831698976cd9d4e882070d809972a05e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h862b81ad50e655be9627d39b5c8735c5cc381007cdfd3a2eff2fb74cbf2b713cdc0c74a7a555205dd2f2f64dcd04481537c4d92c0a2277c79da2e646daea62c64f98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf83fea040e08eba3a227dd84b8d5570a0af34370584e53fe798e6831c07fcafc9dd98ae82c9921a975383a351c2509270049d7726bdd90dc24564d7bfe22b9be090a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b75e0d87cb9186ca8a2a07815a1751c2fe341aa9b97b779821cfffa65a32698f038206da6e5e088bca84cdd04efe58bde1c85ce4529a02dbcd08920474f65cca9cc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h515e5094a37cd6cd526c172b6e59261addb19b58f9b7698354e47d994165dc29f0bb76356903003654984463b17092f3d16b28795fe157e619258c90c88e64c21203;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141883c8695964c345e3dc575372c7ca5407815ecffc627ad168c7a881e6a39179dde262f1e9776436b4cc459a8c2a7d1510a7f1ae1b7a3d10bef7c1a2fa1c2204031;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36c4423e5465fd90647df238f14b24b463e3a2d66264ebda92d8c8280a2acb9efc5a906646f86494139b18b21ef235c1a8ab8c3740423a3b25b2c864537d86d29d03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1604c110ed768c594655e3327aaed84341a745a437814a6e6865a4d6897e042a418dc59409e03a7e6cd031411f848d128c26c0b4f8f2b174b00322dc1cb50c75203b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h255850777ebab946208e83d5d9501f89db0dfcc78d31794ac52b24b77f70fed1a85b57a98c412bc9f02ff98878b0c96097430a9895106793009615633ec0c6e33b77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93f466a40f12f913849f904a20811090517a13ee69addffe3b0cf98c8dea4e7e908a532f49513ee21f9dd1abd80879014e7b92f7a5c39e49bf37988c9c05fef2edf7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105b026ebff65670fddbb9d99558b524f27b6e0f12b5165899f0d124bc61ffddb21b11bed4fd59d41a4219f5e0114525c6e490caa0894376b2805e9a1bd24667b0566;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5e7a78ee5c546bf36545e1895e911afff44af3dccba595b3385970be148c0c39299c349ecb5bf84a1bc27e0b0a736b50315c795a06f98a6dc7360d0a554e82ab645;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18976699b95be327751213a1ff64048edb2363eeec9db83ea82816036512e6a581504af76baac0b5cad5d42cc26269e2020a851a876b91625c5cc2ef294ce37d491d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17274a5af440cbecfc6c2871d7dc0eb15df8a87e3d2ee97881747bc5e04abe614303d6d83c772dd81ed89784625aa5f3af831ac51832b6aee7776f4265b024a29dd24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef9fff7cc9ac4fedae55926c03a8e5a849afba0011dd8cbe381f0ab33ed15251d3881d1a94c1314fb5a03993697132b2c056f19c0650a43e6da9aad86ec8c4421d8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a7124fe5afe03cd92490a0aea63db69783b9c16515ed1484788ca63fc17b5cf00a275b28ec683583c714e2becc84e54d274773c7f2ce3fdd074f2084016a17ff991;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11298a5fa3a37adb12a746ae0be86e32c07a97db6be0d12d2299804d92abb31c18bc95e62e4550b19830dec3f3239194837d957fe4cbcef45621d0c8c311b65b8d8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16230e661694feaf34afe905f77b961c9d9021165db42a7ca9a74b43eb7207615001064210fcbef323f5d00e6c07fcdfc3dfdd1f5419d23e02b58d3d42bf27c390059;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f35731f43feb8f5c3dc383523597335f2a82e622ecb7010ec3dbc9991494ffef538a320e439010adec83bf2ec09d36144b61f05355d350aefd9f2fc2ddc3d5b656f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139072c6c943283d78f777ef985618eed7597e2bf3a0fdf47daba2ee48181137e3b94df8722b7d98d2180aa8c932190e0ea6d3e4c10d179e8597c75f43563b28876c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d27dc91d50c6041d81172d18a79c070411c651bb54c64faff6ee6a062bffc165976ea06cb148a828db980472a85738969412116e335ab43df66c2f3e98e5dbe71820;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134a7dbb7b6b24ff7d50f323a3edae12b8286c41110de7734e05e86bcccecd6f55e3bf1e227fe7788dec0dbda13304a83d18e335fd80f2b663d54e8beafa8de0f188a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19cf69aef11bbd424b451ae918d2b00c39da298dae1c8fee1c098db3e6815b9adff3a944aade691c2d8d32b13c67f12b22571a6a4f8359e0e3130507174d721c43579;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb432334cbd5c0aad12275e266b83d3742ba83530442734eaf2bfa9765d3ccc6b221e9b5b11172308cc496eca0a280ce142edd73771e36b274d81cc9317974be8a6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h446f3253321685d0bd5415e5361fbe64f887d7cf3554ff9500d260912d5a0894bb256524e6663abd65de46f2321daee7b3b2ea6cc0e7dc6f9fb211eb6a0cffcf9ef2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d774d2c03b512f9286d931d3b1bdd5abd735cecfbaa7cc1c2325e33b9eb55a68b6e2435a240e028f67d1bb661498cf5026604849af2d306e74f60ebf1a5075922742;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7c24233ac8bf92f64032d78deb344aabf87ee96735821b1aae5971c042f198f5587956d8dc81e2cefd14d8d78116a5ba8ab2b7731ac810a6c82d25d3b5c4fd13603;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cebcee23029581c351c9a7a4ff8c2d228d7a4b6c81b558061a55669c6df3dbe24065ae050ffaf127be21db710e82804723940d389a0fb92b6f4c97de815da5b576c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd169adc9d339cc6811f13de666c38f7e847a6d8a528ac3197979adb2a78da8d85794d6c9b1fa1aed0f6b3440f207116084abf97fe61f5b52daac977de2614183a9cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c82c8dc53ffdd1d284e31b054250ff243a697568ba9efbdfc4a5581e1701931d1d1dd8f136a010aaba7e394f77865ffc04d2455af13531becb46c0b0f203331f15a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55650573ed722eb898ed59a62e9b46c81d4045c0189c29ffc0d08d6bd758025c11e60190806c74a56ef0c5782218d1dcf3fe7801134b90650b2b68a7fc81ed8e811d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6cdfcc366f47f1e1fc9ec98b67f317a8078fab8bf84c339d7a83a387845309af1905a4200f92cecb3762eecfe95911603385e824d65fdfdda654bffc04b5aa23440;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bbac70e7219e10aa0c39419b894cbe87cf3312e87d6a1a3556f5205155930e9e7f19ef6ba17e008c7a3f34350ed8b4ba61ebe51405a840be977ac7957afd895318d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h570bea972993f3f2056316d927ceb70c7921b7ff4b141f6f3f805c017ee4dab6063edbd59d761b68f26e8e398194f755151bc04f68483a08380962b7fc4168d68f89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4221db8613278ef29c907f191f6f33146f40dc14f0341ca97440c1ac3bd35e32242286e919a9ab0072f94b481aae6f82915258d29ea9e2caa7bd707def548072022;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96acd7d7a12c7373766d25ec1c0205da73ba2f2d9ba15f456ea2e840638566fb29b2ce039d49b8e57de59f0536d7d8b68671ee6fc7727623dcb146bc00b5855fd0b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf3ce70ab88c8beadc61adb6491d2251fdd896f05004c1e70979bf4922a92210092352dfddee32cb184b02bb34cca79a8343f97ee823446997b3d21fd555c50ff1af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0a2a68541c8e5096d347003ab6976cbea5b37bd5e0e0fc8df6b35db76fa3a9e47c33a4305190c7241621898e2d14256fc80e4efa42fc6d319efda11833062f6a420;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146dd7ae6921e6fae33c7a508248746cc9e81f3eaa09a2ce315dc7bcfd55c10dce031fedfb8065f347ed9fbb5346c89ec2de52cbecfc614aca4a30ed50c693cc9d4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5056d79053e69625a854d5728dc0e02fc3dc7edeb250d385d42d7c66d2a21c0146e970ce0dadd770a5dc7be4d7665bb422749bd3a106dbbd07ed37a74b36601f7ef0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86a1783bb643916af6d664a359c3e49d2f9d764f43e64c7718cd8205276a49760f081cdc6d7fed79bf4485261e1ea6406adbedf49948d09630c22df16b19c3bd544b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1361d9ec31c199de780319787063ae91c623c5dfa8c7db537a25d7aadeac2b5f379ab23aab1dad4196e140242e84bc02a50585c2dcc4b76c9368c6bdd08221962c311;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2570ecaeb9cdd794a7a962f79931b0fef9f187afe01f091b1f614b45ba4d9ee627b7527b7b218d6eefd661bf3d2191a97204bf4dcc4ce37d0199d2dc85ff0772120;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc421f4052c808b3d69f87e4e1aadd7077643ccae0e0ca133e6485fad1a3e7c16975a76ffc538e4d26411586118eb8bfb889288ff444612fb0b3a8760c67751a04043;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f9fa2ec0821f6aae69e38294e66149bb485f2be9fd2bb1d4edcf99de214f141cd4159abccf15be1b641ef0a7092aae58e0ea994c16fddf40b2679eb8c36058641d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f0dabe24e9f7edfeb0cd6bf46fdf855ecac1412e5694b1a8d5d5bd8972f160eb6a8ae6e9e1a46f06533efbed5eb239775087d893dceb2ef0939ffb7832a6b3dbbea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170fc1ce742f90d15ed2fcba7ff01c70c37ac0742b91a96029e54993ad8ac5b20a6f0edb57c6e75da85376d01108f7ee3464b2fc7d90eb670428f1f1da42215c2e603;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f81c62a88e86c32bf29c40399925277e9a276a382d78b6fc398285451b2c4bcc91ee80bdcd3a482046a746a539b297781b352a7ffa0eaa42475d466a5fcf80a1c6c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190d7140ca2f1bca235b79a307934d9b430e635f1a96088fb69408040cf5b1ce78d8493ca912b42cf6978d07698fb50d16cd552829670c0f278a1c229e35c91351ac0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd59a9622d9a887cf62ba39d85bae9d0561e5202625c682413b4b4a9ebb83379eecd4357cd2d3d295de461ad4cad915a2a05ec51452c2b4f83b427d37ad41373d31b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c39b55e049d018cb34402162dc77252a69409189c01124ef6a4d58e0c0b7c839f3aa623951dc5ed8723cf41a345481f7f90b33e29f583bdba94dda887bca0f044394;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171e9597498110e56fe09a9d976f0f897b85bbbf702ec72130f599e3b7555ede8cd20a24f213fc8ab0354f04c99d800f8bb1a5776c0c3bc91f953ac6b0abf31930ed0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ea293f431baa2bb1b40238a7a6d580faa81ca2e382e7c59434fa87d366b69952cd5696900455c1dd89a7a09e545ee2af0e785d55918b48ce4fdb24ae977e5f71ca4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96dc1417d183ac01bc2d6470080434df6b2c09b496526b1723b994ce5d5695ed18e89491624904753c34d2e015c43389802ebdc1d26dd6105a4b66055d8221c25c62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1feadb02b2555d60c168772087494d14286b50754c7a85b726fbcb78fd4eba29433cb6e8532f906d2b98e5338e8a07ebaae875b2e54a10e28ea1977e8fc6f8d7b8470;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9f20b425b610be8d9c89de02c470444afe31cbc4ba5408a47af326a3ae90790307f6f45e0484b3029258ad5746cf1b932b5a08c63771ae273125da835b336cde351;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce41ca2be337e5b9cb0c68c065952dc830f9e1948f1ac81d01e0f28739b106994e6c42fc40cd4da0f7b40bd573e401c8311a570c8ab81cc629a9c58b84c4967481a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133f97b471fb0098b684ade0d33b82545db3414d62a0670cd6e857412bbf6df70ca2f29e58599357622f41ca28f536e29e9de24b85eb079687d83a701cd6d9ab5e644;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a084c30032fd7ef69d025bec750ae84439b08be702dc6bc72e8fa98f858e22ca1acbb05051ace56ae9191450d3b2b6ea03631342ae48b62d0fdb5e38e22e2b8077b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3b25dbc55c03f513f650214ac29680a2cf6762188782749f5e1c522c2c8dfb8f441b26e6e0bf7220a4fcf370acafd8e7551dda8023807a96bee4fe607089963ac5f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb4f5b1411ddcf549db02b396f67349eb0712b7701f00513706276f1c1257b433133dad5d6331e023bd02b1571344af9e93f5cfa4f125a19cc874ca470c0f6b93a5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39a1ccfd6e5f685ba12074634513822b1bd1823dc7ceb013ffc6f80a8ba6f854c4c697b88b8eeaf076b30e4eb6ff5720dc86721deb72b829cb40fd17b70d4bb05efd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9eabd0e869b8da3154c3e91659eed6630dcb8c670c3d96526758ab1beba7aaf2c679685331a713c893a59ba5bcac6a1cd5b7df7824ee2d97728642a5b18a0f7f5ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1975abf6bafc0f033cb0667ba42d3c6d6a9012fa07657fbd1e58e5d87ec60dbd4a8946af4513b549d04a13ddbc2f5d752ca70a6082516a1bba581dd91c7df204526c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h433bf1f7e978323bf52e106fbbfbe4c20650a01cadf1e49916549b77c5680e47e6afebd54dfc48fad2d7c19b65ee36a4242e35d1dee5c30a5c54792c4abaa4409047;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b9654c22c4ba6809421e3187db310bba3169dc8fb22f0c2ca641c4c2c52b936fcaf051fbd579e368506eae74839e6b1fc239840486756a5d70e541d7e9d3c9a0881;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f43a5a19f0fece2314c913d027e20630aa9c70753e4b993761602f0345f11b9259ded7da1980edbe4fa999143ffaa85fde73c48e83968a8a1886b438b3962fec992b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c06527da1d5ebe3eeb492ef08e248e3dd20680f828525bc6cccc868d8ad0842a2558861009560e06440e85ef1ca5c4de08e7b0b9fed5f6fde4cae8f014829bb29130;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5c705149ae0259bbf5c44089d6f416e491cf5ea16f0c01864a14902be69e37f90098a741cfa052c37cb87540c6ab4e4ed288c38a19d1d0eec7b98be195cb72f5c34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f09eb904ad8b501848a659abf38ada5450a9af0932c81802077bd7717f0867d8fb06d712fdc9e79a70d7239849a923e788b8b99cf2e401fa8ecd3a5b240c20c2714;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cad699f24f43ffd52b096a4631316ffe4a601a9b06a1056dcc525f0020f831ac9514bb0b0e98d4165cdfa50134f5c0d2a005de19bec627f509ca9114b78cdd73213;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c4bcc6c0a1bc6f2bb98bff71f9c63a0fdcb594c5c71091522c7f78a6f60286aa03e085e6f54d8bb5efbae9e3ccbd8aa994a9e5dd93760cf9b34cc00eb73e8ff135a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19168944066e943fe3248697edfbf346d394bf2563925619d89e449f8ac84407803a952d040e4c19f975c941fbfb577f45f07aad6cbd070a9b71b0b10728f594b711;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140ae14fb220b74068b7d656ae646d1798a963982c4f6020b87588eb60208abbf1a8aa05b8d0aa535abdaea3cd5ade0167f35df2707d30c7b8d487a9ae0372540beda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56d18f6bb3219e231ef6b0ef751b0dbedf5ddf43ed62634a9054c8b72c890f13ddcc53c5d85f905a24fdaa20970417aece318e85e7e1dd3bf9dbb4571dab8d7b5ba1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ac51308cf1b59e13dca8f031ff6cea39cf13ee4a0ee505679b3bdd08c148588818afdf476b96ed45cf3b5f61ac642c3035907867ebfd7e16678f2fe90158728f355;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ea014a8ca898a59dfe99f172ccaf304ba459dd70414445987a4251b109403eb300f1123eb090557fd0849495da86d6bef8e0bdde4cec6b18592037800602177ca35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb34c7542ac96c455547aa36d45c73c71598e36508f2b59b506243122261df80f69bf0cd7722550d7795c470a796beed6990f96c3d9ebf26f61a3c3d14268dc243102;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41488f28c32f5615165d376577af25aa26e0523096053901eebe947688ea229d067dc9ddb6e8bf2b2f20317725e9612e4f7679cafdcebc124c88219cba21f3c2be42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4124d37fa33cee0afedd9b9ae65123d266f25b85b4b476cfc6e2fbd31b26167064ec0c6217f29313a4164239572bb8e8e1bbe7c506dfbaf5e1e69fe65df2e9699fea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a598c9a6e820c5d022cb43aab5d560cb10f221ca31a92cf12753fa168c345f375f75a3f5137abca3842e7c3ff4f779511f1e437834c64e50ecc24b62853ad04055e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f49067f0f6f9565f431a1d64479b843ffb7dbdb55515926e4a8a69841d88e8dd4fff1a6fc96f021f90ab917d81b5adfb9018eec2f07322c0bc1279b84b07522328a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12341ee8b03f0625950953b81c918c696b95a1a1c6ad48f8bce9fca4c9b028c640dc6a60148a90e95d745d1b5b84ea58198ad22fd67eaef8681bdb2598c8900e2f874;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h157f93395a022fa9e8685bb022fb0177aeb3020350c4521ad6406ff9bc3047d37e07118a99ddad92bea935552b14324db8806f18e09a4dbfa403cd78a59d552228d32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fde06184a6b5e8aa735f5cafb4c7dd61d801bc71d747c5b7d0d0d7f252aa305a4a62585ed9182b272732ce317b47a3ccb30abf0c6093ce7fdb8a77df4da9efca4e1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha93c31107e0e214e60d3d880653f2c6e388be5ed0ac6a46269ec6a4273d5ff6e671399abdb71967d3d45753a154ba15eaf3328b8ebc3fcb6d76cfb30b7c83e861e0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6267d8fc4f081087731810865203e8e72efe18c73bce2bfd7068d102974d4275e372cc637956df9313feba15ca260ea559728c7511a30739d0d11dd56c11c9a46a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144dd4d7e7b17f48c7782a46bb2de81cddb8cc24ce3d060fa1dff97c64f294272e5e4bac363c6b393d9dc1cbdfee6b94d34913f3366a3895706a0b0a4e724b087fd33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187d430ff71e525bd217d90cc2a6ff81fd4c95fd0ea21ae340a45000c3c3ce08add0606e1b6460950d22741920d466ac3a571446ade2d0a34fba0bcb1b4c4b2bf6117;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f710feeea52a88661f61d7a5371ffe5fb30b565567433022315248b929fdf20c71746a17b93c304834c8b8125980c507a815817d71fe34fa4eec2d84f31000fd2e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1c0cbdbf4ffeb3b889c79dbadf446d16b15684dad75e500bb502c339a25ffed91e1f126868d862633701e31b0782d7eef9ae1972a1651ef896813c1d48475a880e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ac2199692d7441ac6f848f342833b819f959c9b2caa7ec0671193101a4db6c79131cb643cbac56e9aa5930e5c7a3f7413900e7e1defd4a60e141344f0a15b6fdf6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5d07af064a4afe0dcabc452aa52056119f2c179cbde60deb1cb34ab6e8b368c0675e39d0a96a933da53317ad0618bfa045cdf5d6cd31c5afd8478e659df8525ccd4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c9916aaaa906fe25d2887343e839e3ba6585c44ab2836603a66dc350554c236485d7d9b1956d3a82450f34353bd95fa7587c88a49be7cf75223be2b124386f022b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc70a11f510e58a7665f1050a1ec5eab0be3861e7e6f096362126392915ffe76a87ad156868192c8aad838203c8bbc3f469f005d9b06a6760ea47a45a41afc5ead706;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0b3f795a442d74f4233a1f99155f8565cf7929c2f34ea00e01b70bf6e6770184660e9749b65d2c6faf9cab5bb0da94d35347e485778fabd7e273d0e1512549b3d26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c97c26e06453def76cc257ec817a9fe7f08d4367a420d30401dc00886ef2cb474a96e0ece1485fb1487112a5531ca78a98c1174648efdd3ced600749d55d86de2bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf5b875e83c417c52829021817deca90c325a2b6a99f0bc46fc88efcecd309d58f40ddded8482e8890cdf608294ab4a630687efb65fd0940016f7024000035846983;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4e1f0cba0cbdabed1f714a0fa14b805502fb79155326a2591dea2ce4776a4a8a8946ea03896979ec5e2ac122b304837b607c40d9967e9b4cd5013a540bf1a87fa09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9f535d15ada50baaaac22f44d363a101473f7dc5d8863cb952baa8c2d2587274d550ed9694c0aab77f57e1b25c8d7ef1dd591fda779a5eb65b167fd9b863883d1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99d8cd982e3c4ac6b6c0de2ac59712738cb681deceb66e4a275ee579017b0703feff4f28ac36b6bc090e65f82f1be28ffdf9c8b413073df79bed6839173bc277c651;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccd8f57f2408b78ed902e1529d052746af232e42ae27134443e258ea2443552d86393dc257fccb1960ff03a7ee895a96ee322ccb8024548202a5cc502c495afcbf2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h715fcfd4e384da0a8b4a9854f3d7a2d7f959d1a18d644bb5f047dfcf0fe682c540b1d68d5a310a45603d2e1d68f27280508fbf4bcd300abffa7dc745583931c18a3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13385880cbf26bab68517825e93ceefc138338cf617e29f5d226f0cb1fc33fbec5c9029dccdb8a8ef6f06af0faa2c9a482a1bdb323c3f64c2bddae729f99842d2ffb6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91a63648b9f6a0ce91bd14d258a0006aa8c192eb30e0a328ca22c63e06e147bcd27e1305f09da04bce867039ce2abecbaaecbc5b18ed0d1c9fb85268d3f71ced1791;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc57c1e790b3f38d6c4fd79378008e11801e136f1c115bf88888ed679e967d4d011bb2d26c25b65cd3e0590635c1251016b44f1864ef75c4b7a504d49297fb29a8d3a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6a02c4368c86337a51628dc9d4ee2e00a19ad10463c1accaa54fc3ad71a1eb56f38d34e815f9239a14d768cfdb1d426e1be3ea254d6c705221edc0cf00dc0dbc78a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a1b5e6656369df47c4f95afac806eab4108ae27ec5d5cb1e17c5db22962ddf8e62e3958114db9bb1c45dc58dd734ae8a66de8528a230ed34c7ec78c8e3331b99290;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb885181fb0ed6768126a2f08cc8b4d922792cc0fc8853bc0315416a6b22bd0a986cd052c1dc18389ae1d2b503f7f19218cf1969bd400f4efa289ed6d2aac9a55d0d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h309ee47eb761c34d3063321b1c14f3077e1e5e14afbc71a99c26ebca2a747d79a5e3f89be52d85f34ed68ca5c6f76eb1ef640d62cd2705d595c401d7d998a086514c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd51990886b8680158ee67eaf040c0a8a7bca3ee3bb72f6695bc17d7fd6e817bb6cad331c75d4f8886430e18f80a9fb78aba7d734fd98bac428fec8df8fb98c168f35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3322119f333bdea80f451406bbe322f253c5fbe8d3d5c83fc436bcd8c89939294a6865e529513938bfb217d7df4b2a4c146203fb390eb06a12fa9fb1dbc0ebe68eba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda0c899f84801881cc2a7fa44b3aa28bf34415d04ab2bf523b67e85b19a11641f74e8b2f203d3749680bce0f4bc008abd56e54997ec2ac2a814f7322871977a1af14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df86fc326b27ce30292746efa22e1f7e77eceb04693a576b47c3049023e8c0449ea39d587c671d51af39d95208c0a91560955dd9fc4727ea70cfb30c7e74db6a187c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b84a0099fd047801c1c3c323628be5937f809ea42cf2a183bd49db73b4dcd8577a3bcd1cf910f9db2eb3a946660eee4e967ad08f1ecc49534f70b6401925a44f5618;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c01ac4f48fb631f04f7bc70dbd187c998f7d1027f27112cfa3f25360f04400e4f72d5c79beca6af7aa82f5355f276e63e5e4c858365e457fecb8c70f4e74b548628a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1865ac9b40db07793cec677dd400445689a32345ddfcf9cf01081cd678ec568872bcba2d7ca97074e95637c90822472051d6a29003446fc5151158898afef232b8484;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a54b26558ce3b627426c628a72fec7d3440d420b22a73dcdbdcbc85f404a33b8f6e7d79611ab103dee9547f90ba4283a3b9cc308791f467fa58e939bac98d38e595f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e505ae87ca26a7752e6df257af58689a46967889d3eebffb46056f91cba6fa9f8e6e6f711fba35b4c569b79b1157033928b3cc8c36c32f2b42f29398849006b8e8e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4b4e9a2433a31b81d67425655fe87f7c1693fcfd88567e9ae6fc533604e75756665ca59752e840a9c413ac557336dcee29e7037dceddd6b4da4e0509297e255edb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd148862053ccccb4141f0c6ff3b164fdbf8e959bdd74f4bf1683fee84f5f2cc8c2f4e7483c1a0a292b934485edb2bdee9d2e78334e743070a0df025887458696a65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f3380588267164123ac7c77a8991a3329fc7cb2a36e44391ed89e97828cdd8db1f8e080adff630247d41d8d2cdcd8d615b3f11f0864e469d06d7e78dcc859999c96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa555f9399eae3ce164a45b800ddf9f139b6a2e5f32d5b349e4e6bcc7ea6933d3382f923e5f884b1c31fa01b57933e09ee7d0b60bccea5f3d2b5e62aea3392e76051;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc5e347080cb9732a013ce85311fd7cc3c8b16504e25a122e7ca2e700d51950c1a57f4552f4836381d7cb29a64edd0d42f4733d13323411d36ebe9a39254e51b3aa8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e37ca165918e17458d79445d2cd4160c2e34cdb9eb44eafec68ae65080325facdc4f0946e7ed0577fa581cb734cdebcca9e96d4a2152e04dc5e0b2598f8278e187d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1586886a7c9c5b015af375ccb2075368b2fd7cb89829b7d8b7a52be60f13d196e106a13c72ebde07d02564d94666f01c5ec6a629ab3987ad161a0cefd5e36583f6fd5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94bdaccfaa19e35e4faeb123769be53344ccb59792ba4ad867cb43ad46701e489562e1010c4022ae9d21aa80c3172ec3a2e04c1dfa90e4718c00176b473988e25a94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17347b70b660829807a4dd6446d6bed6e5c6a071c2479777bffb5025044754acf6e641963ec3274b519db6916c8828613eeedbe68cf2fb2beae5c662fe392bd78b5ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146a687391e05b759de96a19cbf9476d269481d0ede03c9b680205492e4eb9aab90b9d22ac0201a56483c2f4cbc2e414f78c411f6d24d4b34b5841771e0719a053321;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eeaaa0bf31cfe1cd88d1cf2c32c70f48a696935a296bd8989af993992d8d2b0890ff7f987177ebb8cbb27059e83515d728e0add2ebc5ffadeeeb2a15238ac3f1e49e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161c689be91b65e5493262ca7ace33d175ece24464344dac9b509e36cef2535c8f8553d5f8d876d93a149b2bda0cc38d6c122226a4953c36ddad5f6b93e7d4d47498;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hceb9455793929cc06addebfa818e346be97c41061dca769d718f950c3a932fd542b2881ebfb3f28cba6a9a71fe1d13a5e0f64bd7054697f5d92748dbc4a8b3960187;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cc1e760f445c3ba136ef6d7e5c089013a56ef97240e693c9ae21766fb2d64fe78aa95c8d795b19307fb9167063a8fce2048f196b14e868264f2c34b4666fd2bc6a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3c818f4d3b4b59a1d205d8679982c4e2b7ef7cf04ae5b83d89338d69768262e1077c20e1bd1eb56fc5ec549d623632637c886b11cb2291f1289989006428ad802f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d7bc7f0e0d0052e7d2526e2693bef9f8eaff4f241714b84ce4145fb07f26f9c49f96bf8caa98fa7ca50d7de4011dc69c796a5b1b35be6bcc7e0634c9f0277b80a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118d11dbbe718cce46e847fc4220757b7f38685d0315674d8b5cacffe8ebb7eba96fc4dee30d38be53148d729dc07f07ab65b97861a639c5ba23ed9ac9a2a4ab5d1a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dc46258ef510dca8945d26ed60f6d37baafe344d142354a5b8f40ea8f0e07149086ee42157b085effd1c3ccd8103712d6243a930abd8ecd65d0d449a3f081d660dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9651954371ff2006c181a60a8bc3208e8cd3ecaf19ae0862b20c0e3e7deeebf3d4572ea436410409ccaf1b670339f9f5b2e800211a3c4a2ea71b465165d6d54d12a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2984928f920d0a34e473578ab583bd2de43951893c0c1c85fbf81f075a0054cad213139e271e995438c2da69e23ad5a05e7bffcde579456a2ddf4aaadd1202803270;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17762162ef0c3d5708112f16381f16a95529f105120adcd4ae4110f0c3febb404878bae7610c6c8c8c98765e9fb342c5461ef3570b810c63d42db270da35f3578b09e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159c8981fffbc9b879b424e5c55c3380e78d28ac307647459a67dc7f654357deca03f9d6599afa4027bc422dc205ee41d7e3f77727e06f8d5ef7e5ff617b6bccb031a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a5b13ad928f1423c7a7bcdafbea79c11db33bf84ecc08a5e97f9a5a6de7398910df82b659daff77abc69c76bc7606181dd1ce7da1c169d627ad5ddf75a94c7c8d7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16abb04873543faf17dcb626d9e6dbdd7cc62169278a13566d483d4a9654c05ad52f2093a98eadcd809843265d01e600eaa8294f56e77bfe0f5afcd5fad82ff53cbcc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f10c869bd08b0512c446df79c69247bad6436cc89c788fd9dc0d1d3a2b83ae6e3cf6ae3ad01b490c3c0f3186c2d5fb353ad45792672029e41f1b7598c63176c3416;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e071b1f0fc1ecf8af85ea2958df14c047d5f7a4f9aa09bfe232710bd0fcd2281d2f6ca51c62cee803831e4172d03f11fd75e306b53c1e014e9150546d1bbc9fe0a93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd2a8a84fb6cff5b97809ae23b6fd553afa84c441426ebeb21ea3e21093b2580d3394d69acf90330430234366fca190dc99138233882434399acaa604af1e179be5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4fc94ae486d6ce50526731d8b4bccec8ebe3846e91e17725249432cd5430aed97daf137b9a2962fd38298761d22fb78db76109a37466424c06d0c30a3c399bba019;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70ee1c0188329321b5c52c3f1ee3d7241e5982142b864d062a55d060af2b556e0c5d30736af113eeabeb1abec328ceefdf0b959448c57bf840e886fb600582a669b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c0f3a5df4abc65a2681dbfed5b08cbba8a63f6a6223949c2c106f6a255c29fe9cc8740e71a8e5f8cb968feb9180c7ca88d6489c8551b085053d9ba32853f249a727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2ef30336634dd6041ddfbed6d66f12d92cbdd9df8e9dc19631b451b5d40f24551dba1ed99ebbb9915ef1516b1afe64a29dc3e005d5a3dcce28cf245a7f5137b4bb8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10644a60ad378cc599ffa3d8b80b8f149c6961ad3aa46c6d0ca3ad4e90127f148f3ff6ad0e2930cd6a1d77e7840c0bb603268e519f676754f955ed64abb09d11ec444;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eac5759f5821060c55a4a00d373a8cc93891640f6e10dfeda1952f8980cec3dbf88265c9061702b6f00023703b1ee7888f2ae0e7ea6a54cfbfe4099b681ae29e497e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102768b21b17e39b0fa6f73c49e60d780a02b46867558fcff53bba19e7256d0479ab7411dc115edad3d7d6f52eb52139160cf0e4876d474c224a69d23a28c5f965475;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8e7cec2fc7f3a53aeb2f9b13aa44444fc02ae0b0deba0632350bd8c3a67a6b10459a13b4c149e21fd4f48aa7952116f9d2f2c21578757c010672e2ed02fa2f6a9c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec9aee6ceb74456a3b3bf01c099fc7fc0f142682819d81c2cfd7aae67f42853b4c1e666c83119610ecbd6e5361053e55fc1b558f0983e39c9a18fd06009db9875002;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ae95c19bfa20ad8a1cb936471f2e5fb89ae53c3ff3be56f51c5e68f7fc5526cbb4ac62ed048df48b4c5e975b3df16b5eef26e2d6e99fe3236492959d17342ad5cec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5bb79a3b33b2c14d8d6e853951261499d1f69611d4c9a14912d5fe4fa1c11f8a504345b1c2f7113ac427322e8d939fb6ae9a2ce3ee937864a9590a61dc14fc1520e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5072b66364de387696ec3972df102bf1f1a758df84acb4234e5bab4e25506724b77e6d73bac33bb8a926e624fe2fabbff33c7f488145fa3f9438437846b9238ffaf0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93ecd6d0ee381b09bcc0914e76763b38a4172a2f25a8c8b97cd47efdb2a863c0fcac23a76df855cd736379e4e116ca7a135b1d11fcf431569ee477ed02136486c214;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a326da022f11a1ad473c16c408e16e3fe24d76af33a6fb81865535400bdab0ba68056c5d9e56907bdb0d5413eacc21339b14dbf7776acf7f41415b7aa614663a340;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9671d8a99bea79992976fef9f6fa6c22aec4fb4dd721f692a22b8c711d9458ad82b6e91c7eae13a572b2c6d18d3945d9baa7e429c9b390947f4148682b4aef3be05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166f905c38a9d9e76a5137fdcc585f99d2d65499ceca3a66ff4ef6a2d19c497c97f2a5ca401584bf1c61ef14d61744e10bda5d3de624ab660df89390a1a542e7ca6a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9d2d9173f7cbc1fdbfb7bc09a7d19087c8f48a70cf38107030ad78e43c8948ebe5a3e1d42b7fc7dc3be7f06f8bdc16cb88ccba305b63494fa714ff23a13dbf5629e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1463b2efcb1d889660a6430660ef6e533c09028b4eea8bb52eed49494f22879726957a6587431bcd697cb5d32b93555bab6c49d5d3175aea7a406bfdc05b1a57ba1ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc11ba23ace7fccbb7dc78110606df54a8d573e90a00e8dac2f037d6b1f1cf1ac76f679f5263b5d16742a1cfa669518a5a6fa96394d0bbec1148a758e143ac0b5753b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd0a46c9473100045b9385730d61d7904806eea6d74ac9c63b21b9bf62caf3f77edd869028adc998c41d50510dbc3119d477f420626a1a2ffedad2d5f083c226d950;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he935733bf6f0c0e2d3bb9b3d36f5defb197de8e459b9323ee4db5a9a6fa7246347d28d86c27211804b1e24ded03aaf89af808c730a5e5d982ba638ff9136055a755d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189c9df626a1e1a25dcccdab7b29a6bcfb837d5f944b71a3a1fc0472ad8ad6e9fadc42eab7201dde0bfc196df213eee493ae01f23293000a79a59a761d2713cbc8466;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c03b06f0e35cac59380f9af3370c8d18ebfbc6636481aa3c909ad969aa0d8310e7b06229c574554b091ccf15b41d56ef4fa2c1eaf90b49892bfc8dc377f917ce220;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4eb5eb0ca840b50a8cb759922c9dd592b1732c9ea63ff4b107218bb02e6ab3f82571305cbc96b14857e4920cfb06a6330bce0f0b48958596f26b267a07c40754df7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9468061b9cf5c52224a9ddb3668db1b748bc9c198dff95842decbc1d4eeead39311ab9c8fc49ea9fd83f8e4b513250754cd0e9bb52d5d17b7277fae2810a6ed5689;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f5308dac0a934516c24eb8263809f7ec1f545193fa5066779b688ac6a597e99ec86e9e5368030dff56b9324ea4e2d848e9b19c6069d65bcd0e16c171eb7fdf6322f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5826918d6ee9d57a56c504c076a5c1fe0da7c9c80bfee3bdff0c220a813eb316fbdfe90369a347aedccf885b70e82e5f38549bfd1d81bc397cd6c5909164d40b6a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc50c2b234020f463ca43d8b1012e1377d5da29df461eaa3e891ccf0a2302d5cc4d56b6b76675126195d3dcb503525acb59dc3720cff9d6081548aa82e67cb4660bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5e52b3fc96c2a9796f60abf080c8775506517672ab68a7551707d67ac1ec61a9e02ea4231401262a0d8cd11470b7833f3cc099ab83a716ff55b6d9b161e65260bdf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17bd146391ef86ff4638871c8e2e9653769b4a12ca94b1355027db6213085871f76b85cce57aa638a2964f99d7643d58b4663e97170664a86b2ddb0b69fd67b14668c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9301ed5e0bc8fd8d5b13147f7002e81a8aa09a56f409950f3ea7f382b6e4048969d9fb82f1a4a162de11f78f98ec5d94c0d23ddc48a55e2dd1154f445cab5f5b478;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1776567af5af1ee1a8c63995d3ad4f9df236a64fc563b33be317a9def69801ba39f54456cf4d564a8745b0e93eaa92592d66f71aebc3c69f893897e2d68be75c1fe9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b89336ec8619ba6247fa0126b52fa7dd82640c8bc3a151e09bddeb885bc53fdbd159e6537e2b6aee1eea5aff6cb3b53a9100942947a544733eed7e8cf3b36efafc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b66b327cb3fd81274325eac3f716861350d1daa91385f7a42af495748c31909a5b40c9c2c1df322d58288607ab576321106cf596af5714fc7fd167f4bf9ae4573aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2ae4d3a365c827a9935b4a22c039b2acd652798cfe12b10364b06e9a33f1ae2f21fe1d5abc4b26b922e53a307631b6d997ca987c07a05b9bfa19dd2065d857caae4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124d4fb2332b8cab7f604df28aea5de29f5e5f869b7ef92aaa531ff550941c97ef35ae5c6c79e0641f84507e0c9c81e90d51bc71c17f6bec0f9023c9da94bd142ec1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86b7c121a911d416bbeaa08b05987188dfdad83f6154a05f4b63573c8fd812b6f09dc4997d3607e486aeb4217b6e0206452ac073c8141d7b1bc60062b622a79a7a98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be07c9e5bda9eadbbc6e95d180cd48497aba87d1e4451a3c71bbb96f18d508e9e1e78531f349025f120dc9ea0ae829bda4291cdac0ffc4bc01d7342fac1621447cc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b83d1555c94201df5ca43d5659cd882a89c15f8e8c3939480b3d9dc8e740879d691f1bf9eccc775d8ea69be4100a15c4fde85abab7303b413b8ceee9235df23bc7dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130c39619b1294ffedb019b3c4ef52bba9fc7db9027f2da2f10413bdd5cc1cddb23167573f0ac0d8df293a4957df4aaa6f53253863534fa5dcafe9da0d1112f7f6d81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b08cff96cb8f5478b66a8b751985962fa0690e0ce0245eb35c7e2f78f5b855db850b35976143ca74b9604a05bf8cfd07921609232ad967c600c1b949ac639ad7bd6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6032c1a646d2ad4de2f27b43dfb661f7a4d4b6a01503be40bd5df6d01a24f7f4f7157fad28d424f922a38a8c94214d2cd85b1c52c74edb6e8402b1c2fba413c6bc9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c095423a8d6bcc45362a006d25662ed07cc9c99c2e88ca303225cd0212fe537889eff60aca3c851136d3bf85891462d1e4c0145462da36c9eca10c46f2be21509b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fe5e4f1d5197e8d1a871a30d6039113a71c0c85d1d4543060920e975b5cdea4a8521824ce72dfe0a9c763bd0422935f516de481fad0745e60657870917728af5e98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8acc80837b7aba7e856dd3c42df1b59b5db6a131ae9e5d0358ffd34f6a07e305adac5054180cd664921446f779bc81c8a149e70bff52b6cd118dd91340b36612b1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b70dcd7fc62872b959c9fec3b3b66ae8cdccf3155a1e2866cb4b21761669785c97be61ea208973ab13580f6ccbdde6026af0a609104aaa331aaf6b0df48b6c132f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab0b8a11631739df96e42fcbc9c7fca6bff537d3a91a02e01bcee4dbd576e31fb143b3e8d6501c1922d073bb7e88d9b9c3678b91ad9e7a9e1ae58d08858c406af449;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49e22c79c352a0b28aa89890fbaede3331eb83eb2b44901ce2a52f81fb1c09e249449c5460e97c7c5003ab718ceea11e5816d5744e4d02c1132f679b3f6440da0efe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185e42b085c85b0f64ace85f9b39ff84a49c6f2bf51dc1fcb9998b77d5c4313cd9ffb430e66ee2a1e1c36c47cf68148d43e1ba3ae3f7b7faaa5f2204f2ebe652612a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d1f71b106394d6223b0257a9abccef909811d29b9694dc6b519aca1239fbf93795f72e25f236375bb40c607977dc8419fdbd70a955efa7d16c04defb712a81a590b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba19a0a76724c2cde8825708d1836fb26e61999eb965df52a21dc0b2d79a70e6e6ab0a21a87272df83705f63dc5c5f7d9d623c1b800cf5b4fb6c41e09dd1b20794ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ec61f03d929ede6c12588e936ce293565793ffd8799a6dc1559820667d68e90b849e50b40e6adda055ef8dc154f039430afe2e5526581a2633abb59397a09159541;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h632fc7a6095180596775c3fe8772030b5e41a4068b737c9baf109677bb80474d00feeb5792d6753d3d003ea7978f17f6caad6cd6381bd48d56c8e459aa8df681d3b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90935dcd603d0fc3e7911abae36efa4957939327b744b0aa1fec2dd3c0a07b50268dcfabba58be10eac378b58a73d3968843f58e54980eab662c1e924e8cbce30c72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba2eaa40e9d649d316cc42743565bd69462dea10e0eb146fd879f82bde5e88b95865a21fc378f96523b8002bb9786294fad85440e2eabeb9a5fa2cbf2009c3df12ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119c932448f1ae67fbc0f401c1bee54c6b0ce35b22daa26d45b11e8042115698b32a1c58824eab4bb5cd2b6428bb0579147ae4269c823c6efa2985b7a07bdc488f5fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e3c4b5270761510affbc4760d83c63710c4281fd8c48fd710795b496aec4161aacde86cdc2b3004cca1b65d776224312922879abd32f2f1ceea800a15d215d07520;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad6dd746aa6b5ef90d2a581ba61b0ec009c4159047897f79f6090c68eab14d45223c1893c058749eec177727c1b4243ad94c14146870f7f35591b56ed1811706a6a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3009e84e34418617cedf451b6a21f7841a4d0aeb67c4936ef9aa14bf79719bbbdf15f55625b5015d473f7e9f749f8152142e70c27dd1dbe06ac5ed30b7581f042d3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf96aaa8849d5531c42c6f8a00a13c8549bf4a447d29e5e077ff399bfd778e493940077eceb0fa8c1d6ab9a540b4c254ecda5e959dcd947df6a9b6f28858b5b3918f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ba8b1ebc6eff65d0aafe8a84507ed4b6fe4bb56c1f0161df7143f299812affdb8a2dae15a4316a5454c1cc594ab906156f7d0f3d12ccfb4fc6a795a087d3ea00245;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d9d4a6276bf5785de60f80959c024c85efb0c44123d1e206913238ff0dcbd41f55fb8aa3f6de6716faa5726481b44fe5f161c8f74531c13aac1d47d7f7e144b0ff3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb241cb490e9b08eca9f79a0e7e0022a0801b45968faa7b235e14aab478a20a9daa05276f505567700fe723f4f8809429a6aaef7e0060828a5c115393cb6d02570e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d2f86744240001e89f92c6423b08fbd7f2d5f85f709797aa59ec5a5e3cb58a04e9915337da867a5489c1452075c02829fa573aa0886e0a1cfa865059d3be53634e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd7621e6099e4ea417f758ff3f2198f0144cada7e618831860752e17e3d575d9d363ce5037d3cef2671c704dd989f634a5257c5f91d1a2c26d8e1d5afa7a574cd254;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18097292baf35d91fb6346fcc1a5516ff245fecdfba225327a3a8d3b6b10545c985c67c705f52c15dba8a376ba114ad79e4df6f2ee77fdb07231e73e19610d17e4490;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80a50015a66c71eddca9b6c63cd3ec1161ec9457b983ee1b4d0c0e7213e9b4cb25199d583786b243c3e815974311df9fa72d2c45f47c21751ba4c183493215c20280;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac8f613fcfc6c6710fb8007d5312b79bbeb5d391e93a6cbd22328204d44f6b1471bc198d9a727e2f901769c54fc1033b7ffa615c23057f076a5f7a57f688ccd22e12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61e5b9aa06e54a192dd5dae18c6d8e15be5c93afc83e870e185544618f075bd671dfa6f7c3487c34370e64b59fbc5823314086c91e0f86cc0f6fc9cd0fcfd21bdf4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f90218bfddf89993e527d40aff5383000ccea54c9e620ab68072fddb72deb0b6df76616579ddecb73b93d7fb6cc8513e264d26032f9cb77ccc3d898f232a24f26c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2d7698ecc373a16f36ea8e316de37a2c8879e66baf19d99a1ea5f38641fef29bc75ad5c23de1199251d329193df9fa94b9db7f6d0f5b02991d9896c8d6a8252915b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1775fe91420f99ad82c4b005eeefae55f66b684e2d626d1b991bd163d23c6d044c4c80a716aa3c015cc4b70849fe17d42cd26e7b329e3653878abfb79d1c9ee5d3bbc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9b37c7e92df2ed3682dee046fad42ad91010023171fdc2a880c05d3adcfd58e187351135e128556c901e907c3b61204fca87f6fc0cf1b33d081093fda839a8cf671;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1710995bfbe759d550dbd144ac3af8fb540b8bc2d6ed21a180045796784e72301515f7bd229795f885718ebea34a99337d3b90da570c031ae7be4384b089645b9282b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd80232fbbafef3fc2515724eb5e86aaac83329c3817ce2669c40c177dc2b5e06820403c7ead87ab61949eda664c8b02c885bd4753c926fbcb56b0afe00d696950553;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df451dfc6a86f2705098b161b52abe24a94fae313e79c3a5ad36957c2163fe4e807d2f1d3473e46b25b5db3bd9ee92263fcaa214adf4e1efd43cbc12ddb5cda969d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81d490062e579e484fe9abebabc9c51e1fd38b5decd7911219c2050fdb94e399b866cccb6072917fd3a44640b7ad05fa60c6eed1e0ba146bdbf2ffdcd1d207090aac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143b992a459fdd78e67b27bba1bde6e0f909c8c330d5bedd05423b0d7fcc4e323fe436334380cac5698134a65548d971245a14fc761b54fe16d8e789457f69a79e605;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ed79f4522ae1a21b1a13291e3ed89ae16119227eb365ced33a2df845bc1c09b92f497a3514f8f2cc21d9c3cf01bad72b7f7b0a41d40c89f06c6b8b4cdb3d5313945;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a103c0bbaeb17834bf8432103e9ea5f4899120726bc8ca60346f81faddea20fe026f3600056bea44f3fff5bf85263c8ed1da30ba93560f0f9715553a4192f3be80a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b55854b590feac0ee9aab27762807dfedc8130536902aeb695644f7a5c5a092f10ec3dcadcf144e63e2982ef476a3ff9368e4be0fc7d6ed3aa070abbdf50719c240;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e067483782a5103f9a009ba4ec6d1bf0d49fe58bf98f7ff6b0ca2899797e12c5b005cca59782aa72382028b80626d96f414a82961c4dc5ca8a9d64354c0712dbabc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c5395a943b240f98dc6b8b4405f435e3cc1182a4a538c0aaf6e9797a594b75589a66ed30a633bcc99bcb2f94faa85b1a692f76feb5f79b9e246c90825bbf0135c18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132e037feb7303543a6190f7c460804575ff8a82e3aec1116f58ea327ed662cd35bf49f265ac0483fb432d4931c0a1178949daf027aab4483d4fbba61373fe2a5f201;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be2109fc902407f829a4bf4f8d7d9ee145ddd444b68e7013e1e5a7765ca6185ae884f64d99f46fe9c69d53bb7650fb30a4e34d72cca627b0a3d80809fe1a40dafb1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h499d986d26d1584273288dde22dc49d4adb7c1c70b7c4a613255d1f6e079d9454cae3572eb7dd44e0a71c123fc8a7e7603a77e47adc4441cfc2379121d971fa6f0f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca441c0c9966d050bd1c588f3b709f3d43a615e806ac89999e52d8bb8501d2b2c602e55d1e6364af79712cc1bceb6ff7f76f1668bc3ec9bfaad20b05807f80a79dfb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d76fbd766dbfb6cf9c57b76417f771ca2319a3db65bc01ffbbf47b78c01ce4ca86c4ee6ec4c17851c3d133eb85dd83ee72e9044bb1d390313db079b081bf5ad8ca90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18054ef91a9265a6bc401d83d5129c97101e5d17bdaeed4e4592468932a345f28cff80843af49648f640648e0e171f8fdc3e983248378e76023c0829491ad246fc617;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb61a956e2ddcf20914db172292f99c8f9a2f4c3791d96e05ec11d4e80ebcaf82b0e1a631258eb6e047c483162e15816cd209d584036ee9117efaacbe97c1e2a624ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0c6241491e3e3cc1291b13b680262b43581d121f39beb74dab6908c51d0bdee642c4a7ff6b70f0f304094e34a8b7b8c577340788e1db6ccd5a0fdc8e144a7d5de16;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha571de0674541c1671e81615e3758c8292f807f912070d7f980da76054d8c3825ada6937c5727bb516d1d60e1cb4a9c2b6b42cdf7879893e271b1f4fd4bdb0d80ef6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146d8f5191b80e572bbefaa61926b7a7c22055d42af3cb3f9e52057ab844f02d12e06d61ee40a26368cc0f4c3d8ed68d905a58c2981748510e16a80b2e4002e6a7302;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b9a6b09cfb1fc5f5b88688bc57fe2d9b10f523d259eeb076dbf7724a314448a539af1c1252d2f2dbe508fbd089df1a73f0776329f3bd5b80b4d92191007348ba3e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2c4eec6a68dc1605acd161f73822c7cc32144d9f2049a9463297fbeca497f5b7bad4ba58d11cd3f5215b4bb62bb5bd65d32d83dff3daac256901691d3b23c0aac86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd1c1718c1c5617c0ada9e9d0ed94860cadb9a22a9ce7b75048534726a80f6e52023a7bb419b90526ec66ec0b7d4297c36c9ead161bb0f56d02cf8e8a30b810541cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb67491d06557c3954591231f1451a1573549a24969d2a775da2fc44f35a4412b78e3319d936e854734a064707872f365c95fcf3de4a8b15efbca1431fa62b3d51ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48eff667084a77c86c3d8c9585f82ffe0d6337e0ba1440376de29e5acc3f5e6ce6e08ac114515adff1254b38aae9b928f75da7fbdefbea0626403e9b9d65de9590cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bdb7649ac4b9cd46b0be4bc3b914f908e3acebaab015e5ca7a9baa1867acd2bc686fff459d47f8ea87ac092202bc31f7d10d898b495b8a648368b33466e0ce9bdd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d39dba92d0e3e5bfb8db397c5df21eab5e9bf9a715e111d729a4d8316942108eb11a9e841876420a7d960d94a675537beb66b89d8da1cb12f7f0602f4e6f4748a51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef7979d3c02ac5248155fe4b577c7e1d4f3c9f68a6f48509fb146fd84103698d9af6c93530157d480d30073b8bd32574a5a6416646c48976e18ce5e41330bf507fdd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa198b250f7343aae5bfd7df192e6e0623c73830df870ce6d533306be3d0d74910557427219eaa83619aaa63af66f252c3587913c60bee5ed9be08cbfda93e5010f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aeb84e3dbb99711b83fdf7fa7e36b43e676f5b080e52132155c34aa12146fccd1113df7e8ffe9be2b45ba52a1e9316dd259b79f773d54aaf54e1866ed5c4834da9a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110283ec7af36afe3bab0f365d0517a4a642615c96300c8aef4dcd9c18299cc729bbf6613728c88eb8666da08d1f70e7530bd7a2af5d2a81a2939c6b1868acca17728;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb1967d079e86c5de6162c7c773d7b1a6d821a45009ca82129e0e89fd1cdb07c5433a0782873f922a5ed168dc92080bf559cc34448a77cc2628d62f6c0ca1bb36194;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a9862ee0bd2265ee58570e6cb0665de3085a127f7fd797e9e6ffb9298d7222a4600b49ad7172d87f9761404e7e85fd74b5bc75675c6e3f4c4f950070c8efd402199;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c11f134c78c50687d279d0ae02d82138775ddc756655162e7f3a0719b3befc6b60de9e6c5155ae8df45e9043df01f52af02ada1d00fa1b07983bf3f027e70db1478;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161d20d804cf271fa424973719c34e62449f1a53ba53a39d3109263dddf4ca1a3a05751b81399ed0fc6c099efedb592d8dfeee544dc65d0cf1b4da755e7c3d5dd85e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91289dabdf8d79bcfcf00a87d3174c0aeab71626ff55aa687604b9493750c415557936ffe3d18e0f535d6ac14f72777ca94c7b009515505fd41aed7a8147fe7ab242;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1714d36e2f7e600e85795147be9d061e6b1510cffb92bd4474d16e840a6e2e0f0a3d314cf72ac407ebb9b55ac49fad111d874ac4f353a01732d043ba86d0c9e35d9b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163abba0a081d1372c926cefe89fa304cc4593d92a23e641e8b43543ff9cedc7cb1277a551d5fc1404c366df41bb9d024deda8a08ff9ee49916f9fad9333b6d0a1928;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf60c1f9e82ae1558a561cb5d5c4af6e98083d4fd56e788c852306edee16e01f94c22825a7ea17906d25a6d1e39dee7776821dd61c6528bde6d0be56b69fd5dda9275;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dd3a249be58b888316edf709a7ba57aae8d963ad2deb7c5ae700756deda545a7f6f0ac3c1cba3eeb7f94e27758d0719492e8cdf2a0f0de0f9dbd54c23e93b02c9c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ffe473036489c59952b381a576da3b0cc86a57a5269acc21711f529b1610260c97d7f1f8117cdc5e79fbbfa94110ab97b489c34a0aab800ceec969056262dcad957;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38ac591fe1c729a1771ab15722cefdd2b83b827a84dab9e37c24fbb2859e52a5cfb3c090f17512f82131d80db936ec09015ea915c2d526faee28ebd415931c59b9bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf8f84347f38f00ebe3a7686bf779b6226077783d9264a0bbfbaf0b348b6c0e7bf38da93655dda157aacbba27ce0f39176f8edc208359ea1cd435c85842d93b7e30a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bc7ffc4da7ba72835306f6bd379c6cd947464d692c4be44133e29ca59e763c2e744d0d9931f0534ed8f586c390e01143c444d37c74ed13d7e0deaf9d0276d052573;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d9a31bb8dac64cdcd35e5c0475c8af900296787facb7085e7fe83b4bfe6fef9d337411a4ed61290b83ae3c7022b42571d01e8fe98c3cb9cc90de2a887963701c267;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h864dbbac9d72a0d65b8779ab02ccc4fec02950da18e4d880ed5630c744ce897416d6530a831bad5731d221d8c9fba8ba73118f2e868bd5e1308212bcc008ca3d5bdf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13981d61178ef7150e6f5404ea2dc53f3b5c164407999e7245a5175a054c6a51bf987d95aacf6f5015b0aa24286c29a49cba6fc9f624015bb40c5e1fec46ca6cc2686;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe0acca51ae9a433f35bfaed2f5bc7524b8b0c8efbd958768f815e4a4384ce87969a503c5251f2626a469318952cc8a0e915f824ce0e2672321134f7b30435ff78e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2e365818113f833a4021927480dda8f3813dd54ce578c57bca7dc1f63be6facc8a72979389a28ec2711fbef1b4486f996ec0b1cc9856890a0770aa26e524d5e67d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ad7465e1ea28a0e4fa5a3471b11e84f506819d6b611f2028144ca2f306032ae4510ec2f0680332bb6bd30cb85a75e36f5f59de0892af1e6ab8a98485abec74db9b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152790ea31d4bc93be42be7c2b72a238109dbf1567164e2f0d053c0ec9c18c50c49ff98f5a383253a652f33435d8985639a9886c1f0d68e81d2a660da8925e1e24852;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1256a11f4f11f1f697f8de371d15f3e4953b456fedce0ca3f9cd5b76566e5712a960c3b38dc96edeec26f9c5359799eb85944637c2a0e90a8e173989d65c63972ac96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1959402fbac8af1f6f8d8e0f2d8f6d6f292da35b336c6959ac656a1af32e3899f645f76f96b66d099b37d18688259d762780e847a8cfbc75bee36bcb01176351d5ed1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d2fe41cc518c0d0fa78abb6aa523218d1879e95ff9d8b56e72510a8c9c5587ba4ba30d5da3c4564649d91a41bf12bfbca86f4bda79f2a63396948f17f87bd81d604;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b1c90d2e287a70c87cd01b95c1454f17968d23f6bb1d36c574df87775f55e539d0ba8ad6f13b59856f6a72b846f840acab936c44d6a3f26893a55ac15187129372b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3398a78c211a82ccb9a94b1bdbc4f13b968bde4c930808c97e2f0015fcac9d573ade797f6898e2500c55939a4cd20fe8835fa2e621014ac1a94b4be9bc2ea9a2d24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c0e7dfe1d7220615fa08e22c2568a7b9b616fbd86f5a7588e03078ed744b0917b7c9d00a98a3184633519b9edc923013dda8f941adf37cfb992f18fe187b28f7bbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1acff2efb68eb0ca3396585d2ed2c51f38fa12f1357186b82416250f438d2b849e99af23be27ab08b3f34e61faf9078a392f61ae4d60dabe3de48be9565712e88146c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f73ae6d350e4f85f4cb8fd6b26db7a8dfeca230719cae8f48c239eb50d2e04517bfde421b7086104aa0bef1ccc17422b4b7654d1a31cb57bc2ab84c2d636b8c39155;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb52fef784404b444759a1744a08f6d10a08e6a3d7de6f3cc6024295ca07b130eb3e5a18027bdad6899173f12ebfc7d20b77dd2547dde98412c698cbf5cffdad39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9781da38c521d79f98cbf88688c0e806bec9d7ff4cb738d85fa5cd7cd889ad1c7971a3b11e6f34f05a2e9001cc08b63e283bb8f13340ad23174beac7c61f67cdc696;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1826eac4347fe9c68b5cfe83943dab2ccffddcb9a246b785be099d2a299796f8c54d09416d4df60b25b9fc21ad88725463137c839b77f9f2b2f94e744604564bd6093;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120394139d3cfff079893018787209411ffddcedf5da36e11c548b7098a47acb544c3a091c9227f24b97da12ccb5d395be394f34ff89a096c23c60f3e23e147b3ca55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d9b930bcd99da26d28a53b40d03016dc6e7dd10b36616b1733970679d3ba4fa438cf74d82f0109169c99058e648b0598c0dd0adb08b367b1f384a2bf4070fd9d05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45b800e134e4b31cbdc8099bee1e0977f1667c4f5fee7bb736b3ed4db390facc32986c8d1898690bef9c118c3009c2c3f2dd2585f56c3e869feed0f14ffa2eaf19b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93f87969cfeae3ecfe85a9f12f59c268e830ae0921cbf7edc42fa2f29aac0d04c1669e4f4113b94e0607939b7b3f5880443ac074c05150a9a653927ff5024b9e067f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80ad17651b39911b825f07c29b6b5304856e0b6d718676e9dc590a22a908ba0b5dcc0a05f868c1c0fe235eba51f0154fca311768d1460806da1bebb59dc5b039a427;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a6b0507170c66e83de4b084844600963264b29f73276dd3afa2398d2663a1ff6e33debaa2c16c966d699f3e2f6d7f5e199e01d7ed9f6decb6959effeb245cae3a46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187d735f7e38136f8fee87f1c53b1cc431a49d189da14d7afb094f62c615420077fcb0cf36f7abdd1f6abd5fe55fa3b7dd3238e096ce7a0ea014f0a9d9a91c6595be2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ae78cc79f59e3a87e72199e9d1a0d09318a65a5053afa63e47055f221b9f3cf41fd85e22540086e66075ebc96d81cbf75d8a0d3589155114cea48279b5af2e125e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb85b0e24f15ec0041aaffacf5b8f89519e5a1cb3eb3ebbd453ecaf1060cc9010a1321a14b2dbc425ff1bad2bf10bb877ab494ac8d2ee5b1646a1a22b3a3cc74322e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7206e8a90b0423d9c1f426d42037a999fea762c96c269b870891da235d18794cc19dfe3ae27149c3cc49efbb329e4a5e4aed796e9cd6fcd5743c5c3609a1c907875d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e4bb2f1dcd62b4a628351b4aed5ab92f3731232d53a8a38c5968eaa6034b9cd1466a6e2bb9e67d9575da6a3f0fcb7a2909fa05dfbe2250ddd89c17ceb78e1bbccd7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7e334709e052b582162cedd8515f602717b9b3e95c6df003b8aeeb998bb459b63fbb4568847899e46a347c8dfe35cd3ff266451692204a93497ffb013f72a8576b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd03bf374fbf7edb003384e9fc1c75d03e336f18bc372f8d3995c8cbd73ccf60da3f116645cec13139ca4cbdab85078c1232f76e68c7cde40844a1a91581801cb59e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19094431883a6b01a104e4bc02a6c75debc96f1ee96948e9de8b36841d623b35b514fb77b833dd38ab3476ea97ec5e63eaee4cba8389027cb018fd3c5dcbe25d0a82b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd614f6e2d8385d45c70272943f61f1bf580ae2eea8dd088b1965a170f2637e7b8766fe4faf7768a9499a8656e82b207173b006e5292043ae0f67a23fe35164d08127;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e21eb15bf724b472c9dc0a6230d5af5dd744c944d4d4e0731d00dada050bceb0280976480185d1df03efa172abc0c3f3a0be035bd1f446be9880e5a88644076fb351;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dc04ce838eec79b32de42c35307c8d0f6f5a152f417643fa52a85835e2bc4291e41b29ac4a5c0d8d1d5b3bce19334d679ba1966875ac4890c7350f08fa0c1f08398;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae245009e2aae345191e8c4c9dc8088cd2ed62ce0958c843f5147f53f61a23895b8604542a8d797b12029db05ab7651cc93b5f6bce483510a11e3b9b1acb8ebc85b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153592e4cc1540146b1320c99875f75f6f4dd6fb40544839ec68f2ffb25158e2a795b4498d50d6218e2aa95b49d1f8d806a41d42c9e6c80756405e333bc889b3e1dd8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haff50461fa4385be57dcd175036e3b376c16dca8fc2d206910f71e042d093e0fb35d6883ffd1a305b1af8c00b48f710b98ef76b4690cd86d05bd7f015c04b3887ba1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h494d7088e13d12a14b3f6d042c3c63d9726f6e2469f81eda68d745007d7ad6cf1994b71b85f11eddea80c361093969df9b9eb72f6369d8396c555beb1998f2974894;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd976227d800abbec6fcf7d41ea8b36978cefa4c7da112526ae48fa7be351f39c6f5420e387cb7fbfc3c6d280976d7858b67953d619ab9c4164b342fe82a21f42e27d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182a95a4057f2b9e76376c182c7528d3fc2154c7b952d46c6c7f689fcc43e31d2e8c3917ffb98f17a795bae03a29db7ffbe33d154d8a09c340ef11d213e239c5c8221;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113ce7e4edd43a3efec6f20d97900dc96825ff18bce33ec461f57e33e095592c9e170fba10f75ed75c2b816d8585f9dce8440c46a49a2018e2e2a4e4db68578a5b4b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h211c35dd652b3025882a99ed5ee3dda6d997f1872c299c357b2a3570b6e2060627cdb4b54ea59f6ebc8e997f72a0d33d8e48616d80f1eacc06c8d659f45868ba660e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1648788c68407820daefa78560aeae71f34410f6ddcd97466cbe2ce9a786bf14bb78d95b4d06b7edde1c9d179eab9df4dccb593798c06c149f866d6dd8c39ea9d13e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc55fc655cf21e0300a4c04b2817307f50cceafc17e2113c5a6668cc3ff796edffc15437123c9c7962e68bd12d438435ab3b810169a5ad676c9ce8a8cae4cf2f458d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b489f6790df308deef60503dfac4305d1ceafe4078195cae2cb01ec3946dde568602f312f22d5407240b6063b0b6f65b27ef77737d26f6224edb7ce360a7e2a0219;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6e73fe836605b687dd4251ac1ac2b705107f972cb1837bdedc95de457f419c30098657df284da9f9fa1cb139950cb58ce4e754bb65e14fe113ed51cc1bfc289c6ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ba70fc058e9075c475f20d028675447e2ff62d73a7e31b2df3f32245a0dc8092655aa2a623456e9db41633986d0e0f0e8f2c566596d6b973cb3b24a8126cd048991;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53458141e018527451325fa2f3799f2eecfd4e3fe1f88d8a3180b3e51f39a63e43d71449966cf72551c03d7d57c78d96b9f426d8a87814c864346d409495c1743398;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad1eafbb119b3fd224a27094430751881b41588fc830f08ab9976769203c01571ab41bc8d063f9ed91dc4582543098c499bb94c75113dbc21453cea5d297a672736f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d234f98b04ded1429be1693637e800b8d7d50378bfc4e26ea1ac62f1a1eeead1a5139b08d41604337def6ad96b905da9a68a3291429e83e22a77a7f9ddacf7f8c55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e003d48eafbc77d6d155d8219640ceacfdb54b4e64140ab7d970624babf21db752361662bc637d2eaee5fefcfdaba23ab7fd99308483c04fce0b1a8184e7150a219;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefae7584d13f35a67eed62e87eafba55af8fd984918698d8bd255ced2e31b96cf338415c114a3b7fd4f85f3dfffb1e96740fc1dfc8c4bf475c46a3c5e24d735e37ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd3b0e0a7a32fa13f10a632320437a1a145540030bc0f58049a783ec1a0e5ad0d1be6fbe673b86f118c4dfc907b8e87e5c5451f9ee31958389a922276cc91eb9e3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc531905cb6c53b154e398c35ce84b8086b9cde80bc9999683166bc5850dc9b8c7e8dddb73fd935806156c0f740f99984844d42cfd376aa3ee2d314377005e628c207;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153d351fe280f1499b230b069ecb82180c041750f02f427cfcbc53b3403dea2299b9eb44cd49dd389f1c37f61909acfe7a672e32118e8fa95c1d9e0c9933b43b3089;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c1b51a8e419d0cfdbe2a0fff9b13ac2edbcb1614fa1e2983dbef2d243fd1d37d0a057b57a9d174ab45535727ce84c5b55f822229a0a5a7b8493e431393eebe3607e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b9a8e129e2d54b3d342084690a9630c78b37752a902ff4f113ed586b7216b868ecae37cf73b0475db5d1c38917afbea7d1782e0063c769a0b5de8e36998182cd0e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha26092a6ccfc3008533dd1ff09b8c9229b7df65f241a3d74634dfc1c7066a5244ad339a75fe1ed16f3cbc3a5f958ecb4abc8cf30de8afc113b252c0053935125953d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ec28a5de449bbdda14ce029cae45f94fafa093fe6411d7468e8deee193178ad1f7f7b6d019a3effff072b96b8a732fc40560925a5da06f36fd0d9159fb760e5a235;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54b5c491859f772a1878babcb52b6398a6db9d5deb8964538d5ea77d1c4cdaf978b964e4d5896e340ebd5db53d916d16fbf9487623e7ccdb2995fd6508ef002ef80d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17985c0f007dfc6fac78b9797bb2bf9b31b0e25f73acfa9a0eaf15c5ade0cde30219f1c486e1fa8bb8b1ce0e56b1c1a425e75d4eb2a3988ec9b8fff813809f843db8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f07928386141e78251f88f5b5295312f20cc40bbfbd90b0460165447517b2afe0434e8cc33f002fb33f9264f825b82bd85714b046ac08f30a07e29a860b4676b400;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfffd8554e5ba8e717565a654f6bd83a595a8b7e002a3134a6041e0f76d7516f29e61100e6cc51f474e5888528a86967ec9b57134cc019e1fcb43e4cf72f9afe6c1bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb599b7bf517f05c9bdab28cda81e7c1dc734d40e8bfec7e058d970b23b2300d7bdd7f0337856e357b70a4c2b2cb8c04add50d42af27a0ad2b35535d9af8380a6bb95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccf901ce43ef60cc5c9f418e067c919875c7400886c8e6f2a8860c1160604d568f74e5231179c0a874f1b4c833f092867d02a5ae8b3ac3d527bdf31324535333dd35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1261c6d193e0fae51a673b9674ab5fc3d7df13a00c8b102465b68273a8a28a5b779389e81ea9ffadb39cd81ad02e9b21f33f692a8700ee500e235eeea63b85b9daa39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ff8de29270e57836f9a61c2ebd007a59c9a6939036099b6674b9f2f71bc66bcb5cfa0214dafa8a22bec6188a92ae80290e07da41b53df90237461d83d7d97ae50ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8758d08cabfe1ba5f711f7fb3416fda560f4741818f04ddd5adc7f48f6489227e6c47558d8d8a854a048e8e2cc5872aac22cebccbcf7a5cf908f6c6e1e8505b9b9e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4fe0c446f65b0dd5b2a52e25ea3e619c2252b29495e25ee3aad0729f6f8ca5ad7ab5b1700d757c131aaf0acfa6bec32df8a030f5607eed11473b8e62ac7b5ff7cd0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6abe70884979ae051cf502e2cdffb3109b54d3e1e23636b170148d9aa0e099629ca8fdb51c6d62a17f42da3910649e335b175786cf586a7aebb8f4628afae87f0d7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a234a6a36ab1080aa7c87737fe93334449e10c4028cc0288054bef9b01845b93abebfae9c79e4bfc3744529e284eb52b52dea39607f1cc0af124a2f780c24dbeea4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9517a1f8547666fb2f2c5976c9816739c48335e13281338af4d5fd4beeebc6fe3e4030f8411e121099fe733f19694d4289f9daabfcc29904e8a9fab65e19f3117520;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffdf8736ba2c8396132b4dec7032b5cd07d758370116cffbb6820b086354c53f0d258ca09797917feea7247449c700d138dbdd45bdadea1726955716c54ad22b0a4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7d99ddd5ed07c4ff9c0689bcecd9ca7aead8e817ba05bb10b637f1d44f9458b7cb365ef6b39a68a1280405813accf70546e4892b956eaff8935ca3877554bc5209d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha43a3fc8762633abf26d68892c32695b250f623c03a76cb288ee0d1b2bb64b0cbcfd0e0cfd249b8d640bc9e9eece800e0a596ef8bf5424c5a0bfc5c1ec61fa6920f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108c8ea0a9b1dfd8f623a7ad0612345c3e989cbc2ad57248d9e72fc89fcc6bec47ae4fd5115a867ec9285e02da30d6f23b96e8b0a5c7b0ebde17bf7d3c1ac8cd83f0c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d1d44308e6e02b93daa9e4e4d436e7f462f3ce721098c32abb784137c76dcc245d62ae2aaf7044552f0e4fef5667ae44b5726f93a871d4117388f2af6668391f84f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc3d451ff7c8e94b039d31623467be0ebda26f1efd6e2cf07878b94b0ad3b443837f5c88aba1cceea96e3750240cebd6188c0c5723a786f6d5a17d6530f99570a784;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c7ce4bc7bd18e44da281423b13bf943678abc2c93892600668d447d3a3245e17688a9714d6f7609de2be56b61094a2e68a1f563c06bb37d78bf11bee0ccbe49511f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c6c2405f39964181b249f4110239639782837018d22a76ddfb8a15d742902926d7a9e09143117c8ca105c5ab9a94c2f9ef34fa17603574c5a85bcdecff4126e1afe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e5a06874aef3ba8bd9dcc74967b644c08f06bba46c2dc28f1214c25b6122afe3a078d5fb60b9efc22031197259dcd7160b0cd9c83e294adada95ec6c1470b440990;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193a9904e2e1f29f795c6636015830b63c43ac5efaf7b7eed62300d866bce1f574ee80c8723a6ad5f3503008b8f32fd3a2a9920f56ad30248d447c6e7d0a6103fee34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa674d5f0593b0da15010fe653688359ca4726b8091c21cdc714f10cd9c34c8ef8f209dd1045f3471b68af72bf0a0d7148f3ba4b97b1eef26f53984bb21bfdc122b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1650514816d6079f256927c1c5bdb44a5997cddd599eba92bc727dbfdd35b2abfa1d7e267c1f73a6aa46feb4c1830395ca0247fc249e96a7836831d2060a0dbdcefc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h216bc8640dbf64a423cf72b0ddbb1dbf1e658479ca0124e7e9b276d0ab7ea926880f2d7dda18cf617b31f240916c17fcfe91886a3f130b9d92b774c7c00ec25e82be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cf4b9f0dd901a7790c5f50780573e6b90d0d0a1d98000014ec69e28f3aaccf6a314de7e88ffa8dfc2973d5a4d7828d121a49fba3982a5b7cf2661d2125202a4729a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9ab8313e78eaba7b649ff6c3b835a442b3b17cd1a2291adc10543b204baad04d8fb953fee930daf0876b3458a0accc0ec1e93c873cf5f82982b0e120b44012cc8ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e167d3910a7464d84d64915ad6271c1b6bd75cdbc44bd8fd620d2855f50e395d15811decd76b376456b61767263cd71629f09a9806a97954da85f9255a4925e9f13d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38ca41446ac0d219b4604d6bc1d10efdd485817cfdfa02c50df46a9ace96e58cfc605c188e24d6a21d7356a6b1c476d430cb6fc3ce591405743339d997d314f09eef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48d86b1329b91e540a7a934439580429c5d34cc720a5e9cd4d8237c5e500db3350f0daef2e8142ee8398505d1756b885b43bcfb1682900fa1641df4b9e69c6925b25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc05ee1d3e58a1c96fd289e4f9ff22e364a974c9eda81365cd07333e11f6a17bd93c91e98e1d5a303a2232a2837a995dbc31d0054aa0c69a1edac2ef4979a787e9a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1100056263b55c6ac17496c1234c1c8fb02b425f140975632efc573b5fc118a5d422b9302ceffa8949fed444c369fdd75ef549e2645b26073bad6bddd1fca975e4d3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf62a28da2c3fc752030c33c2dfb208b81a6eca3faba3e50052179f7635e181bf4d58c08906efd15862210462abd0d1a24de07e387c9565ea524de64c535806d4033;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fec4aea598dc186a5d5979647de86db67129d239179d115419e00b418ad334ba648bd4bef1f09765fbb5ca465b82ea5ede057ce85237b05e8ed8ccbd72ab451aee5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8318e7e9990f2250f22de6cb8ff7d0d8c3f05c4ff66da847b7a40d220bef01e0ffb7043dc3fe3c07b6660e26cabfb7fa321213fc417fc56840a480b9a3aa2c8bc37;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1043f643fa5f8c248e50284201104e03a0a866da97c0cb837d2b4b32dc766e98cf498167a539c9f4f23e6c48724cf53b37ba7517e31d89dc28f3ea1752a1c85223541;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108d06dc655d3a8fd2a2b85d4b9636341109b151a9b759c3e47a82c47a224f81afe74b5d3e5aaf274b1d779c88dc1d08deb47202f862cc8fa3e485f6959a9551c1e5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5800033175586f7f8501cf36a4286d44a6e48570ce71a3d862038a81477508c2fbd5b10a86ad412f6b9d0ad63d8b444d21bb854df337deb5821b68ab9b24463893da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a854c932f31e917368c9b495ee63fbfc34dc8a453d008e8e0887b2cb01d959e01f8a4d6723bb852e157df646213ba272084b744981ed5ce992381b505fb6817d650;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58871e86eff5a6adb569a57b06c0ba72abbb490e172f3c5cc91af0d72244bc43b3f9d01cddd72e9e269d69f4f44ac65da99c26896972b36cf7aea66b246cf54ce930;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1475ab7ef2ddb659d3ecb3f33828aad93e43dc75ba85c4b54182036709d20743d72e20524d562317ed0af0fc93cfb44fd77a0ebe72718447cdbd5b2840ff5990d6d3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1b510ced3dc87b414c90e9e3b9023f71016385e2ee0976c906f117100b55ef44ec14eb1cf9722fb99cff7dda5808f95077680dc709887af9ad37b98c77de887abe8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2904af128428ed152a6d0a434a5ccb9ddb79d27c1aad6cee871299dd33eef088160d3cf24fc75fa07f7efc8f028884bec176b6742c1db44bc2ffd56ee950d84b333;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e12cfef713a49d657f230c9b1c2e1cf1d748ae7a8507718e32dace09af1e2fb17f370cc9e81f76e2a7f2455c594053d8ade9cd851369f85ac9336e6218f0d507653;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1204e688acf3c7dbee5b3554cf09d00dfbef359e7ce6f20c22633096bb466647fc654e9a9bbf577322a4475ff402b0ccbe6c12c7dd3efe327c9b9664d024a78692095;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ff0d85a0c5076733af85afe23474d8d684f526b8bf91e60d6aec34421682fe118336adfd5665921334149017b3d5213d53cdbe4a995b4b09ec3507b4b18d71dc3f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc107bb50233ef1afe4906c9294dc9af0251d9b3de93e34efb7bec4cbf7f47e88362ec006b1d2fc2ee9126ad7c09ee9e98842b43e3feb2287b66fc20570b9d64a3a33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6737ccc52788f7320ddf71dd1c38400177dec74601d83b014a0510d9fea86f96142d5f789fec91e4a233ccae5057aa10701100b7481d4413605b2c1b5283f824fc8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b30660bf24912fd56a85ea149462a82df6a8dd602ef475641400fc1fa812450691316b75d308f4cb6ec46619f833368dd0a79318dd02db9d3e80a5fa970cc71e4ca2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd69a0dc80e1862eb3daa29d29e77fc166818e56c07419c2a0f8fe4381edbb7ccb3909cb063bb701fc04f70605f85577fa021eb4c29f1440f654b3e8e855d570fb22;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1f6b23960cb1763a96aa0db4e18db46c746c7bf2b6370f42c3b664fc9cdee010575cfc7b8c715ead517e0e38d96ee63b258c5d74e8efe7a39213574ceffec61ad78;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc054f6afd8a3fdd3df97811cf3bb14c3e6395675ab1b2ea74fc825d3ee9ec044f6b2c65814a00108b97f3c9729ded7cf8ca32d7ae4f3af31268fbc5f39ca7224a09b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f4feb82adba138e71d58cb6f64113a2f4c2f13992cd5cec9b53b057397cf47363dce0fe23d09043757e4cd4125b9afb387ced7aa0d98f686782af3572a7b9ad1d1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc826daa62470d6e38ce20cc6a0e14eb708c906b0ceef92d8ebc35513e26251850f3844eedbadaf88aff5063a9cfb8c02c6ce5ac49eb5bcb4c2d11f951174eb2bec1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c201fcfc33c5ded69adf8297a3b0ce2f51d873c198aca0c5a51b0336ced2469524f98bf29c31043558a9f2c11708583e11fa830a40f87e28b019f2ffe86ba96198c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h911e5da1a7f2ce9d5e71a631dd736948c7a5327f628f771abf7b99dd9d733bd9ffa01391facf9c399fe48f3ad910d18080356f4df6d79e4ee40e14883a58d9ccbef0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he349c3005188af0e0e6eea6215976cf453ba762a9cbdca0e4d9bc79947f36ebe50ae11c516ab63db51a3ad9fcb6d20d323893b39f27981a45ca47747e7b548425080;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5b3bc1406b0c64828463329e8d31e51e1fbb1553f2a7ee915655f89e908eeab62f494d0a11f7bbec6495c11c20a458b16e29a5cc523205e91c7955a43502ccb1b39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170e7b651635c539950b12b70233a9b45dec22208c5658ddb7ba8e70c80535e5bf44e33a035011fe3647efab85fce6d5b0e9172100008bcd798440d88f181011c521c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19069d77323bc92de3c1353a09b5d3019a30379e91dd28330434bf2a7ce3d410ed89d8adb85932a42ac5a4595e05b447462ff0fee95b7ec16d4ecda38d660a9da5366;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183621ac953a19999f5b6774a10871ec864f4c4df29e1dcd691ff52e7eef9f7d68c31a1d960c09cf6f615805e896484ef2e8b31e282872df0ce4afe2b96383b976874;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10069277c496bdf5089bada27d782a15dd5d115a37c4336e20a98e7da89e4e2e471b525f8564ff5c9fe6beb61025bf42d2987a2a5c34744378d29a18dfe4c585ed1af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7037a3e2ee74fcc9ac2ac0b92d34516ffb7ba23f5cc17fa4e3ea2006eb895d8c31f1e5703138c03375ada177997093b1a83e5499567f95e0fa0d32dd6c71518a706;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9c952481d8f31ab1b8f4920294c5b8fdbeaf64272a560f21d7dc7e48b4451c8387b17bb37dbc19e079d5671636095d312e9f62e3c4309f97e5047822ec0ceae4538;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f09754abd07c6359e10727ae5150076c8466da36fd6beac778d4e3c0e8b5e94554c89180aff5ac2619f87bbea89a2ebbea962e4620ece7e44892909f80442101898f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fe20e6387b9c2246435f54d048b7cad84340d1d91bbd3c741b6c08580c0ad8c5b3337e5da18d131376187f4a6727a4431291c57c9014e0ee5e965da317e26cd3723;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e97b8393e96d15e762f17f66fd54a5610d13e124dbcaa8eb95258bebe014eeb0ceaf7c61fb2636d5f31251ab564784ce1a2491915b77c7bda1eb1e61ada0f360fde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48e91101af40365058b90337e09ad86ddd9a27050d7cf55fedf6c9e5636f7007f941a07bad5b59cc6e3826200f83080584b0949424a532d53f9a038010c49b5c7610;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2dd9aafd645d6b629c9ae7a620cdc88b13851ce614132384407cc581d8d4f481336dd77f15e4b04a393b243e5d7ad8690fc75253c0d9d512a25b8d26c1c059e6437;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c98704727b687d1786ea98dd6881b874a187b4cdaf691245c5bb73e495f6b15125e141b1566469e459fe3a7f04f9421410fcbaa145e79b9d1ea0d8685f27130d87d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e136be93171e0cca74a81b32af9cdbdcbe89248abe611412f330ba044e011bb7c4c84f68c97171c92cb4aca03b00763892de14ac5d23b52d528d5fc589298a6ff2a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce819821de9253dd432cf9b12b3b64b59fd1fc7715c0f1856ee720ae169aeff837f1c53912f5b6d11e305be4453d11380bc3ba711b8793c27b23c2ab477efd1077b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cd2ae746ada7114a5128a31656c9ed9dd6b37c7be78d72b08f3ed04aed174a31fda91fd9a96b13ef4d48d250f8afdd4fc0535badf73496be8c127f91fac2eca380;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6208d66ed4bece189eba68ec2d9aa31795d5e346330dc6b9017175b8a1cdf7305709954dd8f9eed30430337a72c721edb026ea9842a2cccf003e7fe58665f942f765;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9db2e97d9c38d127003d446cf36900dfead0a3e7c538131164f6ce5057b429b10be8f22767c78a20564b66d264a922846288b9bab7481898cae9ca16fbfa2779423;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f624b5664f7ca8457a8076f1388e9508caf6fbebce4d8d8cb443799294e1a02897ae86c7b0c84ce96eb9fcabf2864a660e6586e8a30a2703e82100bf805ddf54273;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49c363a8a0c2ad70cad8d39d41b8c346f79632ea00bd79b2b77b0fe93608c2122f8ee858ac764aad4b67d55f811aaf3243f93e5b9fb88eac1a9ab9adc24243637fd6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135f7924dac71e2f4995ca7f02d2b5dba4c176c28b7325b39cfbefe777695b3b47cdd90ac4d9b7e02fd988ab306cd3b45f89a37a357ba3b1ee3dbeb14b8b58bba75ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1870592df502e57dc1aaaccee0b02812874e12625ee60e6b5c37cb937334656d9922f487835931abcf7b7cbeaf3a91638c2f6db8dc433de3153f1b9ac3edbdeb07d9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae607497cfb93e5006296828cb87d3073217c84e3d1f72a1d775602abe02765ef2c3aa7c26efe3ffee6b07bb6227521698c5de9de8bcadf5b0a85c7598061a72515f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa22f2396153c88b064f4d71dc6d78d1d3b6d2eca591db80d1c329ec08dec54871356a83d86614023b50dbac7f4b5097a8cc7d48e987a9be574177ffabc3ef8f4636;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc3531f1a500574bbf00529ad5c3165796d24b3dc7c40b9adcadf72ee951ba54dbdc907dad185756e28f9dc34062e755af2e65fa0c6a981c078041401b10f5220b1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b668724b3e2137e196190ce9e10ac5f5c75ab117efc30aff4068efda41889304cfe75ea2c6249a4ae1d3ccf8eb888466c242e891eac180c5c203144fb7a4a947eccf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1202af5c1a96bb784ae50f4595f3917ba44bf58d1860e96ece48122ba5c61f822113adbe36a299eb61a7a63ee3bb7b0f30539d4db0d36a805195754bd0492df0398e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bed280be86a1ed68d0240ff6160bd9cca604934024a957d392d66d8839a4e4a759031af4837dd56527f9931f5d6adec408ed56fcdf037053985d538282063f9526f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79304d5f38e57e09fa68c64fc4b858e46de0ac978b3ba1e6085e0fce63f461ab8f2090856ffff2ee42987fe6a9fef7bc5e43c7a519da8daab027d961a50bdf993ae5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b5b1e895f0b2a5f53c0e9f11e81eb5da6c7b4fd415fc0e8832ecddf13bd25dc0b354c1875aa3c900c2504a43b13e1f82ae8afffc76dd8421ef0a9f3adf12729980f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121f3af805b95b7a8dc0b52693907b760768cb91213e06e9f17b21e83d2d323837af5dd1cc6d24bf4eebf19f809b16898482b23857bc00d134742899c2af352486368;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3b521e1e4b23dfb80148e8cd6ceb5d7cb9f37dd5702c8e3c0c0b0cfbdd78634d27d06ac7395b7d5de02afe36e9328e3252f62bad8cab813c7057806d0ad4c3e606b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d6ed68c73fa05cc021e405c395d3e30b44a6f611ffd8b24f7e5c4de6c98c86d9161387f567e7406a3d90eca9d4fb6cd97b8167a39d25d174bd20c280bac482b66a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4e4a5a7248d26b600dfe9ccc410e82f2d02e77a21e9604c08fb564d34419bb9db6f357c9a3b9cb9c7cf49198e59427abf8268e802038cd5306e8e8e96985352fcd9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h495d8993532fa85abac3e46a6bd540ee3837b1031d362a57044ceb30ca03c72c00aa55335229fe3dd1c469e7d6f183dc5920f2b95789ed262545a4bcaf1bfec38b5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1792aa4f9f157e4f91de8ae6fbb832708a82281dab83f42fed6a589a9bfdc8beb5b22bcfd0b2331adaa32c8bc564be7b04a27231840504000af5fbd5ab9952b33224d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1785e32dd4a88e50cb26730e97053021343620cd4ea48edc524d54ef89a141a61d5820515cc7cbdbff91ea08a380fe32fd7ab06e41016666bbb92d93154ceb7d9275f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110874973b0e787915728cf893c2cbf62b93d444f2364d19e5cb705ac7217e4b38dd0cbf062d2d4b6ffb5165922f0df574ded7a85f389f4a346a7cfb20fe59c0b1fab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h521c287efe7dfba98131bf2f0199782bff030a4c428f6271fac84ccf4e00b222d16214b2b489b0f9b6e036206f50b76b06c1e0d4d5ab420ccc5ce4e2fda1ba0650db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb23d079472fa9aff8112ed307b5cc2b427efcb4199be5a59fe18f977cbe49f81c9ed8198d8b544b6aa5266396c428a305f351cc8371e2a731f79ecb43539a53cc539;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h503cf7004c0f2fd4a4d2a206d7b6fc1b7aabb8a1f279f3e5c922731e64da8797e7076ef161954cbd4ab2d6ac7d1c863a5137f5b7ad43430a20cefbdaf61a50018782;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd7471ddee2643a32c2824819172e56b9ae900a5a46528ea8c2c0d558e214d6c2c30d3cb36e95e08fb875084adf851b84324999aa93ee325e4edc5b391948eb8e028;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had5fa44e64fcf0dd3982e6a6bcd19bf4daef54d577a95389f94c9b044d3f6798d0804faa4ed8f101c9eb51d9700822c5e2d1a0cf6f112bbeac774318008c6ee1b543;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68c4556333e0695902b85c6e892a0d8fb8b70d3236451c1d71a7ecc4df4fa538925b18c6c3b370e0f2db70f06b468ea2eece90987c82a57d629cd8dd1052b1e02226;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1318b8225a760395a8b290afa260150ae94ba83f3c2aec90f04cfbc5556ba9eed9d1b2930f404dde27ccd771a7482acfe1fafa66007aa98d91d72a8e2024508060856;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d0af8100ada8e1b6986e4bf82fdc71af2b23f486c3d846cf20ce30bd2c29a4445922bf75020f180a68c371773b04bf8af140b207d60ac2b76a40392df18a982795b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f663dba1aad274ca01ca0bcc44474eb86c50de78257a80112b966ced64ac39d7b45cdf06a66937d021808eeb968f48b82f8f1fbe18d14816f8bfe99114728a83d635;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1613d516425e99e9cea8a6e1807f56ee9ff94b0be6c55b5c447be79ad9f997bf10ba2dafd6f1979bb13a5fd5d63585af8c3a69f7bacd95fa3f97a3c7faf181116e49;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73992796cd57a30bb9fc57d1a6e83c245e7ceb3baee568ed83ea7ba0221961e1134fa6855d95198f5b3bf708b121664c2522fbb98a189e32dd7691e1b0910f1453f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5c8869e58d7fd65032a359cad38e0252eb64e4cf7e20221cd4829128f439141fa3e507c407006aa8332526d2696de307ed3839bdd4b7c37c3aec88c28578e521f7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154d919d556c3d2a8071e03823bc86011926227574efa319ee5ebfe09e17ceeac1c7db1daff77f202ad247de5f4cbee876f5b9067ad627f33176700adaf2146fabd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0e516240dadc6df2ee321888950f5515c595495c74350797be4ca8426009f41411eb6fea1224c0b3cffe5fb4ee5fb389dc267b8ad930870183437d27a16012f8953;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee09d35a315d4e2dc8d37501ec6ef97b92618fc2715720bd369fae45ac10ef4c4bf8611d1859c7191ce035823298a70cafd9ff98d6bd297bac293ffe8ecc1d3d5685;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha54b175700bba05306634d0486a4adb7439151252c68abaa3a9da23670b14023b0afc8fd93080155769bd6a40250c1579b08eb5c80513dc6e91b9c4e3b793e0c9921;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8db424847f51e5aae3a40e56c6955065351aafd836c2b92c4b0ab2d402dab9c0ed428726a0f4d466762e604a1bd373efb35a0973e7b8191f38b7fd1cca6523941830;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha39aa867c774e7e33e90d6f3cbf91e53ff4058362fcbe9a8a6a7363f8c40ced175097b07250ba64e795a00ef33267007a82ab0e5a6bc84780e2d125a39498c79ab36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da3a3d19fb25c8c707aa59aea135a60523f7d4f38e4e6667998a79d907ced6629b075b5a538b9d7d91bdcdd936d29a1d47fa0b418784955985d5d91b2ddd1a1d2991;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f4f092736526daeaed8be4152b1ebe986263c557c453a9c03533420e56c145df0d9b12477df7351d799b5e30ac0277b1d2f989ab814c0518fdc803733b45173d5e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db4a537024792efbab76e6301bf7d771a96493b9ad91cdfcb5b616d73cb07943e74e28dd42e75515608ef50bc45a2dca9be922cb69e88a5c4a009ec71245fed4bf75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad00ae5d4fe69a572b9306d846a5521dc977badc4bdb66b3af6ac7dfa08d7d88f97d99077040527826b6d39daec19fbe1ea87ae916fe9c53a053c381407f3c21f0c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfa6c1f065ffe57911b101574666372eaaa2a5b9314115494f4fcfda66790f5eb3b0d8364135300686756919d7a4a324805a896de1910510ae4a532dc52ddbd00d9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131c733ba2ff79adf40f5d3cba79e4c8f5cd84d2ef1b87eaa5982b3a5ff486ec816c2b3a222d9e5b04458bafcadca246377f7ac2de91d4395ef73fc9ed305b43c436f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d66a8e4b645d5378734e2a527fb08654370403aa4592fc5c67f32b12420ab74ba4d18adfee9057259d92d2137e32d509df8ded6827866773e449586e850e1025723;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2ac8d0f7e77d52f07a6947b7e6b5a6c9e16ec1845529f7e8091446ec3d684b5257a8abc1cd44e4ecc4c4e3a2ce56bf2471a4dd00a80af2e5fa5da5a72af150bf603;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d374edadcc519fe78ff6947f1951eacb975488f7686488f6d116ff571359d1ef50bb4dadc2b9af946fce990045b10b177c0300a209a48f8e583f5d7d82d27885c1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53b8641a3ef6d81c8301e235b17223044214830d158c60339999284430199519e57b5905bbcb6a4d9d6ffb702b7e97d68e812b6bb7442b58cc5963f0e269b71c7bb0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a258c9817aec5eacdd2f5a4ba9ef2c6d8b88cc0347b1b7ec081a7882c64670199773038d561a8a0af98cf148e0c7bb885826b96da69625d8fd09a3896958fb5f005;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b9745f5d25ac84edbd2cffb2f41c3b8804edd137ab3ca00e6a1f1d8d88f0ae19405630c2417469121ce0b000b1a7bec176fbad15b68aeda47a5685c37ff9ce00a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0914f5a8cfa3a3de21bf459853ab5cbfeeeb69a4ca3a0e920c045e92fa2fa5ede588766611253461e43753491857f7578086756e746d2344ecca07c6d29db660570;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1deea8d500a49b7836fe9ff7beceef647b0375fdf8360f07927e6f129a7b6205410cb1a4e9a0e23ecb48111413210be8d3b9fcd20e761f598946389aeaf0e5b4c1c05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75eca23e3a2ca9075b0874ca12eed76040329e4142bc9dff2d78376e4163b67c1a24a2f9596ff308c1cad5edfed0fe28e2377ea86b6c640c77001159d7c1a8e5d53d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3d2ca511d02283fa8b20239bdc909b4a09982d454b83b386e60376091214fab027e6b33786f7d8c720e29494745c92466544ce4c7fe68a6881c43a0862c4715954;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6a33ea2340f08d7b2a6748cdfe6c82797386a13228fda2879f5a463789cf58a94df11d9b575b082c17d63f99f477c7954ea557d5ec9ececea1576f938283230dd0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1dabfb309a1c48a72c1170832f2dabe74d03733928a82a04541482be10c930578aa642dc3cc6e67f48ebdbabc5ce85510a9b588d3da6b6d1fcbec369c0ae6f53101;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c44037e95345c14374932f9b123edaa011f17f522b207e9820841a0e48ede2d2c1fdc451a41da959e905a0dbb72f1529e2222815f97421d7e146155b3b53ac3804fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e86b893169c27f64dc109dd75bb19d1d6c4102a2345a3311b77a1da3fe1b427f0823ec1a00d96347fff979f3ab3081a1d279911ca1594a12c4cb086bcaabcc82dceb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edff78d8cb3a5f4d3c011412a8205322cb6d295e48fb398bd8ad02436400fabe0d0db1d0bec4ecb7ea2da614ce934362d6cdf6a35fb1c0529edfe7c3709c1f6c5939;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70b89147904634c07e1dba921d3c8d1886b57a19093efb37d848dc5b2141dc11374777b6488edc718897617e41e049dddac24822e77c2af491e61ed6b395f1908c00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108c90ea935273e090f611e897037e16d47c0ab00bf26261d7b94092b0161c54f31c13faf160b2cd2ebea27fadb0dcef67b5c3f79de1d6dcaab0fac58ce0dea889f1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e49e72fa7aeb17ae51796fd4d1b06da532e04a81df8f7fb1d6d6e8e21403f88ea96e0ed678871c423d88b4377b5a354bbb86010020f70547961f176bfbd58401439;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e81008a9f7c46df1d6d35031b683b5d8815040308b59537b582c02e86a84aa41c55308a84e0b5b1f6ca3a59f972d03dd0b4f6dc0e1fdffcd47d8882772cc91699ddd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4b6c8b07711c5d0d7195f25ef022812704e2aae8d03204d6be759dacb7140b3e617f8992bca98c38e31c984979d53750e863d28c7deeb855453bba2809603ca7362;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10dd34e1a88a3f10afa11831a09fc592afbba3ab0f491ea489f835bc2336b7a32be2b64b094623ba4cf5625c2297230281e01cdd40cd4481f87927eaadf4fd07cefff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h506bc21d3decdadcb2731b7dff85b4bde13a25f2ccb2ac66f8828dcac7cd88da885f62f05876185ed91c62656933950f3cc33e07790e4d7103d09101a3a717a01c18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c5351a56546fe0d3e6d562664ee4a77b07818e59691a63cc43ffe2c6b41f86410e43eee4364715907b203edb242a8453c98ea45486403f63131a29c8b5e5f153b8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1226e8a6ebf4a51215a2d709c8dfdef1d0e368a5d89bac6a1ebe47ee862b504badb7662716d2bb0e149eade26447fc47ea5ed5ec8fd4c3bfe1d0a06f4516a66790cf3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118150117460e7a46f5154087b8f8f035dd2cc648c52f54afa4f65e80f045c80bf8bd7745ee9030cc27d35055dfd37a38af9d5d949e020eb10599e44a04a4a41fd9f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1838d1302f7551bb5321bf0213743b2eb3cc402c3566be503306023e90bfcd2a29db35367af086540003e0d3459a14594fe8ac3fc26a35f38fd3e1b0d6dbafb81c9ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6d5e39c51f1032ed504ddeae2a8e65776610047d59f0801a5c89426ebeb308f6dd6229c2465967fa374f5bc43b7b5f748958d5f6c0126ac478ff89ca85ac7c55ceb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1394ec5a86813dc2a0cf5507eac9ee650d53b78a485939c275bdd19ae30ebb5c018207087d67bcb93807c2b1426394a2ccc653284dd422eb4cc3bbfb1b925b7ce759f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b7083b923495aab65615d773373554189ab74c2d3b0bc7bd70672b4141ee297149011f928233757d4cc88e839592377242262a24b2f54472b3df0eff4f06503aaff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170f0e4e22bc15fe9732c8e63288b9e6bdb4d8ab23c219804e0ffafd7f7accd2697da2dca69e98a11f147f8891d2fd1a286f88079b0fb69ebd7573436fd45e0b6fb6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f03ed97f98bba32f0dc38b745ae397f5a38a42068c5500a343c008741742b7fe96d9b51083e1178c5c0a663a1958877c4c6b54a0cc3cf7fb177265ca99d8a8f0536;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d03d2404d8988514a60440b7ca68e71b6d991f4428a46c4802bee132d29d46b5a24182d0cdee05edff20dd1931530dd4ffda28a9c2dee3644d1489e9f3f234f30d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ebad3cbebc30e6332474e3409486f2858814bd7e561d93b37c55809a69fd5cd2b8126f6374577057ee2496b010852a6fd27fbd4df62182358e28cbe9ea7b2ccb4fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46de784771dafa808b5f5bbdbdbef74a4b3a50e7993e03932e6ccfd9baa9e83be1486385db5b9dace544f1b522b389f2019564edd01af67af0aa369f3894d47d0896;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3af217b683fffba314c2060c788256dc5b9853a9fb5318135f407b785d6c849e9ae12e95bce17d670d5198dd17e8cd39bfa458eac6e3dce7a8b71feb18fd76f38d59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6cd241a81cfa7f50143b7a8a325dd9a288d27665bf748e5fd565b8eb31658cfe9b25d25979975caa38177b493c0908cef1185f368672091c71ed5b91a9d494ff216;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6dbf798dd2a21ddd0e227f92af9c5b35b8d5d7ea951f5fdab863e0fc67862793decf9f2819edf959a1f12c42a9ccd09d3965932bb43a37542a288eb536714e30075;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae2cac91edf2cbc5ecc9770da2af62202e3b49240d2f645aa296ed1d8b4b48577dab5e12ac8a2985c06a149833f24a9c1cb389ab2630f9957772c49543fdcf6c531f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40689db1f93836cbd9a953aa73f72636c397e7cd2e8e7f9b91c104a99a4925b0d4d559c1ef9d27fb3c9ecc78ee8c8e38a2d3abf6e85f2e43de0926698c3a06a6bd52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h633af832342fc50a4fa787bff547bbd004bb0b6e8570c00e8c24efaa40530a4fe1ae91de1443e2203d129f56fa644dee0c3460409373bb9cd454c00a11534c3fe9f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha595a62e49d42c8aed171e5fbf3ef8e95a0758a018c583a3186ecb5ce15e81e9733c8e1aff9192d7df841a2f0008f3dd50006cc2aa311a7df4cdbd21a66b91fed7bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1657230320aa70f9bb7a7ee19e740116cfaf1b88acb23c6a4e04eba3eb8faa3d076f112b10ececf56eea9151105362495eb4037d192b987f8b7796fc0e4f8d22c0135;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8a5d7d556e77b72723f12ddc5c514de3cfa23923d39005f6ba6881c1e29c0a4dfadb2d64d4647424bb9f0f3ada4936217fa80af63a516aaf71e5f9c520a1caddfc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he208331211bca7ee9a52320891e205694000044aff626a29b352bd63acac164316800bc9cbde128e5b2ac992de3662545c0635253de7275dc81f92dd13b542761658;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3944a6f48329ab0297ba098d331a6b8b8679b07d35d2c8ea28686be603930d2c62f667b67a7491ca6806493aa7b9ab5c35db7233fcf5ca3ab140abcf98a2cc1a5f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16faea7be7a85b5429e7d640be4ab86e4cdebf5db79bbc6308da39dcc21bf62b4285c31249a61502da6b29b3ba4f9c6be82dae8d8dff444790b9458c8b17980cb682e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137bfebf65041da10037be1c505a936354e575be5fc5e07cf48f88ab942c83b3424428d13d18c14d12997aa0cd71cd6f59f9888d789414210624468bad6d7df61518b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc55aa62375234783b18a111b4306cf332e5185d927abed073fae682df1441d612c35178bb1616b6eee656aef5a16867ab4056728b9a61bf823c8afd81e7f2f2c6bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14232d4ff02b1e6d817a9e98d9027961ebbbdcbe081e325a7b179be663d692ee4d6a07a94e74b393f34b3c82022b0e0b9c6895c307e9dd7c5526df718b54b3818b682;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1763a475cf144fd100563630e3d4a09162371b7ca8a4bd10be413c9cf8df056eddce15c22514f2ddb8f1762d4516aeea20f8b145232bc2a4fd85cc9636b875d4edc34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31a2422e445a88f208652280e16c76d997b56496f7dd27789a471ac36885dabc23d788413ef8e13210c6a4e5abe94c8b0af109690343a7aed5bc71def298c986a998;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d1d4655c0cbfc7606bdebcb46e342d3ad1bdc02dfd2dad3444dd8901fb3c32c6539165b69b3285f49de51e137fe51ed858a429b05ec63934abeda800e9535403182;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c42625136d5f7e006d4bd1c3e83593f85f31a02d004269b0f5b029ba8d40d1ef3fa4ecd9f6068fefb607afad8ebcfc2703f54d806ccc1691b4be3419d23fd355af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13525e2703a4fea86d0ffd4fe91671acff1a13fc8ecacdfd920d72e20e37477d716ff88182965d6a00f502ee88fbb57ec530f6e322230f1e41f8da3ea20026776ce09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61cf17f8c627a6e387985035ea4747a66e47304804442acc9395ae5e157ea4fbaf5e565145deba329bbe6f2e4eef43d9c3117f55f00b8993d8dc6e69f0d53b6177f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8c26fa8354695a637368c18c2fcd288fd7b52780da848bcc3d5815192b364adeb63343de560f51e456d5984c228ec6d41cf6c7df072944ec87b7c0d491248829035;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb373099eee4bfd7fcd62864c6411bdebf76c9f30439b33ba08e974a5a0c4c038843592aa506b06be94ddd5acaed096b7668e28cfc6284c444877abcae0fe3a363e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf63c9ef5386195305356ec0aa26b751469a98a1a62c2afcd114cd5b2b6fcd31894c5ca614cce7acae2cad3abaea5dc7f5b82d75ff0babdf97e055231e2e80158ac15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a305405642895a3eac5c10ce22db558d24a35efd0feff86dc31756be8bb6b75f43e8cc89a21ca1ca89b4ede70772901c34a85ff1bd82e6f3db6a811eb4fda488360;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3c4f9a8c9cf9d7ac6e7d14e57d8dbecb210ab88e189c94ebc7789e8d77b6c44d7a09d512cb637c89137077a047c2673317c72dc0e228e83b4bafde489a5734b4838;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd05f4e4bf7e6f69c001ec8c1c69269940e3542a5a62d07f38b8d0097c355d55b60181abf82836f169656ae8dc6a7b5fca70780f4c96259db6180555a34e5a98ccfba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f25d7cab19e21df8b22de0c0730d52cd66d2298b65b0e9578e2570b3a11503c850d51224f5cbbd422d85e211139878cf06cc1f4fc77ad4826a759118e1d4359f4efe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9950668e6b31320c9bbb386f53e74b8e4c8654d46b0ffeb8e6f62af424ccb94ea97398c7f8307d226398600062cba3d0762db9997e91b4e25128e144b1b4769fc81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf87dde196d5dcc586570b20020e1fafb276dd1763173cee0281ddce31663f62134ec5ce8ff95f1d335e0fbe727b74fb9107f38cf3a8cb3c0d0e76f5384654856be00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8f4f4fbeb05d4cc7e111d07689c5d041d128bc93c704cfe371ac4aba0a1d28dcd440929c5720e9f76f96f90ea450bce2288546be813c91487f7ef8248a8f4a37809;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4660cba51eea762b7c85b070b0b35eefa4ee7faae3b7b8eff31896ea5456f4406303882b965b13085edc600288730ef7053812cda9e4dc71e9aed59c13d3ccf72c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce4820c2fe007245e3f8c9246bb300c11f7cd15a313a14d7c5d132b1bff93d50ac9d32c3e8e85e451ee19404bb9acbbfaf6a9361b1eb4befdaf203c319be8bf088ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156d50dd9988d9ef4c9df4f35785fed15af05f6755c4508a623b7e1cb151a589e4ebddf770539768d1c7379113d1f3eb630fcd4ec216ffccaa08f0314e6f4fd435345;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139700c9267294553e4eb87a7c06d817cb601ec181e7db5b79ecfbab30049ca502f864d9eb70fc17d3cea3f2116e864962aa71907dae31fe1e51e314862716eb33b14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e8e15f960353fdbd55fa7e04aa503223632ead207b259998d33f5a66f92baea0d5d14a5b64501b5e95ff1c04c369807e6d3f54560a5b25281d13c7a016621966ed5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc7f00e22a17e526ae6f83353ccd1302d08f145f7eed9d01f8a914650513585588fe77c921af130677bcb02a877676b0a0313d55bbac496212f9b7c2ef2d2aa95860;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1299bbab1c169d478ac74d150f73858c2e1f5b37c1835cc8f1037caca17aa4df449e5be5272f0218e3df9decf1f1a3a131060f264349027df742ba92b4e15ed9ff171;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156eadf41917590f40e300c0b39a85be1ef6fad2dc60a1f407f2615773265501f0b9209ddd3ac5de8440ac94c96e24f2a0d99e599b43e38c76fbe43d206be79166993;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36c9747092ed5b2b9ef3d0ee9ff9eb43a2bb65aef62085d29c035b4a5fa9035fd23c15c80efd2f110df1a1ba2ae02178ced5a79f0de440d5dd8609ff128dc446f09e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc61190cbe51139589f8bd289433408a4484076f55189f70a89edc4e70b0c15ecbd766d15724b64c30e8bf23bdf2de90f0fa8c3db32aa572ebf13745a6a3436a73257;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32a140e1582a2ee404055530f6f4d94d66ad763c3f4958a621941d7dfd87a2c7892c9c51e6d3ba6cb5eb1ec151a59839f1c4975f357335fb6d22dfe41119eef9fdcf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3ef5c1d614e5f36bb299cb6995c9337d80f9f37821708268a561111531c4bbd1f8170746d5ed5cf91a9562f6012be178abc7b2dfe8ee5c931d20a015929f7daf951;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1591a0b64305a5a0f3aeb185f05ab5388bbf7dfe9b42200ac0681e77e904ae8b56f83a11ea6556051e14d4f804b9323b9ebd158b5fc32cce8e117d7736243f9b97e10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1191605f9c55b949d6ff299048309b15b1d919a0aba3c6a634f40785b35559ecb87a9fc3b531a2415e0f87d75d0029f67bc7c83a9223a187bd7c057593cee3c1bd3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4a5bcecc10d23cddce3ee4d39a09ec9dcf63481cdc74404b434871f5ba0c15b959e76f7db3e7884ea494deb232dd90eeda84273093d88de27d756b1dd6b01d7bdf6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110e09422e32f8d7aa36ecf5173b5c262ec3687eb32f8042c1dfd490c9a862a1210d4fd2559b449855f392e2f252160a91ffbe8cdbf7dc5d0ba641c908f40b4ae1e0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bda75ce52feaf8531442edb88ace4a2c67324b43b4f691e4651cd43f1aabd107f9c87a97edcb69130c0d666a3790a087e8e6d40c34ad05aeeda6b57ad05a7c2e94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9e4002b0df54ecf8f558b93804b9b4d59104b79361bd9cc569c84a23c5d5656c358fcb16c508071b2cb0f6ddabe0231823a67e0f074189c63cef95372ca62357ae2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b8f1d63af33b68ad0e240b03f749dec2d6cfa2c7e8b0e99032f4c2d6582c97b7c6bb11c973000974724b92aa09270a6b0aae6401a798e405cd0de860320e9163ec4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h835799ade61bc6068cf1a396783d542a33e77fabd3f39f297fc8a5196a80db7db4c93bc8d0e242eeb4648f6e7124629df0ca7c379595e1a28731be3e9fdfb6a3c493;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80a75d4ac1f149f3487758e07986c34f39bf2cd33e4c8e47ce69b3da29d4cd7efd93652f1ebcede8b1a499a85b019717bc003f3f6027e8571b71ba3550a022843df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he240a48ea6b8e0576d4eceea2a32166533d99a13a7ed5b6f5e90a62692709179ab3a0ffe7d0a3ed68f08da9269bf248373605b3c5b5d197ca01392f91e12473605fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c5c185f35126e913a637b6d0e17977fa884f89028d09d069099428c23a3e7a979bfcbce8002d4e55b3ebce1e94f3bdb94dffe9336033299ff11984e56977a5691b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fd16e12b491204a3b2b02c94c3c7d46c1101beccf8269e9654975467468fecc5fa0b33bd4f907a26d7cf280d434302c5a4b05870031fc775b82d695f8201132f8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2adf71756b743761455e6311511844244d345ed2537dda700ebaeb00e90ca0d32e73b07a83746947da82bec178eb7a492a9ba7da075ebb6b25ee517e9ca64d00c7f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170855b6ad7e71f96740e26f6f64fbc5c514104a71d4ef2718373ebe3bebd907e51880b34fa4fd646f885684987dcda98262702adc85643b3a2ce779f97463c172255;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14dc61c19e86330508c9885f62e33d7e7f44a31dad94096ae4e4a452f945e6ed3619726a5b7b4664fa52d7b1bd400d26f2061a47817ab2ed58768629849f9ef0f5cde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e35aa1db3b89c1b765e9aa0ea8144f9bd7a09e0c893ad02db3b11cf3675dc885fdb4f807cc99405bf95ec1c86e118d06c67c370a75df6d9981f818b66dfd3737aebc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd588e0a9318b8aece4a237fb157d34f3beeb1a0645fd811675ac0a5e888b6b93d8ec52896f14a8ef82b6c77551c56582caba6179792b737a34cfb334984c21541ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd6cd53bb5e8cd1b94203532d3a37a18ba17a384f41761c5022e67665e7434e4972c5d5bb3a6d2df3ac3dee9a57adfa5974180a74358f6563cfa945afcddd6af6176;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84bdc452ed890f96c3251c3faef6d4dd2878273939095c6166816f32c0ebddefe94dffb317eb41b6d7c2fb12e46b9802ae6f9477e73d997e3698b692500eaea4f56a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19bf83f2e951117e6d3711527ea75cd9cc8f21940ecb42b8ed1eae3434855c26b54dc5d93fce586513bcccd5336226538b7f47566413f4db2dd43292d39061d09a0dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e03ed64c9ee02ad84b2d88678afe563960ad9eefe6f98741cbfd0526790aae11d90f5a06af37119a9a9a5e2ca2b1a8334996bdde7d8f2aa5575203a272d776656a38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a225d4231e29544ab6516fd537be1df7f6dcb83026051545523a75e374cc79a44968755767be2de6b4cfe8cf5d04547bec7214f3d44bad330b3f5fafe5653676c110;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11295e5b18a68d6392052c35feab841171f86d0124f4854b6b75b9fa4a8328d8a6562332a1bb2bc68107c0539c96e887defbd7c30252c8c94c457c19e1dccae462d16;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h990c27aba7a1548eff051d2cac705c4d822b776cc53d97d010afc72a9659862bc67ffb543ad124aa2d2d782d2f76c25a10f5e2508baed71a33501590ec9555db2c53;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac6d1114e6c861c5e55a53dc9ab4d13cba0167e7e024b76e570047d0e20cd23396044a72f72861af0fba2ab9ad90a40aef5a29e93a31d234c943b2f0c2d46a2fe9a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c2429437452d45f97ae42119cc719f7181d4edd976287ab82c0228ca8fd7280057e8ed5d9dde2b5950506b7851a2bc6372fe9252cf7e29b5868c306829d6126f64e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf580dac7f371851ad02bd05de51453c6fca568eaebef77a8db11c448b6186dd5becf76433d0081e4aa01d5008a9402bb87f131c04e61c58fa156ac57792b5ac9299;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1304dc11e2281884595dc2694c238ddbf96e77c256eee1e6c0d4f9b76508adf0f8a1c9e1054c3d6ada633b085733be797c829992a7e9e1496e5345f67d842f81e2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc53862a1ec8436951956c1b49dca7b0068191aee741def1d67cd25382d653595f1eba30da1a2f8a9f6d99ae8b866f3eb372b5a977c272a7600bcfe052911891d00de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3d9f810fd981e1226fde048df6e5bd5d288ba0ac1efdd56904325d7bb2c2577efaa43a38b015d1f27ce6a05da0c17d8be2ef0901bad95943cbd309a962b268cf0a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c7a88d39f7ca5f6fce0e88c991975c27c263fef3c7c984746e2e3f9056bfd0fa3b8adda132e365ed4147c18001785a0b8e57bdfe962315b8917b95525de04dd5293;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc795874f3770699b11a216b02cea12232106f322bbf8a8d2a528efe26fd50bbe3f6cf65862517001e032edf2b3332b51d2317519906e3ed68fd30e821c222f6751c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98c0e63ff8ae912bf3bc69101f7e09df7480a2ea41104e969bb87c89e13b53f75e3c2fa3fbc759fc90d5962a5d5a156e7b0bc9e9a4718d46dea923e72ac1dc735337;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5ca0c5d93c2dd931b19760159952d277274f18969f4786858baf6d052ada567dc6131e6146ee432a3600fe1cd257bf9295e678d2f3e08e64cb5c847fdb3eb1c202e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179dcdff9c905e51b06580660e592027062de9195116af9e6a6876c61993fdfadd4d230848f162b49a8d5913a87e528c5313d7e101c466e91af0aaf17c7db8c42ab3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54d20f480496a4d739757ac93ab5a977da41fbe7e5ed4cb22fdf1bbbbd94021eb5a8c352ac783d29057577627654323bdad1cc4fecdd265046892510e48a41dc9a62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e33bf4fb45e9ff1b6b60efd8437578ed57363b1a9a056ad75bd216d674ad645928340872d02dc4a46c2f950ed9873fc7bba671a7c51530d4568ae61e698aabb56b14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4f5656bc286d338c0b907feecab53c659cd3e1daf2396da97bd9922505215bea473fe2254c96236329815c7f788d53553294b2ce63c6b53762b07c1840982a4ce8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cde60517ba7fa6905a654ac934c5a932db7f82362b9f99aa13ce6f968c5a42ead050319a90b413d0dbbd091431ce2d6372ea6f9de4f66482b07092b8b667f227ea9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cfdf05b8321e58ec6eee67747ba11b7f9b173e40baae9bbee7aff7c918022506cbfd89cf83b4de20bf9236267e040f97a6b29e5e7f43c37f1fdbd7ee2e4443d2424;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143f3214496ff0f22c917b6a36fb29f6003668ddab80d5eceb05334912d348c2eb1c30d3c7f2b6d186a35cd2f8862f71f2e6cf0b2a98b65e9173cef7895dad052fcca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168b3913021109a66e0208b69ead8980f6012df1a0a89a10a511548d4bdfd054f0d52e81b75609cb62ed63775a8b9484832e276df64b783913675d2fed3a21a43f2cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de2f6659391dcd6aa6e5edf3c52866dd00f09dcd616f3e879283bd156c9493a006bb32341feeacae15b6dd724258452bb7a57a4705a666a49ed0d9b92d3ea0419d8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113382f370ad29156ad5d89d144571117657f1c21c681e0565d59b16f6df7e215e7e555fe6cb72795f2266e59830e6536546a5fe0dd432dd0081c6334f1ece289f25c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e6e3551efcc440ec08e8ae6141d8acceae254b76acf79c8f67fedb59d184630708135af2fe4088d437bf335923d903aecf4ee9ef78f4dd0acf87640164799b20f45;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd67f04675be325765e819606e61d6c0d7db9a11125af985423330414f6a1df68db8c8cdcd937bce86b031875e0d70204e7dfd5f124296f7d5e315b033a52e6278ef3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f5e2f0ebdea03adbec04f873242fb8e4ac84ec37fba9b31851accd00d875bceda1578e06661a3f5e53234bd520964bbb1938da28a0de3ec2c022184cb3e3b1dc02b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b204d8b4f973c45e9dd8862b0088a653b1bc521eeb043e2f298757acc728eaa1dbc1ea73732d8fc20c09169ea8f086070cbb722363c8039b93d33800e1eed9a9c34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd43812562076bed1b54b3d879c2e0533fb593efeafacce641270ecae24dc64c130d4cea3b110e0754815722f28b9ea372195452a5f65a311d14d12ad87dfb3f81be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2d5014704f3a015e56e954fe769d88c6bef55df0f708123d20899ecd911593db5b38948c4c482ecf9a23c8bb3a86c194c2c13756362fc3085e68983b1156ce8aab3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49614a0a0acd669b910747c9cb6da1f1b04aa19b32107764ad39e58d27f7509854cb39b0e46863cdd38ad2ac146750c42bd07da8f50993096069ac926fbf6082dbd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176fc714c659c9c641ee138a1e2596fe08637eabbce3494435757859c4d230f30161cf4c63982e31932d6f4dabe6e9ecda43ab816d01c20fdcefbee9018464f87a440;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1092cf0377544617cd0de83dbca08ed9ed947b94a7c85f9ee6d6326e3bd8c2b87873839ce756f4772b66ad9e6ea3a63e7f777ef02c76d25cd31c97272d3d2c8bb8de8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5beb5e5df5a6917a3ab1f550cd43172ceea4532911fb73cc86171ca041bf3e9379c1dfa199f611db704765578ec340ff5f37d6305ca9786d10a9757bced8362e7c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175b6920793581e9531bc66ef8980084ce150b5ff62c5b4169c2fa3fcb279270866a3828ec1966a4343ec93876c5c830dd63865a1816d2cb665dd65cd7df69c2f44ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163e772f5f85e19187b0d7408029b03fba6f2e7a2afc3c5814bda967d13b1532f83b427e0a4f4ae347de1aca5007110f938d5aeb070da0947bf99d605e118ff65eaa7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h619b2d9f3096a9246644675299cde7a203ea95d9b80d37fb12c459de625f0ea875e41109a21db4b461a0e3c6289408b95d256615025e0713db7d8336f30f6c1aa27f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1256cd5b1f1a17168f4f6aba6b8156d645f0b9017dea3f14b4105a46028573ee6d14958e80fd319f2ae521f85aa9378e9aea30e98cd172a53d524fd2d4dd2ce1539e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a7ea6ea5eba09bd33e4d02258926c2743d94fbb704c1f1523bdbba1a1789c88e1aa61244517d71747b730b4c7a8b355376c40fcf8e16ae164ed4bbc20f95b2d94d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfff354c223eb50acdd7feb2c209ce8e512811a7dd9888c03346c81fcbfb5cee8aa89efab95ad5dc7a20c8f683f7c37e772afcd37228ba08237c0c5a23f17f8a2851a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ed615cf622fac7f86e97272b648d2676d5051d7da71f6946382c00a2b3aa630d27ae980d8ee1cae208ae1a95b2fa707c5c3d51cc7e0e618257c9ab7d1834efa6875;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dad4df733d3a8a2abb2215fa6f72d49a153a386a62fa7049f6eda50c85f74d6d26a5817da1ff32fe91f2eb79fdfc0a9fddf5ee0fa31010afaa779094f99fda3e3b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c881fb2b501c5140f2bf54181b8edd53681d4cf1a651f7e2a83126af6e47bae321eb4c410a387a9a86167a32301d4ca9f03b1f180f9eb1fda44f15b7d770eacbb447;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4693791ec61f4631f3c769470e14dec31ce554cbe7ca629a2d062fd342cb823b16e0661015d8c77ce4474f880924a7cee5b968876324646f89b89d5a781b7d3ad6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ca6620fd2b27b5e24ea5ecbcab7296579bbb107093251923b1c19f8447cbe49f58a59f1b10ca472e73a0f65c312d9bef59cef52e0b0f78a80e67c9d1496c92bebc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1153e874e6c6afd41135da1cb1a9ec5dc1a078581527d996aff9bded92bf3ede658a24b7d2740d10204822e7391b0208963e0d2112f8d2817bd962370163dfa1cc7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe0868f7a7f8b15b4156bd1086caa2e5cb4abb3114ddaba045f09335a46396916af4b47fb6bc2418caf1bb43a4738a587b4ca479883c16c5c1a1354c39f299896ddb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc6bab120f1206ee208c1e5151c0f8dd6e621da126371f200774ce7674fc47dfffbba9c8cbca35574506c54a78550e0ddc7ab938b0a8b2b506259bd6a857ac6d1646;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c62c153ad83612fd4de5dbadb06563de0832e5d0685b5ffcceada05423c6540c6d16d4fc73f786d216db69daa5d91664fa3e5f02448309f6e9080bb274ed4356e66d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h246bf547259190ffa30c49cc521403d3676e94eb27dcc97c37766fd3b185dd0cf5850e3157217630ac70ad8d25b924862702e5ec22b304aa68b0a7cec132144c2354;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ba6843d58529c8ea54a74a8e096e1ee30e9b6292046af8551424aa43bca7e6bbd1f0c00464e7f857d52bc109cd31a06c08a802ffcbec1d800bc0acbe79772befbe2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19154ec65cbb2f3266eeecb63ef55e1bdf18a5c555d216877ad1c6ab2989002922cf4b8b23852892a819a68c10e7439439436fd9fb663346a5632f8aba9f3b7be66a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88c495e3ebaf739c293a65cad4e2e2a38512cdc592dedd2d7ac2744956b72eab4da119a4c65ce312e69d3b4802eec3d157b306e3d65e3ac4ec73a187c3328e3156b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e50914c49c03ed5d6f4d67a7bd91947db813cebe0b85cafa2fce6fb188f6f48dadc0498904d0b9ab05907c38ca771ecabf2052dae5b6fe5b0dd5aa7c920fe45b63ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7a6fa7ce3e795d6712105e3a9e3e0bdbb1e24e65f596ba279985d3e072ced1c02cf462aa77d53b8892afa81901a92d66fe36e2646479059d573590eaba79cedb15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25415bcba21a12aa065f513ce47ce36991d54b9ae12285662fffa5119493f4b192df5e950bff7a6c1ccea85981834af79abf099156de19957693971af1e5e321fe96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d7d6f52dc4ffc3119230c1d8bbb10de071c492fc78ece89f5189d886c3a22876d712b8f7e9d363614d7c2080611fc313ea84509ff0605f184ed7924064b4c54a432;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h429d40cf0d4e4c7c1cb659f4828482cdc6d0812ca3d6b4f7692c60b70a6d0f071939967c343f6abd4b229d2597910cc6b3bdcb9888465771146b1cb95954b8b0a2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35f6050eb20b6d94216102d171ff167ad8d75ea2b5bb9ae08e23680ff1c48f4a63052351116fb75600535a76cbaf632b8ec9e4397869054f511c4ea17a79ed13d37c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbbab0eb0aa69b28ea16e2ca1fd9a188fde9580f5b8b5f4ecda9b3c2b327638bd4a0da71d3cd4bb43061521046a0b238f42d8030bf2f833548fd6e5dc95154d4d857;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ab4250443fa1a4e548c2ca1618c27e9653b8d8255c1fcde742020fbc0d52c36e49bafa21c78c41ca1e7f6bb1f1272fbe0a7bd2f2ca53e29fc1495f668a249c71f91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6db21f664efb8cd2c82af47ca4a77425f7db283629db3eedf8fadb69edc22eaa8ddc71c9fd16fd90814a2aaec4daf09e2eece2d78e76daeacf7f875e984ebf4b4646;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bacc5ad5acbb776692021f17f47b2b8d85cafe8f81fa42265491bc3b4e2232c45ab3367c0a32f2bba5a44a60cdf8aa4e30e032b7292a1d54279f90de437ef7034142;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbab2a166e7ca8a6cc420a5c0a55dce2c446ccc8664134fa9dd58f8339cc00c605a1fb763bf74c63c782b4627e769400365c539980155aa31004c3488e97f3566fb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13342020cdd6eb7b61fd51683721d89519c9f3bef699fafaf7521424d4b3a2346343540c2f5d48f5f38164389038c6d36cab7f167b27c25f9443f0a02c3028906ab86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c13e43308d4696edf60143258262680b83d4d6103fe7ac64a2d1a6d75067c7969f2a558b683b50c185267d8e2f7c771d18bced9d8b2e18a843e291aab47e9159efa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19444fc88b210c88d0407e739953186f0b6a281c8c3e7ff7ddb5bfb9567aaf8db76000e547c169ff900bd887f6b2823ca1964fdd0d0dc760f4e07656308f8d7964188;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67a03d2f01de019b9a3d57a6ed6881346c50d88c339a6da544c57c7dbddd8767e24469ca3de8da40f1931a6fbe81a5346212a52f48bf668d8ece799adff37450faa7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2123cf2be518f4b6777df6cfa1f4a921473bdb210ff7e851e10b40b26562bf14ae35dee8eae92a0eec7b34c5bc264bb2db2834226e62ca6ded4b1e7a16248eb2e59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb8f3d6055640e305553fb9f347cbd8f0bb908b5926d0e02a844fb68fece4bae6bfdcd4ad0c85b2c0b3010914384c51d07da07b6c2e0ca6782d4d43f9108b83197ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b20ef92ecc8d43621f7154c665b27f290403497807cc4a093692085fc2af49a2ec26cc6ae4161be14c13629449474aaddfa2fb56ba566928c54a933b092450a7c1e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he792ebdee126c0363dbfa130e42ca07f4ed65ca7ce5ae1c065f3c50ca575a28ddd9601159f9c81edfa1c004a68a4836ae1fd7f54bfea830bb7ed6a4665ac6c7837a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he77c7b2135cb77f7c04420b146622d28b47c19cb817d61fc381b1858b32292cadb7b0b4dccb03e0939cc0358442900d354af091a0ea9c8de680a4746c5f1d69bb763;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed44430f9fd985b54d42fc65bf698c86a74ce69d7eaae8046ac6407657d61999e71a5c59c54a87905da39bc53f990f3907ef2bae80f1457f1cd6a3b3a8b57e76f777;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1284352e79371c02a20cdd470e3a8e2547d25d6b4d9b60b0e17eb1e2cc953f34f55157a30100b8f47ef95e6ed3cb30d8f654e474a6ff46edbbb6a1acdaec771718b99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc35b3e3c94a3c363ea9dc27e0efd79dcb85d0efc491d0d49f34e59005cd6b159acc157294bfa55df1f0f6e745e5e7668df1a35b98cc7facbd3668a1b0dcb6d2cbbc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1500ac6513ed67c2d315f42379ef6fbf754ff887ad723f825e44474098e5ded6ee398c066260dbfd77a1b172571068fbb9d11479acb50d933cc3fe190376928e7b2c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa84a0b22ea9745411afb4a24c6bd51fe76873f6de8a0b7f11d29f9c6ef4bfb8239b98c0f687e46c2b29cfeac3a0e1dc645ad32f239d76a8359acf130d4936afe16f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5a43ae9f299c68afc879609a14fdfaea4c879c77dc02fa3c77a471a3690b79109fbe4bb35e3b43a63a5a351025eb2c87f0299f38fbc33feb926284d03d27ce9258f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a71fb24fc7902cc482f54b7aeca452fa23600e90c2b7cf15ab256634b3fe3af7b9de1088ceef42b00d0559589fcb476e31307ef5a30c8cc9efd95e4ee1b9f921568;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c32017debd3f695d2b1e01858d41902dbd12cf0ce2904be1ca54ef94fe0a25eb29132363ca4056d648fae970759d7693658ea0631c33c12fc05bf1f8e00ca0bfcae5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45b3661bf9d86e791fdb5f77fe2b1396429e37da81ea9ea0ea97c981b1de4729d5080193485827762a9a01853c216fc1c7dd929a660fff2df2e69261abcdccc415fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c87c7afd61bf122d4a1c1923659ee5202def26fd32868db2276c70b1389b88f47379af59a81f90e26cca9cef98bb51db19ad94fea19ad413028dafe3a4c55edec1f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he81910a244eb47598682a8ea0aa52aefd73b3bcc3beebd25966ee4f1b4d16b7373488572a2472d7e7ce30a3739932ce2da7455de864cec0de51b371e0773db432011;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f548d2bbdb3b2a34f72774cb5fd71a546147bbeaef25a13c9c0c965a15e313dd20a8d43222619c8870b3e6433a0ed3f8b13fa5cc5491521c3b3343e9b0b6029d0acc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df2757740480a9e411020830d16e87a1bb438a81d3068814f733ef4df8df26c20fdabe610d73a4ed700979a133c5bd9631fc0ee893f048632167e49ad7fde4ec4819;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d3f1aadc3623d25703d55801012238692eab734ca31d5bd26b07f72690ac673922733b6b04ba5c5e3615edf37aebfcc6bc6d9488c55716e8b87971804ca91952605;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h628237b696a1aff8dc0aadf501b6b489f5713d524c526d78c7595365adeddd9b8eb4f11801ba1d78fa77795959a56ddfa699c204a0b93845ce78897a3984d82c02ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7dd79499f91d5223f8d84eb242240592496f988b40740369773a7d327d28c5a28b4f01f3598e581ba221cca4ee22e140415d400727c4f92997c2a2169c2537c1a6b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5244a19d8d905157af0628a4d5744decf9285fb164e9d5ef0fc8d212ea88f705f37eb9639f69dcd5ebcbb9a6c31bbbb5773f89f0fd13c76f616274f91ce6c606772;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121e2a78bd38b0a3c6bd54ee588e3d2db7c13692fee17c002b7bf3521aa2bb041d27d87dc6aaffde8b0eb9ad99d7ad182fbea252ba8cc2ed59a1e0fb9b8845d95d32a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc6c5ca29d277660027c32525cce949dbe6ce55b20d52e5ba618e97e07ae6eba363e1a88e70ba8b196c2be0d33a56f8a9b01f479d721212cc79a00c2cbfeddcc37b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf036d231ab15c7a07517ef8f49bcafeacf096da4cbd5f5d5b13097530d8d440fa42a66ae3510fbb393265e11b14876d2e6ce3628d8fc81e61257007c18f5e6412fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150328349b277be4f706a93fa0d09247124f348c50b7c898a10f854f850400e59769a7e2fe9e9d1852f4b509f2ed3bab68c190e79a3df00db9a54ccea91d6173e1c0c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha248cd6319d4aa1c79911e557719cedca9cc864bf63ffabf6354250498eae6127133d27278ab3cf5443e21848971b7323c80d9adbf84f5cea89704e6907cdebe635d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f0cb114144595db08723e1975841fa068d5e2d80b9a8b2182d91416376b6a90ec7df34277eb9ad0aec6fc4926b8503160745669e0268101af62338ef76805f8429c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4604df9f6561f8607417b87263a49055b7dc993a263ebb3acfd88266f2ca7763eb305000dee94c6d53947be8d280374db9f259db26678fabbd382890df61771e99b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc5e4de080bc2318b236d19e0b4ecbb77ae0fae959bb0049a1764a7a42e83701b94c12ccce0ad5f8771f9267225fd3d5c9e5706e7db82ebc94b63ea738176484e412;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a995142fc7d92bd9a817036a1d37783c8e2607227d8f331c2265ba1faf67326c442f709293c787b3e02042d6b5b085e6ecc28ea13c4921e71ba9f71ba0b2ffb8e0c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb98ed86f6059bc09f48d014b36bfb4b77241ed980783202e8dca5d04ae0f96d8fbb1e3e1697bc5dc3e0cf3f7e21f35a82a9ce63cf9c0a37b05aa953c2dede2d77726;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71ef95019051b0fcb9a940d2179d55b3686318ca09633878bf6ca4a9cb692ed6bdc06d58961b336cbece80d58cdb7b5b1dc620a7ef6b9a35021c3fa9b00ac1144a8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hecc24c0cc842eed51fd182043bf869bd7cab2168cf078ae3ce7f81cc143354db9f8e348cbbc16cfe97549abaf44b7ada9c78bebd047e4d7c0701411b59cbd18a58e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1e9789ff5a7c0458aad2d3e4747e35ef059d6e88c5af242d58694af2312c532a23c7fd34107e2d2fa0bf9f7a4acc0b94f8c4c13823ee29ca81505b62bafd792667e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefc8ec802387f2f23a64d4394b2016a44b6f1b55cce0eeac14a2efa7131a1f6bb5e4905935a945a9033a3b7ca38f6cb83a207396d080276cfeddb425204bf6917a56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4214da3a045707bd99315ba55cc32c7c7d076c8d33adcf42052b49fd58a01c2cefaa4c9cac1a873ac057fc97965a6bf582c013690c15b004558e0ae50083bfc5c59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30ba9db81fbebcc51cac43d16b03f4f36bae97783592c47f82bad3d9c8dc9d4f7667272a6db88181341e6eaacc94faf234a1fcdc6ea129ea682e6c8f7056f523f27f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf79b4aa16724eca7d14418fd122146449474b28e36535c2dc8ea9c1503cea31976b4f3c1188b889865555755a372f324637ac041a2c7e23795ff5b9a0b0d8bd72d94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7a419d81aa08e0928ef2616e180fe11fb90da4eec02cfb3f2a85600c94bc6d88328ab42580edd780805684aa59dfc8685bda954c6f2a6d1937a22c011df1411bdba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ba0e5e1510f1618e6190bae9c71b34cccc6b5cdbe6f716b54089830a23919dc411f11160d30f64a06b73cd15919dfdba41eae2f96794de5fe305c09d9f33fb05fc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79a67aa2c9fbf453c93bc107c8aea0d58bf0aab4916737974f68d9d9933dbdf74e0e32fb4bc6c72550ae0332784fc6b356eeb185434d37aef6d6e61f3127311b50f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h640e89cf11768608cf307931fdf233dfd0e05286c0ea876c5c1add8dae723eba5c72a4b190f0a5278933826f40bdc70f70d5df516348122a88fcf0afa174648ff560;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d9913c66be105663bcbc9b1712e9a65a7adeaf71b0ddb6d498191dcd2bfca44e6b8c6b4499bac3861f0dd1a63c09dc0f22ee8a2607464901162834537b9ba92ea71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1251bd6f5ab683cd2ea085bfd987516ca068166e4053327bbe3299736326bb8c7dc2a2b97bda7464929886ec127ddcfba756e4903ea45e81079c897142d351f60b489;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af0f2c0d766e8c1b350a66b70e24b15a52c74f7166cb350b4b677d7b98d200a65ee7f58869b2ff84ffb72dc8a9b9b81efe5343738937177b50e61814b326246f090b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c0cdbe2cdf61c48f24ca7f5fdc0cc5a567b84eb715c9748aa724d7a436e5eedf89db6bd5745cf786ac03cd2c618e0a07666fb6fb40e3056bae7b31a3fd350230fd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ce300a821a33b5f3d948fe3d72ecc41786b1c4b8f95781d301d52c4dbd06143d94be258ed0b9713d47c58fadecbeda49e40f2aa43c29016eb9ff4e90669ad4b0572;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173729733a2848106fcf796bcdde1484232c232c3282397ece2ff558598020a1e91b70e5a6848090da9bff0fca03a82dda4bc52e552825516709fa692e3e5fb81b906;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9783dd829fd10f9212e24ad5afbaf3f7f00b8d62cb9cc6c63784d621c49542237434a5586d5e1977e7d64736b8ae1b79f0e488956fde4b2e76a7bfe62d8f891db3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1467342fbd36d905ee918b4b127e37c52a65a68c1a9692332d3305c221fa37c71d5eff2b8e801c9588e1a3237e7755aa73abfa88e40045454ee859d7b5299fb39894d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4118cf8407a2a35c5da5ed86c06985fff483b188c7136a9d268daa893547d3702e262862a62524fe59ed1f532e877febd78dcf116a3db7c03862c6f8e659b270a60d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba95ab4d166d9346feb197b2ba86e168d4ddaa5d6b55ad5ac4a5eeb9e784b7de64a7bfb7d71d0b31c764f33e901ed5144d1241a965af1eeb72f143cc934109efdeae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11891286d8421ac45dfe2bddcbc2fd25b12374d6763c726ae3fc0111580d5545c8495e9be36672f7622daf4b3343e03926f29bb6de0b9522f9888cc4d70ca6c5ec034;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140a2a339d54a1ff1802dcc369235f1aca75892d3ae749d3742cd4ac63f0b6e3d511e5fcc436f2b935245d05c71879267d460c5f416968b3db0637a41b7445ec0e37d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2ec4fe8c45a10a786102e28ef5ec830778c22fd93926d4cfa1cfa1869862aa8b33ebf616bbe8580ed6ed5a3656a072c91b07437aadfcc6c1ecd075904650e3bbe37;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a99c19dd52413dd04ecc0e5bba9e837419f8286d474697cacd707e2dd476087ce1864625a4ec0905cb3a315c253e150b9621635bc4926e77e3185aec7c4e15aedc95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8d26685e90b94e453c5808b6c0821cda8ee78a8f501b83bf2a0b13296b1e291f45817ab13f37808bf627acc2dfe911e559dd5cc8c86584997731f77c8a714cc4952;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15eb8fc128c6ec65886a3a13e09c26f92b6611304fa20ba567e76465236ed181c3381b7f29200b3c3d644c66d6e3654d8a4927f15f2951a059ec2e2f5f9832f4c5fc6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb844ff2ba49818a337a0708f28f0d4ed0fd5abd15458fc062fcd2f3452dbf183393906f13c79ce5226175deecf9908da48bbcc9175179af4acf5e77d18888ff0339;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198b1556efe7d8f95325c83ead46e2aeee73587b2ec590f262fb3b0ba05abd8d7f1eda07516b7d9b08cc5e2610c9ee1255f0d6e4ce46ae1e057e73a73769b73e1ea46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14601950b74133df2a29e4343426eca3d16f1ddbe7f4e4dc93b4298964c0b92ac104085c1bfaebcd1324e6976df473417ffe8d6a51455c2e6197a61bdbe3952d74227;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18193780b6e5dd5d2ce6c307d92e9df3c2c1b73f5c1a34c9bf66acb440e119c092c07d4af39b7c8d5c309f9438ef7669e551a8512ea9c09483e915ee819f9356f26b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c282a1f2a975118a60b4d8d7f7fc123cf0f92e2776639a994092974ae188bcbeee791fd9f364c8bbd744f083fe1fe419f62ecf1263fc8a9dd265c6561eb04da100d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13af49ee805eae4c5883039d08dfd507cf8847dbf7ced324cd80980262667673c0b9dcedf6bce281fbea0a224eb2b2179ee14d4520037faa707b07a1bd027df9f3447;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hace43af80157c7ef927ec9a6cecabfbb746e6d029b2583533b27654588052d043df4c83e06136d7b6300e4980a9ed01583a056b203b1edb433b9b6064dc6f5ce33db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83cf954929e9b263a4f884d9253fc300d2800cf2a3f3f227600e85928a92f5b8312911694a6ed0d3ab36cf59257d00ec6340a9ca1352325499486b6c5fa905acc986;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfd06226d2e22de71c8bfb8a67b1dc3f3425c8090a60c140784658e1d7bd53619623af3129309f8c98ffb1a3fe4fde350c3ef2dc552796d967bc54f3f5d2fd4bbb52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f88dbae3ab0ba3f4aeebee0ca6104b6c33812651539ea228690f11af19901520d6edf06a5d12d57b283a90172b0d814731ee9723c52000e74abeb6da45cd8651852e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e30ca16a5f5fa790fa5507074c631486cca13d6f111a59917396d0ccb10ca90fee9d34b6d482a0b4909f186e93b1dad4212084254652940ef3f0b693f31d472c187f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154800494895eac76477eaea6078e35c06b2dbd9934a969ee1b9a87c5f3a3b6d24423739e99e195d769fa90db099a2e984fbf0769c2cd7af99e14e11304c3a7d423bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e9f38c068a3d21da2eb3da4d4845b7b1cec15ff4d04f7dc9a39b025f02b98f59bf056bea785669c7d2bfdb2479ba50ebd56e0820a4956c2541dfa77deeb726e9cfc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eb1e2e066b9443e5c972fa3f25511eb3995e51f58df63e3d8368cbfca9a27d1b25081e0a8f24bb48bbb215708f21e736610b43d9ff564817e1d626d5a17b4245262;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d70c87dea239cd8bdb2d8755779116817f0cd74e0170ca0663213ae8d9f28da1bbf21a95dc5655e514bbcebd362eb43a0a8c69d2a1c8b3a8584b9a5504add4f5ca6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1526c1e0a3b01ca3af6134b251c316cc46117f35031737f1a351318cae6eed384ab48aa60aa2e659f3cfb48a727b795af90a2cbdc4357f7f925c71355541e56a1403;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad1c5d43338c49d53820f70803cfdf3fb80af14aa9a81ee16ffe12ee1f599c4305b2be23836c7f8c198c1633a9d24e7e63884ff980e6ca07c9a283a1ebbef79d8e99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83dcaac792aba4e36bd7bf1660ed19dd4ac19aa24f200507d58ab57e1ce624b27094d3f946ab48c105dec9f24f7b905bad0ae5623ebb84e534d45ebe1f0855b5bc6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3bb68067ffa852e5b2c0871c5aa0c198d994b0c1d0d43f32450b3ecf52efd4396073861caf39289ab2ec809c9419678c2853c8bf4b9fb1905ee63c764782813da02;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7dea084fb932fe9baa29dc00d83f6e048a5e14c3103e58a243153a43a5f083c80a43aa5fb5b484425e2cdf15fa4352cdaaa0bb4f30b565d8142ca12f957876f39cf3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fae349daf826f6dd78c98c0bb917b1f5051b4cf441afd24b17f765d5839f2ffd8dc5912da41fec6f183d5a007d5f30ce9b6b1af5e44f75bda03d4125029ab05a65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165d4ea7b380adeda7fe1c8820eb9f9a51f4150ca682ed870b729603aeae636f9d39f1f022b29dc074f5184a9adcbe63d97f99fa1f547450aa579662278ae08fd15a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b2dede6d8e8426e7b5332a2086d05b800e03e435c074b0c46ddee87f12ec748ec6e7321007dab3267a7fbcabf138cbfa45590daf54a1a1fdc4860d734be858ad44f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3b5bfe1e88e0b737f31a7b3124a768613bf4063c16e32a32c092755c82169bd14a31e7de0af30c43607c0dbaef436edfbb179b362ebad981bab29aa1727d97b0488;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27289c25205c764b167bc734bb540ec92e052d1a4ad8c62fad2f042b262db25aebd934d2607ecddefdcd271e66d221e9c5863b4cbe80a8e22c371f208edec072f050;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f6d5791c1cf2ae46dd7208acb48c03cf15467b5ccd76f179b8201c949e0739c91afa6d55faf3e9b694dee496ec44649a550f03e0e8b41dec1dba683b8313f6ea9ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cdc336dbe330bf741c14b1bac260eef5895091568aa97b63045907414b088dc6addda6b3ce461678d91b8c06c9566ffb2ce151efc6fad362897dd8886e9f4e4fea4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3116bbce2e32da1cc1395119d07fcd88a61732eed3d48fbb29f45eba3ad727a459a3f4a7de9506fa1c771e6a4d84dcaebf86e26df4f43ee06167ee9a530b85e08dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h660b559c3cb97edd820a2fcadaac54ee53834e55bdf90e74d19d1b7853b598ea331c5d9e55da9e728944d70410dc9464a6b1ed50e8e5630501893e835a84ca7a17be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef81ce5202e2da19d87d8a4f581a4e3a688d5e58fd2e4ed638f7679d918ab0d6bd96c3439fa7a6343ad757c8ea062472eb15813eb1971497866fc9b6d9d3a5caa7e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160800e36d080798b8e7d2d5fab26a7b035d61f03219629ee32fa439a7896fa3247f515e159b1855b04ff99e3c6dcbec3b9c42a0bfab6405538de31cdb2389c050556;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd691ebf4c0c14296a3f95162b78bfe6c1d56e007650f292c358897d3cdc256a3953a71115796188f40963a88baed413e2eaed60530e83d63431dc8b131525b30c5a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a92bedf7098ec3a2041567bf3488acf2830698aca051de52122376f9869887062bd178685ad420e47fba56264213a591d362de0425fa24f9082e330c609998d84778;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc1e948a960733ba6fc018f493a9674f9c7971febfe373cffd724fbfd31e4afcce18907583ab93acb8d796a4c9d14286fc8f8d0a1f3812c36d0b12ad07a9cd89d0ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5629bbd42ba4743a697c04a1bd8d70dd9be550e5eba498a3dc2e004c74cc6b6776b28d1c482525f96fb56dbd5f3c259754caf4b35a6f55c814e0f05a66337e2e01c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h944e435781fee93349b4c9ea0c758ad3e3097e08c6b38ffb1ceaf13332785ef89125cfe3821e15e6c9aadb7e77fe69f337ac7ed2fd21154762dc7f66e715f1d4a0fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b1e493117a2d9513e702b3c340b02817219a6699c602cabfc0fea10fe80eef80b5da71e3ad95da5804285320d3fb1527171146c645bb49c6db7a8eff925137e399b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106d0e76c11d416bf8aa0ad933ec3994c0dcacac6e3832710ed38c5e3bfec2c5b9c43682d7814a489656bc4db8c15d911de9cc213d8c3fc38596586e346e39c8c9027;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1036f636891d000bb8e9109edfe144d51161f7795c1b5846b865c381c8e9aeec4dd2c7681f766ddadfc61ed4ecf7bcd79b977808a8876ed91cbd28692d857561d1fe2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb439b42909616eecdfa084169dfbcfdaced51a90025da7586adc4f09b4d2849bda24b40d1a561894fc0ee454fc4a5daf8f4f37b4a7721d51b70081eacd832482eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1483b0051df1704753d2d419b14441e64e2b670ae1f1ee4211fc1d4934ccb1f856590a619137296eb3384df57b61736871694a83d62bc7224e72bacb349a567c6bebd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h997cfeb3653588316fd2d72d47571090bd3ad3474f42d9073bf11393878a32ef0336fbf8d173c2e398d5cdfdadef0c879dde7ab8e9bdba3da90244fb4fe975fcc382;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd642cffe0ddb420a194b7576f595c78e7506a4e985fe43377edb0e6f4e0213494b19e959de207e9fc118a4a8665bdbba5f6d8e8bbb6d0fda08201a5d6ed0554658f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h634c5caa37d21345e8800806bac1ada8985ff136d18773c2619a0d2a011ef94dc9737e96f44bbeee073c04c96478480f38dd3c3d4ab32d95615720fdd9bebbbe8f07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1175b7b2c3ff9d96943d2e88a726cc6cb8ae4ba23b2d247872db11d760d6fc59e964102c527fc956dcfd99148d20240a619128394cee7a607a1e81446ae7df825f7a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120621587c542a689d21eed8d7bbb32e194b353c40dbda875a25b7a73539fa49d6009fb5201d0a3ed7fc14f93ca230b33535279a8e580beb3568011b5f6f298a3cbb9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1922729936452d955bdad3ac4183ef409e74022115028407a8a9e5f129c33fa161387cc915e92fa1eeff98c439c2a92e8ebe706e4a1acdb573115a7f7644105784ef8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5322d656a70bfc8a05d21ef8680e95201d219ee430fdc5ca153f28f7dd7b06bf1d90fac6d145a8bd8473c36ccc24efc2f189f5e00ff37f5c5a4c64b98c0e487bca82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166ffe00d54c33d8c05a3de18687c6d58a26016574dcd7de33b4664ba38f68ee2f5fd342f4494ad38fb28e8da7c3f0924a45748df83244d53c17c290160dda878f90a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7facddcf6ab603366475a79ae9a9c898e587d25fbb687eb252cf7411d6e58f440de813a8b12a1913a9aa9b2ba2fd739a15d41c170fabe5212e6712b63f0c5fe51068;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69906842b47bbbf639620a6daece9e9d069ae732f1997a20deba8320ba76748e9e2a86fa3919504181b012097c15cdbf2e215245d40d7b7d625c7d8bccbc5a40da4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha18958c6f44b207de44856e85e1095cf8949c8cb6f3f863bd226504600d3e8ad2fea055feed6d6284ab4781ce9bc89347865cc1cf156be2c33a20a1e450c7d8863c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a9fb4653a6a28a7558344ab1cf039c06c9869c6c2ed06f1597ad94d3976273e0ecb4d7b1552cb3dbf86bf08bf285a052543aafa356a20c466ce0dcb417c886e2e1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b120b8c4758a9bbcada1c2bc039e5ccfa000c48c1d9bbdd09fb55cb72132bf0b3851866e5ca2f23887419b3608153f88edc7e80dee602a7d1d3b4adb7368ff87de6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed6fab55572a3cfea2dd844ef63a8e7e89df285bae52aa5e150405fb887d6a370f02b2c9486fc7464de3d607ffe99bb4e6797d5e890ca2ea0f33111a30ee8ba09000;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a3d8f4fbcfc488c9842511e9791e6b648aef717230a60d70ed4e996b3d66daff09040315c716e2c91a61c3a9d311c9273ddd359acca5732aa3b44c4e99aa7952248;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cc2a6992da4d2a7dd67c11d6bc7a6b51e716cba80642d7b338c2e487617e558375c7838f2b8d903f7e74302b3788ac713fc5aae84194d8d461efd0b0be7e2c9f91f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b4093b87d60419312dbe53416d0770b1083236d725a72a7ea2b49c16fea1ef838f862ecb97faa79b2ec015c30ca89dafe556e4d1d5ee61a39a2e2231ea7865e3706;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f6b473df3e4948debaecf4797d0eb5462dfca8902fb4c2a3e7efa5aae487abe2eeacba10fa42c7e72c11e32651d6098b884dc63876992a641ada72e9e588d92c9c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbff5e6e3cb01d729fa9928463c8e014b8a4135385ec93afd3691167722575e2073b66771719daef7fd494e0e09d094aaee8893bdcf48bd48e494bff2b09ad5546b57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ff0d0e20943d73024e043e372bd0a045ed3b3027647dba2ba8068ca422135fab321ed6ed260d684fc7f28a8263b393841403e60d5de5e7aa530f0b6a12db39d02e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cbbda5c28eaf726e4b6a6b1848c49ba22510d04a89fe7e9599a6164c840ca66bcc63671c7e47318b8ce37ca5af85d5829ef846b845608455477b583f7f052ddbac7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125796f7552b29ad5f6d9e70a83a363f3a3a3f560edb2002668eadc288f6f1d49adc990b73ee745dc168334ac15ac1de70559488a919413a8162114868a5d787daac8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b6c68559f500a23bfe7f37d301ce7b531d9b2a5f91f6ce82e1872d836bc578918250a321e934cf8af5d8064380ea49d13c3dcf9df0f5918fafbeebaf788885fae24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e576a78f8a910d1f7942ae58ad6ce195f0062aae16c38fea517d7eb94ff4c6561ec0be3fb760960ef254d4ce929485d6ab001c180f4a18aaad455c4ea5a39841b22c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64265d1f3c0e9d8fc8201556d8f937dd3d2e86ac2bdf300fd15481201cf0c2a1b4f7984e294e6f1dae07ddd859cce713d0d1b68be42a103aaf15bd423ae5b77837cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f7e320c60a84e4f223346a174725bc95697c2e12421363a509c6893581369557be988e186351bc8d15d1cb64a9e0b1371bb890a0a71dff7fc4aa4caeac82b83c401;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8208756c3d67a38f86dd886ec8dc137568826def7316ba23ac56ca688335217c51819bff3308340f48563f86c935e0378b4978777a9ed3348c46fc64cbc289345c22;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b74a28991fd81026c907b8ae58e2fc8dd27bc6605e58e570339fb1098c770057dc02f9adfe1ad2dc90d7aa8a9c8fade26d635095a265292e4bd86ac9d3e3c6564a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d65bae5e22d9c822510feeadb64cb813047d152f78bcdca422d61fee2a49650e3777ce46f0e3992f773e1a77deb147676991f936f318cfb0f815913a1806d898887b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcaacc6c391d307d7ae1b8de2196dc153cb2fa9fc5539293cc7fc9a50f93b8634e98284874eb3e8f706c1d3f236ed4bacb870623c1d8672bd346e12451c8dceec1a7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13765ca80da8ae87adc6f544a80ea94d9b0b03c9559e279b8993b70e8d7efddd7353bd29456489c5641af77c09357ebf1608fa038c6a697dd5f8fb039ac6bed53cc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c14782f628e8012818a17bc2dad28d8d31288fac3ea85a828d9330f883db2e3e17d24774baac2dd98f0c47d353c6a360e8b8407e71e9fed48900e812a0eab4bcaea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf855da2dfb81dfaeb5691361ab2919605156268fbcc5003a915aee34b5a11c5e99185f24f604138281c70266bb5f31f6c3ee735d101dbaa5780822c234c27a48ba97;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha866f3572b01e70fa8b6a197c9b7b114cc0ed697b32d0bb9fecbc06028c91210b69abb7a62022282ac5631ae9ed0e40611b7699411248bd79d8f67f4ee18eb3d8900;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d52c30fef8012245606ce45898dca96687423e64e24178f6dc0d9f8f8abca7af218af72c1df1a0c23c666b477da1d69d8a1dc90755c202e2985addf49bc51d3b9202;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101e44b5824d6145e1b3b6fd8493c0087057a54f716626275b64856bb2cd7b655d59f40caf6b761e76eb88361821b68143df6a9ea4fb4d1372b3f160599be317c1da5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7b191bcff277bc9e2d4d840bbb4383f6804763c6f504e782f7df008b63dc85cd81423b2bb89d7318c5e1ece07425d48f504ce9a0e7e7c702f775906b2f315131d21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he89be814fe51e712a7602a12cb413903cc27e0959cd6b2f0e77133fdb2b4e3cc8e7a7ef7c2d72e9c38f226bd154dd7c0037f7250550cedece1a7d0fe7680923fe26e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ce6e398d5b9261036a3c70dff1fe909e9207f2b37b1e34fe58b33308b44ba25832f52e9c166d31c26a751b63fd3c58a458c263d150a0e4389f2cb4043721f7fd33b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6c6b95c476a5b071436b28adeb80bc069769ad33884fc6da1b9f031a935c2c5738560aa52d5a6ca7fa32dd7a532765ccdc2aa2408e45996cae017639369afdaa4a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167e78bf3d9ba4d353436be688b6ffd1a5da0e2ce41bbba0fd8dae733de4dd659ab3820160d7cc70a3c15305c67fa074c338adefc0de387492839731c780d0aa8efb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1689977cc05d2cd5aabcdc2b0aa30532c0ba42e2a9d6c6e18f4f6e7f3279cbdb174cc98d5e3bf2604971b26da3886e1286bb36d5ee43a51304796202c45eafdc81632;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h995877ada190b9c930b4ab831defde6edbc340e2309173630a13f9df09a800a101a1fa69a9163da76d6d0efc6b07eeb3a705aa336679930a7ab6d2d219ebd692a243;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156e13e78bc9b2518e573dcc3ff04fbb4ce5babfed0ca8e3f483a1a05c8696a8381b19e1a78aac577162a9d0805a26653f50ed58030067bc54f832f508164827ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b7d355768755e5a168e9476da3d3c9cb611468da982776db4db101567b6b4be455c20abecb54121404f00dfcdb8cfdbf2983f64b36dfb8b2e0f3f1cded5ef4454ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7789252b00913dc6e50b832ff78fbcaf92da45c480902c1dc7d428f43fdbc7b425f92931cb8e2e8a6ee1238150c4372ec233f97945002d3a880997269d77192c7bee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180701b9a68816596de99e8ca28be68516d55eca71319529ab2d735ebe3bdc2c42a8814c91f9bece988e9bb7094b598b0df07b40d2fdc4060044a6b9c7e2b0179e519;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a15cbce2ab374d966888ff8edd070f6348b44d1b97788e9576fb2339cf4765bb428a52d4509bcc87e5117faa967b35f48c4d281ef58e6ba520265c58cec68545bcc9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c452684c38cbdb0f1cdcbdf87d1e73f30c3810e2edae8b6e24e1d0fcdec82179295e2f6b99d2b4b24e42d340beac2828ed87386e114c562898d0cd8f10140d2edeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13002521af3f11d2fd8b53140b9a61904df4841ca98dee84b2b5c9780cc735dcc82940e9698cd37d3cbf710fa602d7e24b4b9962ce97951aa02c9440f7e2c2a3f8cbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff23a47d639f43d5bc538d935b30d1ec23df44ee95c039d34188cce0a097f79dc59e36df580a25f420ec627200a039089432e3291fc5860f9b6454317f734bdedce1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146e295f610a174f67dd8076e8789ee4a641eccc8097dbb62595e39e50d056a28a84266252b3bd9bece3b5cb622c3afd7db0eecbcbbe0b3ce6279500a6442fb33c3fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101dca98ca770cceaa71233ed571a5d9eb81fe8a48f255df8ffca8f0d632a6a723224dbc41fb4c3e58ea8bd450b613c60b1b29c25ad08aa07e6a8b274fdf534722998;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86c59b7ed5678054ff8b2158913f5b4330be0f4b10b56a0386ea2bafe688a38a25bcb8abf9d2ce87ca1faa8235482096963ca37ee44f70967fa3c60cbd190109efbb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h197d7cd4e672b09d62485c853ce416e348c9934f28b14f4b8bfcf4e07b5fd9f08fd7fd1dbcc26c91a21334fb786b9d1b93c69f27302c15f875e42a75c87901cd277c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8a53f475c953a0f5d2f01fd3d08bb3749c3338876e43db243f11fad527ade2a70cb7be590d1b14f33f0b5bb628aab29a5ec39aa93bcbc515c4d8ac66116972ea7e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dff10c643de5087e889a441d254a4e4f992a758f991695b1603266823dc07c54d3a1bab896bf45226e6f314328e5880b7fd98f380abdd6013f258f7d6538e34ca14f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1132f0d56077aa96b593fb8494942d2bcc55fc94e4bdcd1b96ecc95e1d3b72911ed0b3760457dfc1c2f6f94f2dc1e76ea5512bec8f9ef449231f9fc44d0cbb90e1328;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8486cfd874b30dc09079725bb32b6bd24d8dfac41f28ff85c61a6c15989e6b5522bcb9e81a55448c39e482cb19aa6a227df3ed0638ab8f95cf0835c7a246f2fb6a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1233132ebf38441bb7343122e34002fae4473f902339bbfd7bad3edbe32b9072c88530615b3da75af7584cc11805fbd15526ba94b6376195fc6cb41bb72e79bacd8d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6f929103919ee458c69ffc87c963df239ae36469adb3f3474ab8abff2997d115f573e2fe7f7fd67fb63cf939c32babe08a8e5e95c15cc51c4651ba1a69a6c1bf949;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bf3ba16930545e323ea132019b25d5675ff938d136cd613a34c39d71ff1ffb9e788c1dda9a01064b0bb7aa5267259fd076904750d7396adaa023abe34c915b82d3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96e0839d4bac104b2fd87110ba051b7510af6e835c3773ad6cac84a2496e7bef67947e28a1ddab97aa7496f428a0d4c0539cfe894e049532d31efd60fc361eea1a7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a46215d4b5d6c035c168c86541d32eda81872a43e64d04366df250e6d037f223beff557daebd5d8876230e4dbc5c4bb8d88f769ddf7cfdfbcc6b901ac9cce50963f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11846c725b468e2e03cd85ff05dfb603041e2385a4be2a67176828b3f8283da42cb3115f8024e0ac37e576a610baf814aa2a0b906665963aae9df8db90e5a578b7157;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19480fdea919944cb417b74d94e0de92ce436cb26d29c349ac71c29da2c6b16f127a5b122942177ce65ba9a66d5e1b42d56345b3ca3c865d4dadd3717544b8bde8fd0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf5dcdbb2c1e9b8987917c0ee0198c540160c57d18aec2bc899f4010d0b618537d0e6d52b2a7770f98bb7b899ce37738162099ea89fdbc690ed6a84f63e36231b3fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe15a7143522384114fa0412eae966a303c55d287784fb01bf6a891f7560e5ffbef5d12121b9d6dd582a04bd5a862f0efa94c801d2907b445afc0ba10e8c67a10b9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6b692eab14f9be3d990aa86a28cea3b06d35fbd4dbf4d40812ba502fe1c71f501ab404b0d0f6a183e12ab57f2889a6319abb04c7eab00f88520e98ccc4ca9477eda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e43c7c1b7994fc035837d7dc4041121d803b9ccdabbef70243c578ed94966710b75e1a16c5808fb61fe75e8a2e04da3bbe8d461ef29ff7fb982e7cefa78f5984fdeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11dea93f7048b4a616f38f21dfba8881e6967271cacbddb8365afefd62f6b17e3d5eccddd3792cb8434ec522f325da667ab432a4e6f067d7b98e2c7528eef10619b8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12165a4d095092b08fb42eb0d7a9eef3e193eccf73bc60e3f6d73f002e007e07eed2c1eec205bacf8611bcd40173ba5ae2eba7a0d238b8172385364614a693040921d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ee5ff6deb06332ec0b51c5081604670e547eb1e5d7ad1bb87282e07ab5aea2e2625a71e91f44f21e1112825fc7f3c659f8a62d8b80c2a4afeae8ec453490bd95802;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68e90e1b295b01d7a0d7786b713c257311664acdc991341c4502e47ec5883d3808758d28c3a8f0352d97ee396042e229fd2f9a095ade5c493ca94185ce9a116ee844;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117882fd5155cddeacf386a9776494db5d35ce88ad2703f703d53ca4871ceb0eb458e84acb6c08d67ca0318b295331a9f4f65da1b687a0982b6b4e655d1816c10f0cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ce25fadc1576be359df18b5857033fdcda367c6c322b838421dc6acfcd03a7d5f2d859f1b3146ebf1c8312aa7a1c25e9f725c9d1792367b163c3faba9887dfab916;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f4f316ef463d13741e286f765fb0e4048fe43793404f6c5070338caaa5c5dd349f566018dca30a6870bced37debffa61e28b4529e12bdfae0ab474870f04e858363;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a8adcab403f8bd4900037a142be378fd2ae0c3ec905dd0deaabb93b2a6f6d96c72fcc6312a33d621a164239df48a756dd7f9ce0338d4a88ebdd2e704012892f9d81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13acf54a853e88b50dea7910eb60f189840326588ee3a7a9af1a3453042fd828afffc1d7ac6545a086c3c883f474f2e7451e4960dcc7fa92c39278c39614f5831f930;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1802b0c6f18062e8dc7ef492475533989d34131424232e00d7f0ed00435083d4e0c66f07c56b572e454c999663d1943bbef2e4ab45c8a4accf78f66dd62b0b4376663;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h940d0f3b4817876e7f27391c408a607cc01201d10ea285a53d767d8a7f5ea78720fc7f1470a59c53d508289f3bb048ab9cb69469c13a88bc1f5e40ccd44f34b63a34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52828034d913aec9809e325104145e699add3d78c15b1dafe65602de76d4adbad4974567c652e6e4eb8b42846ef889a5a87f82f693703c1e9c648f968852218916b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebce939eb2a962f4a290d48c025b6d2a1ab59893404662e77ddfd71f4547559857e32a0387f07aa3aeba6065231f481d14c9c32af3abcd845e95fc33045ae122893b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h480c59658844313fa50b8117a44b9ec4a4d36ed8d71852338a26cd9b72bb202475ea80e6c270518fa899b8563df8c9b60375b2f5dcf970426046d76928b5fa8b0cff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefe702df2f7165b4d030a07708f10e1e748826d731875455d9b9ad328d0142c99bbad311b3d87180a1228a38f46ac774a36c0dacdeaed0ac0d658e7f705f04b850a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd2ec669baaa01f72454891f0afb937c807ee2b1f218a8fbfc6d7c9c4f2d31b07d267329543c2d325f794a23241d23478bc21583608371f1773dcff77dd0f0ab55ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfff98ef1fa97add529410fd7620942a812a11a347cfee83519d4ba09a4f443cffad8668419aa9d5d8502427eb4b25d073b21dae00a5367fe08e7f7e6e4bde415f4bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be6952108063abaca110468f51c07d44ad7ad376d709b1b7c9d30f0e251021f792b8d6349ca7073c9db8d9b861f14a1b469ae6dd575be0db7a4bfd9d227af72f4d6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1267ce8d72774285f931c595622ecaa090a8ff4328613a2ccde0e984b575f619a27aee676876659b89d62b3174ee205c96360b92c9777c1bbd6a656937728b11cda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14571687242019e1426bb22e148a6c4c989b45a02405e3efbbe51043d575c3751bc0b447d4c579eb018c90ba3a8732b450dfcbfb101ac89f704ada3d52ca36c07f798;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d88383703d2674decbcd7536bd520839396f1ff6c1db48b7b555290e3062c539cac62e5c00a8c43c97a0d394a6e1151126a30f861d7e3f39b25c1b5c3d6c8541397;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186ddd913cbaade297d5110b3286952f5cf2fb91fda51e004253878be2eabbacabd225a11a6ba30dce54ebce55124cad21830c95c8081e728a332f255d622902e253d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1894bae78ecfddeaaa4fa2e23e49000b4f9f535ed1e136445f2f03610c5c5ca3b3e82f7c557cd2847d71a54cb1b4b4ba3d90af1e52430e3859d44fc3f60e6c52272cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae630c55a02ba1569c3c4d6fbcee3d19147b178e21f41b48b6da37dc130720b1b94649a0699fde5c3b07c7d86346ea7ba79b26e5cf81a641a6f1db51a113f98422de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4810517d8991bc04cb8faf2f9fc69b05e7a279738050fe32e6dd76c16a60ed7e14712ccce829e3276c516d6ea2ad56c85237e3cd5802b164724aa54ce5e50635148;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6e568080bdc2b681ed3b1bc5e03fdc65d1f295bd2d470f7b72fe47ce8a9a5721f6d73e52b3db66afe5a94997587cda8bbcc00c2c1a33de823de4adb521b5bbf5d4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf7252b5c91a6efee5006cd385ca651a1cb7c32f9325c6b707559893cb4ef8c86c64b48918209e107b8f017e3179ba03bb6abaf3640cf3ca7fece0af42f3efcd1a72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155e366e356511e8deec9458ff823f793afa3c00083d93e9337e5d6ae85ceca75005d5c7f4b9ed1e74d306865b21b65c1e088fa76a66464a6f204f6ce0930ae6e0690;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae892c75cf3db42afbb572927ae69f1f91cd66655c7ef1017360253de61dd9cc15756d3db698b3ed6afba07177fc8dc71dc8b87f684d7e814bc39d33f8cbe47ec9a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf273c381682ea8863185671b1dfa80c639a879d96eedc09f6ce5e3b8d52fa6e8831dabaa3665a163a3d87b755a7ed3bbfcf47365adc957b0a6ad1b4158d888900e4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50270a3adf0d975ef434fca5b12d2dd41b2c64f659a07fde4916083e98909dc2400174a8e0b52c6c5a5795675499458a5fdb86c83d66706f90646dfb1cd8e9de5cc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16135fcbb05083227b12d40f8a434523c6788d80ba4397b2bda75385284405f1acebd04739193f3bed6e3d1a8719803aee3476c081cacb57a0fe6566f43f3fb399a26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137af23d7e5584a5c31a011a942cd2f5703d147d0c56f846f4b32860ca9504f47baa23d5d3822550b62ed5f301d24cf48fc883af0cc1dc7edba94c083fa0266b094dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccbfe1b534bdd8885ac8679833ced8ca8088f69edf1e4b784e9dc4d6950ca6d4e8220e1011286e02be21d40b70481c3df0132b3ef4b17cc4f8ca40de741ac403dca9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d7743ece1e55c97dd0c08bd8bf45a9f44c99e873a1a19360187d17d50d0af38a2444e41fb199fa5977039f890f45e6877391b44a019d083c6686dc5a2be7b8dd337;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b89975b585fc99cc186859afb4b90be954eef22f62bcad47a4bca0cffa88a2bca2196460e41a74c80df7caecaee5880b1276b171e95f64f33537322e6c5aa12def92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1330619f0103719762e28f11b8f37794e6ccbdfeb304f4c1e34a4ace8c5691cb7bad24793a33be2fa3362eac0e3c7304011d876e84576067b4b2e878c1145f25a9b05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f925009ff23634e24c867e42d61865bf5115c4ec617b443dba8223e1dde434ab3de2972ade004a2af6890acb6f1c3edceb5f4a31c650ba6de3c811122f799451f615;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc123fca2657b0859d66dc76149e26519b072c729837669e390d7e2842c111cc46ad5e2c60175a93e5581282cb3bf61990e557bfb458582431c7d12f58639631b1225;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ded03d792d8a5c532bb505380f7c5a11c60f1a89cfaeac3760e1f4b9fb059006dab63e698881b9fb0ea5708497dd0c94800e98b397794413713dec9bb349c3cd238d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a2f930a68254dba4d24501d10941579f382955c45441f68b151f59ac151e1457e3de7a4cb9a049ebc86c5bcd6a78cb3b5628022420ea9a3c3abf892d6b686be533a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a580fbc6c094ba5e2314bf23c80cc73be58bb6d7ea9bbc93b1c50693b8e748d3508d5fc0d099ea7c8c47cc9d4f8dc965dd3b329b3a9eca0719659ae46061f37c00d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a54079e2c9fecead7a0ff56adcbdc4b027ab3491047b71874e3cb9aa9d67a0c3b83790adbb542ae9aa96cc016d0de0e6056af1a16d3b2da62a97c06838c3ac64d03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e47a742ca4f27631987ba82c43479c3123deba86cde807da960270fd812441325b5dc9f48cb144bbfff224edc62b5de2b8e7d501e874c6de63b572f5949787cd207;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4710b14df57ce126eab333cf086bf20e2530ba37a8047ab0af865aebd39b1479501519498cf03eacf37892bcaefeea36e07e0b764a7006dc5ac918bacc75b0b98eb0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h572e824949a4f36938bb547b05374535a6023b7f5c25c064dc570100686541da30aa17d4d9679c3b4003272ecd7dc2ea85760bdf86a690024c479a7693679fd23407;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2daf948b055f23aa9d845f38b711615ffdf2a6e1dd78a730345f6a0ab43c38c64532e7b0e74cf2ad956edeca938bb5a13234ee26b1afadaa8faaaa64d40753db5e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d86cfecbea7f0544a340d054bc5b0c5d964cd77f5a4490fb803d263e32d80b642c189f5f69dc282f691de0598187552c4a6927968cfd256ee5ba165eb7c5fd5ce19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80cee3e2192e6d4fb2e0f29c2fe3316617f9d42f9640699757a02db4237bb182ef2e89e3dcbffd022f1ce4864dfe72dfc4b13e6b68a2ab015ae2ea37e47ef5b3af3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4d3fa601396367959f3c9ca644520921e19b212f57a6a98d4fa956c16397d4795fd4d5fefeea03daa0467a8d3610248350c2a32b1bf9da4d0d43e6230b946578f50;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a5bd2c1aaf0790dd1547bb57800f966820cb58956b90cc8bf4abe473b01bf4fc69d0a89f56b6fc265f4f468001eddccc25b2c314f4f3d0338d67a5b37579c695ef2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd189f2202f593f5cd926fe4759f7d389fa56516631b68195556e92929d9000651ec2447e046f59e9d8026f22a785377c84a7bd926f67a223e1115334c6614c45cbf1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b33c9fd3a8431a2e6fd30773d18efe199c4f31431c9502842ebaa1d2277790657e0fbff29bbec773ed1590a6b873d40be34fddd1d7f54a060c7346c92848aa2a49d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40ff0933b66fc842ae617553d08f5345b14473612e42936dc3b70b4eb1e1f638876c8f56cd7915c9f643b5c24eb6846041016715cab1c7e65f905e310149d5451192;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134ebb48d74a130e9cfc6efc21cca2d1535db8bbcbec1f1401a27fd0d8f76a89a06761dbd0d36362bffec02670d0d34b591cac20aaca26782da97242abcfabfdc8ec8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132d3e67124c888b02dc9c42c90bc4e0ed7f832ec7b501260de9c573bb2718aaaacebd97a41a750177144fec4aaccb5a2e9491f26d13fbefccefa1d3ce7655fb0bc55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e1460c744c62d46e5d89e2fe1a13999e1b8fa9fe2b1c241d0ebba4e951b3c333a99ad75ae33ca7bf91c64e697ab1a173a34a7c847e9e72e463f2a2d1357eeebfdee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5d8c2b67e854bfdbcccd61789604842171b5566232f7975d27ce1e9cab2582a8a1c464809d8588a3bab6d19352360ab40239114146e806cf17b8a4b985034062eb8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3176862cfbc88ad48beb46ee83170f4903d1844a641f359ac7b517066dbadd49847900dc8bc62b792ee2deb09db2fa3290e36332d1a0be1d0f1267618eaa55bd6c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f678762335cc8dee39731abcd6e9ce11123f3b9a2d999b73e13073a600f1404fdb142db6eda9ba728dae6f2d376f67b81895f90404c2c7578ef8e4300a75b311ffd8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c07d805730613d35fec2a51110b81ef721cbd82ef068bc77cf7ac0a8ad2ddcaf40676f47072a4ed7a0d4c0fb1615904fb5065c94f9cf3538087c63ad71d2b07e5ff6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1719838c08410df721c9c9704fe4941c3dd364d2d950184f38dd60286bcefdcd39878bd667295c8f25b5ca2e453ad1b974f8383edff522baf835492cf45a805e95b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129d82cc83ec2eeba6e9c2b1252dc75089a0a04bbb34af4b1062b146c0bf576be6f64eeb89a06bac39db42f59e2c2e4a2503bf619935f4cee8d4c6284325b13a680b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e16bde1b4ab34c1d708007f0fa59dccf368ddfdba9b60a51488c358fce8634a5b11f9712de04caa2745191857e0cbeafe5fcf7b2e7ce6bbb61dcbcef7be5a2285e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7ba2b31eec94aae5d724729e95ce7f43708dd485e7bcb14ff04315d23badf506ce1e091785ae1c4ece60c61700095c41b54eb6ae4748e9221f0882e8315c0bfab8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf0eb22895408e70bf86687a3b46375e3da9fd4de98e4d10a52b3280d131b4d64deaa0f808ed8e00d930df957cea7a7b122faea077f81e597530f0cb023cddf610d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde48948074be02ddeac4d696de5c1aa29d5dec103eabf391246f7940f05eae61265be4fae2455cbfed07144d21caddd63a00d6a1dbc1f1c696c7d1d4a8969eecb73;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165e06976c6760a9d9ea0dd92a8cc9fb511993f02a6a730fb980798f252dd0ea3f89d84c47683e0448d187fefef944aa248a06571f415cc238234c9dbf1bc03eedee3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9b14fb89e6962cdb5fc6687377504b68e3d04b1f16b58e655ee461044c418054f78da04d4e172988f86ffd9d554a6e2215b9afac092e058dd96c07ef7163b445104;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd24992098bcbbdeb935f02c48b585a56291f72101ea6a00c6edfb3485b439bd4678ac65626398c102f858eb02ec3d552dc1bc894086e11b081967373ebcbfd973d9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h487a40b89bc7dd1af301a11d56238364ce1c9d74c9cee3118af407ce365d3a86113d88ec7fca863684b92589ed4caa88f211dff07587dbebb1c78453c05002e6676e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e69f91915a51385008ae59201da122df4449f9167fff812ad7deb8c51064312f5a1ecb22b5e46914ec1f072d9d22b6483ea8a70e5e1761b8c9a785f4f729bfebc6d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbb84b2453c554bae8edc4e20965c7a138eaaa8497eb3d5d709971dc06a309f6fb090fb8149d7ba855fe1f2b2f17bab765e5f296d49365223944fe7529038254ac14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4c7bc31d42df70823594839b9aa70a4e74169b3323eac1ecaf87a6a034990b806e5730c59f981af6052c2a0f1881ca0f550a01945198ec96897a2012c8f22796d01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15151fee4471a977b39d7a7d865c994b29e0759dedb43998f6bad8fd9297ad3c179641e1e2c2adc4236326b0b37b4fdd7478a6d65291e20a5202584cd7bf7b2b60f58;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1795823d2732976773b5c123b9f7275600a97ba71a2bc7db0363ccd0d8acd31ca3a94bad306d98478d295d1b2193e6a577f51b69e336172e71cd6ecf1e922b5a6d618;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c84737ec9b45ac1595d7a32007e3df5ffff7dd7a6aa405d8219290ccffbf72c0dab4e1b7c2c1c32ea39c863f4f8a7f73d2d5f22fe5a9f9bfccc332d53a5d9d922ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7d6d30f98e428c93bc5daf816aea6e94a6bf46862aa77797ee520bbdd2d0b4580c9b95e4c3560194e70483984101e359b97e7c2c4aea2eb1d9e694f8c11aa9843b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec23384353e44e3884bf1922c012081af2fc9850f66d57fa259c7e5c7697644f0d0a75eaa14d447c93ed4f4b97fcd5a2e1710b628bae4c1ccfb3f191062a712338ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c01d9292c2f80bac25882e96d18f6bfd100bfe4aa7f6af11ea0729be896371400f8a16cba720e08e24447ef4fb3ffaec0b8edc56e46a0ca34120eb20753dfb34b667;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16568efa605f29cd605d1c52479564c15d7709df952e1f66e2e8a268c57d2ca6c4940426cc85a1a4bb93418e75298b50a82dc2adb9b96b54be69d24489576ad505f14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcafc69be87f88a2236d431321e8d732b6c4bdd52f20159d8fd02558138bd63014aa0286b5cda6e710adf6a48902e11f36bed8e9a1010ec289f11240fa7e8e28e5902;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103e34e46a48fe0f68ebcb76874b0f178af960f3b9feefbd9240cf29384f9b65f009fee5254a9583046908e30cd8b5d1c89e3ffd2e320e3cbe2c72e063c983ecabde7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c44206c847e28452888caf4bf0e19ecb4c23f04fc1148ed24eeb3588726fa2ff807361e6d079460dbdd8bc1b6c0e265160737ac07ee80231312dbfd44f9c07f1b99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha72afd6be9c60f12063a80df560a8b3ec2a2d1430837fd8f0177dd239d77ffc5c7d737a2a3bbbc903001fbb428d7b937a6c309916992089558e33f1e471f62ba6457;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7e29e287891bb94439ca81bd8b7c0b7f8dc33f415389dd46694d0eccf6e9495b6e4059c4eee1545767cb718959c8071169e2744888ac802b96190e86907a6ff2aa2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da4735471c0f4387836ad7e7d6988b56d4b6d6c813810a079f3accfe51abb9e37d575cb7b5d155f82e6c33f4216502bf9fd6c1c66835b028bce9b22781cc069d75a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habd5bfa6e6aad307850aab2d44f7927d7181756914f03b9a8600a5a4bd3b93f1a2fc8e6790c6dec0fc1d67ae68db5e9b7e7ea42617d7d05ebbde412fc06b133a5a8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13730449529ab59d4dcac7f2c46b015c55789aa2e05917a95057f75427a854df4166c3eed83f29fe70e7d0148397b1e24e7e89e0e6aedb9c05430938e33e618d9bd9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9f98e4b797cb70666b889fc647992ea804938ca4d7f478f4dab78fb21ee7129de9964db089c767bc199391acd9932568f0f7ae43f278d1c65759072fcfba203e67b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14790ec5b651c44eb462b718b4fa0339a1fdece0595217c8898405e280b91e1e6b3ab6d44d14ef30fd8e44b80800f1c79f48cd44fd38c293eef86adc6386af7639c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1fcc27067b317d8e32eaf0a081feb36f41a4e02b93a26b9c9f8e666b6dc9cf321ce7778d76159b2ebc756cb6cbb59061dbc6886163abbb707dc4ad9226f6b88fb66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cd11a5ce806ae1c3d438ceab1ee810254eff4ff3c6602a76eb8b8b2409ffc6afe657944857168b359f51801ad9b02dff6936bbb0d1e311b9209b8241ba76ed42a84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h994b71bd6d5fdb917069a5a6f09a5f7eed989934579665ca6981d2b94cf888f9e4e34ed29b9963c9603d632218535e330b5beaf5fe715ee74deaccde737551a673da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e27e3c77c83414805dbca24869341f6de9663cd9be06f1fe94335b60159732aae11a26ba4994a2986945e6fce0fefca2d2121ad7a7c604db9338546848f557c0d46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4faa2b4a915317edec5e77b58282a21f5f16805821a7430651a9fba6ede8d10331f21f06065494d53c60ace09a0e300fea96a40c77a59eec11f3439201e1b592c6b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2c5b101b2450d0044d227bf6f957ce0d7922cb34349a23642971e13db9815c82598c83378c4eac4f06b2152cdabc0937704ff1baf2a716a5a6c5d056ce78b7c7a48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139f2a33fe6ece6aa70b9e4dab8a2e831f0db1766870c00651ed55f956dc5cbb4809ca3ad642d8217a69f780a6375db87c2ec56c3f88bc82366d96bfcb550309b37a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h925438d9175fb8acfb2baa8d10870e83ef8af6c1fafea0c00db136aa1ce98ca44ff7ef4179d35182b4e59f71350bcca3f6153ad9b37114c5cf40a0e673ab70c36243;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83f889211a4007a9aa5b8639e2f88f06ecc39b2504cce9cfe1eea63bfb0ebcf8e8dcc6dd89d845d91946e94cef0d391e12bfd0d961c333eebc25e65abff1055d1396;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea0dc7c6fd795ae663f675fdac807af5ddce8f4ab90c966f51dfe0b490cd9812204b5b1e4f46ff3a3a0c658db70e7052a3cb2da011f7e3bef219b9f14d582e86f740;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef34aa0b90d89eb48a813cdada97a442089e6ba9dfc5d2bf0921d9ce4e3c8b78efd4de998d0512a945c2aaa0bcd27d2a90364a8d76e554b53ad88ca9b6184e55984b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h493da8ec107f8bc9a463ab070ea2cbd096c99b892ab30573b216233e99fbb2c5ef34bc4887c1d6ebcc1a03681f813a443d6d39ce944252fdeb65238b7285ca18aa35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71af7e0b682a7469f17fb14806ec88a2bacff5be999ffe8aa3301ef46408c2e2db8b322deff569bd94fd93ca172afdd05aab7d10f2f54717f88d2527ac7ab6199cc9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196714eda72cad280ce60c481d9fe3c71a0ceccdca8e7299bdb1a38e11fe432eba26f1fcb119cbd5d7b277e66fabf6533a053441e358c8ff862d03a7136ef6e4c5d73;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4dc95987063dce3a4bf92a315394c9e5a6823d09d5ff4b5bd8914b5b64b84609384c711687248f5ba0115c61f4c85734e00387bb1e5ff093ce30b57f4e0ce9f48ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e8ad7f44e16820d5c24ec2e67281d999fb8513fa5cc1c29e4f56a14030f5087b64403e24b91fa2d3a2f71b8fb633923f955f31ce7c28bef7739e70b88b22d5f74e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8673739f0bcc75d52f6c9045ebed6c2a959e95249dfd34d92406dd89594a98ce14de54166c48493233ea4f7b606b3c8a5630423a8bf70ca4eacc68f1c8b7433400ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cda8f34161645c61a2412acc0dae58215ac6a92dc852b72b50cefbde11c12ff7eda60951372b392569c3f472fff83e88ee43ca525a5186f51a4b9e87eb760441b79e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c3aeb57e5031fbe170c2162ec2bc1cb2c3a464771d30f7acb796cfef206265d19662f6b0dd70368abfe03a003fa0f8ef776532eee9c52507ed332a05d751d55d3c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8647aeac06b6c2a8d5ce6702a6b180145a8aa69e69c27d733595770ff3226131599e16f267f9edb6fe3387493308f8bce172ee02b9702b91db4c7ac06d9e3733e0de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf8b791db7fbf68f3eb570f2357bf138197ea7f7c32eda9aa75f218a9ca84963c368bea7be2457c03bd74405340f9c675f2a089550ecfa281394a7e46a4ffab4701a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179c88a9b7fc0c2bc8073659b77fb45eca90c59c4d03be2114b4982779b27163bf3a91ca8b6009690ffb61653e64b4e07a08b20cc73c9f2fe0a1e8d5bcbb18472db1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h471e7b05d0a96833483a35669473fd92fb191aae04fbfb3f96b6a06b9a61cb4e3b482a38e4d3283d09a796438d36829341cb0dc9cda33f87905d4ab9a7da69c1aa2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf34e25684a3b577877b0ac6fa698d737ac621e3a3b422fec572695e9a3fddc869ed75b84758b96ec0aa9e1ed08d9e9c31b277d466621566ca8aa99e577e4fd7c004c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf74d981ecc66ca33ec95d0f9dce6aadc18a0a9699a9d8dfa7d838fc7f81bfb3e7e08977a35583a79f1df8bfd0b50fd47c1f7f8b95bfe0d948d42b67e224aeabbaa59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151b9256e6d811b315a9e71e1a7b19e714e287c1efc320972b6f31e0fcc3e2dd4960c07a9ceff3add11ed61ed91fa7d94a849b914892aa838f9474469b159a440ef39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf80762a7312b4fc4126f3b91b96b1003de2805583b875550415fd777491f6d12d92bc9c598994aa00915c3ca5281f62b9037cc8dee9cfb343cc51348b061de53de8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e383f7d9f421c1fd41f585a5d6c1acf9473ccdd41fd7ef54e189fbbe39d5d74005ceaefb7d7b53d04cdb242035a844d2b86befd4c877ef7aec3c46e5582c1f919c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15035bbe3082554d9cfa3b274ff13ee09d0fab34bcfe3fbe757f72b65ba46ce79caa30069fae9837e2c6a7c093a586ea604a4e74a5e267e83e7e8885dfb11b05a5143;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1446e515f036e1c669a1ada2c5d3bda23a8708bc00d3eb57d54a4a14b0294e0758ca068b2b63d52970414ea0fd457348d8d8b42eb677062f13c7485b7bf4549e94174;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ebb81465f5ae59fa1e4731c8fbb16f271d184495f77225afd83ad832a4439ba320a864670d82bd94c2de51902876b2456db402f161fec4f836da9e9e48854b1b79;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4308aa7bdc12bf720e06e64ab7c70d151a32c26876270ed11dcda2488c7cfa512c6e35e994e0897ee1210e62587a43d93cec86ad635cc8a6beb9b30255cb1a1aa0b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b6fcc7a66b9bf9fad679846fb8f6c4ff63cdab2d9a01269e078ecb417c7382e0704c79d3d7a4301f25ebb6d4e3b1740b3d0b8b5286907e0f3ffec88676624a2069f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1219d8bd19cdb4b4ea7f953474a40052d99140b17d796b34eedeada056d9fecefeaab944305b8d179a57de8a61fd373a479d2ba21687868a61d17483ed2be4082df4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42e72c124e46c1ac666b6b9b1320231862c833619c8e6561d749ef6c612ecf84f35b5f8689e12bbf75c4b5a4d63ca1540173e86e55cda5e9bcfbd06b8cdd7941878;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f570d98f1dac421e176b009331c30d870ab6b24a6020d32bb7ab5c8452580a6c125c4aa07a8202333eca34682fa458da7394e78fd2a0dae47580ccb1544f4d63169;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61824a61c6929dd720a8a0eb9c162acf176f8db48a9214378094392ab8d06d5ff1982cb5a7acde36209ae47dab4516489c3aa0fbee40d983aa6109dec73989f23111;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f19900ba79ac0de1099ac3a8fbb8e022c03ed9eb6e1445ff995086eae799066612dc80e8e476c6837827ece25ff3a19f0fb003a4c79ef6c9d2bf88bb1c203b01026f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1400ae15f8db8a3b1b5d7cfddf93350771b30c821da603d809ec8ea7f7475cafe89142d9575fb3ee6867e2970f57a82b8aa4498934ecdc9b65ea89b022040ff5bd79a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152e9ef94a33f66f3b81d50dbedadcb4fb306a0f5d062a5299accb38d1af1e446ddf9dbd2c2eab9f3b0bdfa2f4263c8c91138c361ef2bdc46d3771eff1b45bc56434a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7dd2cecfebfcd4ebacffd6baca0e8133f93000c4af17bfd6035d5690748d3a067f7f82b9f5e684e2fbe71b205a83107410d14296c03d8ba05a7a9bc89642378133bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c11448d65f3680639418d77f551b4561523b35a21746fc1a892c4c23fb51e3ff132c16319e5e38560edabe3e7583012ebec13e15af32e5fa4257f0c2385ae51edb6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0b8bffef418f7b2e7d855add30b28fdf43d1636b7f482c4dd445748c0e0b06c771f570e1f315b95b090b06101264bcb044c3d66aed0105ffedc2e36259caf0d863c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e205c584c82acf6c682dbf004441287e767905fab7267a4da41d010d3de55f9f99139be229b447bf37da8cc57a60ba78163ada12e7e76f6b4b80136af1a25e580ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb106c76d5fd850bb23c1e9c294ffafa543ca2eb0e87f48d95426171f66ce7c3819d7e0ce5b5b1ea13ad06f04587f513952c5e4be753e149d167cb480b4957cf0772;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154b6b2671ed40eb14c088cb0ecb6f2f289736e6655c84d41aaceccc1cde3cb96456d8b80a6e7baec8417220c14e2558394548c1fb58c5277b5995cab87b1e8c52618;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h827b02500f7b3b0631c555ddf95220bf7ff31e15c56da024d9f9754d80b777ef325a1c09addc987a15f22342422bec6d38552dae0a418c55781e5d5af08a04281982;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dbbe9e08eddaa46275278f6a80b3cd766ad74e8268c187c29dade908f17ee535f57f764dd28b13620f377036b80c931623255ac82bb76d7540f4dd30c87f545e49d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1577de5629947be9453b3e66b877c24729e6aae67e81c498b3d409b9a980c1ac087fac771dcf8cdd67300654586c50cdbe9857a1b8b55558f09056a539c3b6ac01240;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafc22767d47b6b20e5ae8e1008d433bf2a44304f65f4ce10bd25f371297f49c6a202ef8cfa68ce183836abfebb200b05508c2800e4f7d89280065ac733c243bcbe4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e89c865720a5a05455b62695653d3e4597a098de1ca72fd5acea8c5373eabb791e9c9285ed445ac9501af69cdc616b6da8df110cb1f32d4b30020a61485db82d17e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad95c7bd7a68dcc1325e1c276ec94b814bcf68c3cedb1c6f02e9d09cd5136eadb254d2719d71e933bd92d13611b76e6f2e39c2499e1bfcf422d3374c2d3a085a2e07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13949b857756ea13fe1695a9f4496ce5d7f89a940983c8a442ca631d277bb281294a2be3ba6bc07d05d70a28ae7c689e48c88a1cb0e78aca83b356c5e83c604cbb073;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1d3d5ec848fcfb5e4bb6f6aec659ead9c14d15b21cd9b46720783fa93b2843ebc03024571c004b6c2e7c753fdd9a28239b6529ae0676a69b9bd2483a165c6648266;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118b31e2a3f8f586473117f1ca3f146c47782f8776a6f754e30a482673f294067ce05ede272576475261ea1db38400ef5c4a964c9f7a484bb6eab9711ed524b7603dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154a47729d225b1145bab700a822fb068a5f02745cd2eaf9cfbc809df7c82b33a2710ec9a257d244384b6bc4690ea598d8627669ead85970c352bfdb6344d4d17ab19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc100daa07fba3916bc599c932fa735d54ca91da9359e45eb2f876afa984da5d8ec710731061fdc15dae41a76b601f1792dca43d08bac77ec03687385225d0bb43d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17356e4d8dd086cd180b1c4f71ef6de91da7a969ec48ef6c81286af4625a9dc148dfd1b960597b0bf62c4035abf950703740211994184c4fe889c374fb99519280497;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h288e8ffafb3b4ac559f7f37b74c40cf172ebcb60f37a828dcf3e3a6bac255dc7160ba3f18192e75bb1b686e76d416918b4a0f37dbf455422522c91f8f2af5af8b1f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f221c4e5964efd1c54d7cad33224a6a4045e746c6187368733b1b5a196010726d7aca4f4ae1411bb2456d59a033c8f42cac050b1757e1dbc8b01674439d12f88d5e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a70c06c14cd9b3761d4615c49b1e58d7238c08b7f73d4d73589ca55a4ee27dd0bab01aa70f139c35f93b6aed7c5ddcaf56b2a7ae2c64d49c8e931468af83e872f38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd675638cdae1ceb1a3dafb72580c790ee8e55ca04251eb4466d1df489e3fd4a01a525c9daa288f72a70fa6cf0bde75dfec779381e1ee7faf2cf4a15c2bb4c2a021d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97b97d8141e90ea187175908a6bfb127266caf2932564d7c42183b60154d138e9945b5521b3463d05e169789e0fd3847591513268784ccd0e6958113d1307b876d20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b7c0647ffe14307ef7d0275ac8c9e0612a160802c7759152a0a33d26d25b99d54c3f49ee3f5581a3b62afe51d8917adc26fdd965fb03cd24c7defe8efddc4f6eb27;
        #1
        $finish();
    end
endmodule
