module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [23:0] src25;
    reg [22:0] src26;
    reg [21:0] src27;
    reg [20:0] src28;
    reg [19:0] src29;
    reg [18:0] src30;
    reg [17:0] src31;
    reg [16:0] src32;
    reg [15:0] src33;
    reg [14:0] src34;
    reg [13:0] src35;
    reg [12:0] src36;
    reg [11:0] src37;
    reg [10:0] src38;
    reg [9:0] src39;
    reg [8:0] src40;
    reg [7:0] src41;
    reg [6:0] src42;
    reg [5:0] src43;
    reg [4:0] src44;
    reg [3:0] src45;
    reg [2:0] src46;
    reg [1:0] src47;
    reg [0:0] src48;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [49:0] srcsum;
    wire [49:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3])<<45) + ((src46[0] + src46[1] + src46[2])<<46) + ((src47[0] + src47[1])<<47) + ((src48[0])<<48);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1920e72fb8d8a8f01bb708160fdb652b05a5230575216d6c6b79176cce72586bb869f26ac96ab73eb2321688712b10f3eb33bcb19c9fca1b65f883e5e0ae6ab5f4c7f073d3b074bd17319fd877cac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143c056e669e580b25aed3291e7d06b9eed1e89d6bd10f8a32fc300e1510939872bef0c59cb2709c3b0f5bf311a48cda6fd787ec363019066878209ed9b7b3d16cf5e6e99150ddea96f7d2a3a82a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8012b7f21618347a11be26dfb938343f966d92cd43ee3937d083ba1c446be25a3b1cc6e4109332cd4c1470bafd83fe55be8c49d594529ceadb6e11959920bb79e00515ce846d84632dc85bcba2b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10bf1b2e6b2599927c3a2750b7e4838ebaea57801a101616befe909d95fae6f4ceb92fe7587350afecab494f5cea8c5a23fe45c49ffc4f90ecf5696e201a3cce7ebf2889b77f1020e7e749e271eaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13603769c75f4d2ab3c316c36502fd8f22f2ef6b8380f3f6efda515dc2f2e8558ee8671618ae74170f31021d14dd4574f1ece11417ac8e2cefda88c59e626282c4004f2ab93177d4c5fffd9d2568;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bc2609102f920d360813adb2ba29a8b4b745b33ba522043daadd10b05d93db3c6c58049632df75fd5f4b346cf0a0c1a739c0f0f03e0bed4ab7357d431ccb6c11770401d7bcd4f2ddc2bc5db3998;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b22059b056f28a2b0b6f62717255576657f5cca15e1e239e1ff6f6ee2b1ff1a76052b956d96325dc53cd8464f54bdf2e1b2a46c51f6bbb0547383a31d0d6d9df15ad28b22351e3dd4804e0c933e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35fa7bdd3b2610be88e94b97b1f84c07e54f11c3fe48923fdc61c93a663c1c7658584fd49994f9ffa872630997236a4e5dff64af4796135cac93645698a82b8bd0f53f14a16aa0713c274733772d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cf92caada7248ba48dec41e05b8d73debed70285fc6e5509482505f2af464d52c3a6a45d2bd5af8cc834d5c4278c784af5799f0a392f87b83673fba92d5cb65fb6beca043a6d35b8af8ab344dbd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h151669e2e15364a799ef0c5ce5f9d71e82aec544596f5421b95a611f088e2be59ead99810bef70c8dea93654f0b56f1b7864b76fb4055c8be2988d4a8b9a2a1a8bc053900542b7218d963889ec8d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1098a7c38f649e1ba709eff5b9eae8699eb2a0eb5992e191afdc131b2720804e586d13ec39da9d521f6482138a5f50639c47be44587c2a420f3e8d68325779c0636871f3aaf72f8559e172af2582;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a2b01d4f8e891ce6cb4bc504276d6f95109a2964ee4cfdd225c55b6f58be4d84fa1deb3f6682a534227d7b240eed49d145e400d93c4171b99964010fb6aac04ff9845d6841fc814577e60408be6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44fc8b77f23304de21625516b297d0583804eb3a1d919ee515d2e5bd9e5e6ee0c1cba49b3610293b4e9f74f96b77060b463033f4a6c31f70a9c21211f3210477ef8d80ead9511c990ec23f0a471b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6c698ad89cdfb60db5bc83e18e5833dfea0184803b05563a5f3a5203cee668c2ef50dab903d663aa5ddee23c8dafa6f2e00348b14c2094c0ba89fc8c29db1dbd17d5c2ce90266c524ab5de5d59d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29c52e4b1c44797402643b0b184729b657165d37dc61aebbe0ae537ec03a8a301c23da1084f59bff6881f4ff0695b9233c86b0c45fe819afd70e164f97459b7de4f511aafa31aa0ce13ea4d84991;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcaa260697960e5b8fa8f49fd9fec23c612290bddaf361a63b42d47892d90af6d1809d649b4eebbc159846976c39f5ff73542ecf1f46166b36f4bf8053a69fd980745378506b75159453ba1aa48e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbdb469a55aa95750a480cd5325ab8604480586f6f7aba411346254b73d19ac461304f0ccb978c3b2d68e3d997438ab00c5b743f0d07fb1cc548499394ade5ce9156eecc60a090c2514b39342e2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180301454ad4fef263e4c4bbdc321ce353bb9146ea6406f0bf0b1e33b54d1b37975c2993a33eee0662fe7fb85a4fe9df064d855cf686f214fd14e6547c016e535849ec3319a2fd8cfc3e03f080827;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c56354cf177bddd16c96d9cfab05826dbef39e3dfe4bdb9af9efe1b6474c034bfd88832117f536320c31696ccaf71dd84e707f2dc0104d965ce2e4a848c124e7bb19c91f221323b95f41cfff134;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183a1c1c7eac473a1bc1e9bc5007030ac75c7b48d22f17b4b95f1e372074ea67c6eb0b21de4518116cd8ce524f82eebaf44ffbb230af6ab642d6f2aa1b59d9f99bed59b2528f907035443556573bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1085540f6f25f25743efd16887ffad11eaff82a9617c415a679f0560463d26e9871f3873781ee6d021f19c43fd411a3b3a12a2fe2f59f4c73ef3da0e0d989d1e47524bc05851350eff59be87edab0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3396a629b514a89d8946f14508384925da6c5115c4345d556d8b9e7517ee378033258a49a82c46be2a88df86217f16b8c984db1f3e237d3ad5c9549d673c7dd66304db1e07630e9737a3b797a929;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e047c7a58eb5049fc28bee54539d9c5f04e646282b22f2cd168e4241d52910289b45ca8f2d0cdafe62fd7ccc444e2456381c1fc9cbedb462548313a3873db77fa126de874b3554f599cffdb8cd3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbd52a8433c0e148a934c4754d3f65a0a409d96bf9e884d22496cc9f86b05aad5e53b9ba99fd2326770d9ce672359f80ca148aaf5d0caebaf328961badc6507f1524ebb0af47d98536085d74be8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143fa482df8d834f16f2cc0949d84659028d6becaed3c333dc0c5ceca170df119ebd368f73ae93d78c8637c9ae79d698cf5aa08088c662a59ad48d12f38b549352f77e12e4163f000f2841c1f8c52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72ab8f2df92736a264be5493850aa3c18b170ab9a132d431e37b3b270f1f3bad684f14072c704d01d2f49cbbfd15c7affcad05255fd5179bea8cafd9a0c787884db140ce4a83b21445cfacfdf532;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e7e1c11539a460c0952a8afa4e2740f4e9b17fe1f5e823b5b19643b7df7c7de68045b435657798a4245f8cc4ec9103882e517972a2490b0194ebded4f33b8e0da42e92597f2db3e088f3ab4ab09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2264b8ae73f9487fb138d1a0465710f709479e8521033d6f8cb10753d91779dd3478a8f4e88a6154bcf08803d80a620ec8226c1cb11ce25cfc4e9b6970b00b3679aeb91dcf069f5cb840d5ca7b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b18ad0c4e58215ac72da7bd0f383f2f698c61ae08dd96b24a2a214d61d0fafba98f7b2eb6948f03e8ab222def2e0a1d99129c13edd96f8789b368471070e380f85dc2bc65692e1e3f689e4e9f70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad7da3c76280136d006efc04e130fb9b017b99014f04c3b25819f69b53082967097d0b0919e9af25e6fd0c5251f2f865255b2e618ac1fa7ff941b719ba89688947005743ef1f56cc8564e75928a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcbc2bec0b9984ab6baf6496dbc4a0e46698bd8f8e81dabfd1e99eb2ea9bd2ca9565cc7957e040d19dec9bc0b049b29aac84b86d1a6fddb8514baf6c60b03586a931f59b151b04191f43d3281402;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b82c0f10859541a9fef5916e67e4e2eb41bf3e6beccfbc5bfb2473946d7b7099644794ab0b44978fd969d5d0c694cb04c62ef9412da12efb7f27f3a9a796b43184b530c727c428de8cb82d64e5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he808de7159e20603c7250eeb79fe6b92a61d84eea3105c9d54b0578239ce1e774f0bad606f8f58dcfe6b536ef4ead5b845648f54262377a6d5772da955c649b2619c9853350b440a616893f194f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2338d61a7354ed31d30e19e5b3552e8af7440f1a52d33f285f7865f92d4dc0756b68bd5e1d3603176595a203d60c5d36b4e107106ff49d907b82ef760c8846d3991b0c54fa5e46deb205d2679a9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h586dec748dc77fabc3626bef784dee27b3805b31db8f5153cbc4930718d737ccada10a868953afcaf4f2a80543804d32f4a5df89909f02da0a8694b1efe3372b5f1d316dc095ab7da38154a0456f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b64409c58a4d0aa1004b8b9254f5dcd8421d0ceba584b12490a475189795a258a7743bf03da4a80358717cb6a161cb1cdbffdd863d2851f24e5155cd702f2e75286b6c5da6fde5d87fe4e3270fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5336ce82a1925b44e569d0086bf013c931389f622b2fa5cbe5c5ce7d6bcf9d35f9e7ce45cb59427620a19469e3a1347888e62e57125330a80ba2ce6edb77332041f36dc466ca629f00766822eb0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdbd7e36ea9c8f400a5748e058d36b06f63c70a787e7504d6120393d73aac61740f32f5788b30ac671939910ce20103a7c8364338aefd98d59e432d1565a2c566387dad55c95c56747c5845d973f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137d31495dc533ab369a7eba865adac347bc969f7a1f1b8f9cdd35dff15b25c5537f0c20435d421ad7a3174579ba7f7ec5e8a20e2b3d1e5d40ab598eb10d77f3e856b8320818a78d6ddd37fd5506d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e94d0d3e710f57c9832290f01ac3f2163147d30d744663d616969318ef79167a8ea7e849896493853e9358d07d25f3dd98413b01b978cfff3387eb3a94660e15c72579b9236082740f3c1b273fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12947094b045d3b805d0689fd449dbaf2f012735ef060ad85ada9a58a2d1771c5eaf9e568d39f4fe160fd477ec811cc2ae19eefc4972e31cd1e4823e277116e61194a1d0b2535026da7451ca64c28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3bf0399115c627430ae8d736d639882172eba9adb0513ede6e1b34486dba3565afaba9781b309b0d779806843343757dee28f7a16ac8ba1e31ee34f21a500bf94a07f7db479438795822539fdbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f68af4f558a34408e8fe29c968b2cfefe16f0fed3ab7a4729e54ec6487225e9bf6bf385a34952592fe25475fcfecfe51a690cc91cabbacb612cb67634489ad3f6d70f91ef7ea6134cca00ca59586;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137e906ca3a7e98591e2f9fe6382cb907a68aa467e0554937abfa75bd7dc42aa29c694ec9ca2d8289a1742b65e00727af195b7e6001913f266fa99e5c2d72b311b2ccd4af09623974d5807bce0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ba6594222798ff57a2d73a949bc23d73161ca9c98fb7469532af31e17e49dc8f98cd1af1328455a65f68954a6ff54292572f035ac34e462163d2a9f13e9a565bdda7066e5509e228156913abf55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa28474367bceedd68e1aaa939e0dcc223d59d1aeac07ec304cd05ef59b341781157dab3481613c1b226dd28a268185a16ef8ef929cf01ed684ffb3f085f72b21b849b886659085cc886f20f9c90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5730e52f269f618d24d96968766010504e441acab82284f22b625c5e2b08f5ef6e367c5df96958b10d61a520d7b3ac5eeeddee8dc79f771a4875e67123994243ee4930c1fc3890bce737de1e9616;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hccfd8feaf5bfb49eb5110d88a805e463c89a30fd713d6389287a38981a26ae163e524fcb05759a008765ff0fef0f581bcbf41a0e10953a1a4b22967f39d34428d2da0eea52e9e75cadd45a2c50aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e0770fdfdd56d0e1aab9af0c410e37d5a93bd72065664e1c156ce08b3d9cad2eefde12f13ffef7bc956e254c57f25fa80320ac7fed9ef53b28f513eeb8e0ad7f3dc59d8f91cecb4970761a52b55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc823ac1744f5981f692991d8a184679a73a32a2a7bcc5bedecf7a4ce51e38ae7b38910ae574b05995a59889bd7798c07fd29619b1b8ecb5dbc7324ff9b8c6f89b18e12447f02ae6c6ec80e33efa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc5facb652de2f10c3e6ecb852749903e682ccff5a3a51c17b839416e7728e616f06839313068f9b97f077cac7248c5055399d2ea71f5b3e20cd5af49e04ea17d1212c24c0fc4cafabdd63083365;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30406c4badaf02e655a0bc152ba926b3408a1531440c1dc603fa922f91f4dfdff50efb197150c86a90fb5a9fcb48e229dd4446b6cebf32e2398347fb67b9a06227f1fd1009e6f2bc5d721aa21d9b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaab19110f7c3931fb73b90ecb2dcc83f94fe71d51419b6d2343d29e8649c4bc60b62ea0ec2a0a32d7c0c6fdde7eab6e45dbcedb355a97f64010f516a7fc5e76291ae7a17f7637b484aa8d51c1ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e54406f7458af9a40f5ca8a28a10dc223cc03c1c87b569d905697085f768f612edce064dd3da8329a2071742f89a039446299b512dd137c941bd1d8f0d792a4a6e5a80ab629c5468cff89afc2aed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f401160439d923fc392021981eae5d119d2393a9fb9002e7b1a01d3e497d50f80b0e5aec329d603c695f5765d4de98df4f9086243a8037db9d575c2cde14f2671348a356bcdbc2b238752d0e102d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e7879f751aac25760badf3ee36ac49b26ffc31862ceab68b290e6a2683131dd3b9894d84d5cad758798e00631f6c0e664b11bbc6a1c504122f499e0973f283611385780085526f5a3d4658149f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88dc5f4c74129fa0c08f8e972f5848e1ca9cf7c72e7ddd4e1b591f9a5cbf46a39a05a101dd650f4109754cec4a39a07b32e38b1701499987ae9159a278b8b2f7dd207e54ee0b2a06814cafdf76a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acd0a65aac4a8f24057c21ce0bb2cb1cafa9e62ca4f7152d29af30bac8987a0ff9f8ea793e3d9e5b93096e34c399e4034e159d964b1f0ab7891a710ae34806535296e6149b790b3ff2f97ca4ad62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83d0cd3da28f74198cfcf47673ba0aa57e20c4e8e6510d059f4ece3845df4d8f24fe0b23c628b341478e38afd5006b3c51fe320101baeb1a5708c463bd457a609019f99be9c0a4ba9aa7ec566c7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h852da3776c8a7bf70da451b5d308d2d86e05ecf4feb18f0e374a38055f13dfc8a61dd3addf2170324fafbab2b1a20a1aa0327d539add47f78077c1b06e93b8e766b73effa0c54006dcbfcc2e31b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138d587871547281216fd2f9653c5364c4be6fadee93fe7442b53b7eb3b0f2eca45807f127dbd72d7936a1a3b72b33a772cfd7bbf4c70a23ef4714523d8de9e489f9e950180206c8210f1cde025db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h675e490f9f17b316f8f9253bb1933127038ea344ded8a5ed0688201cc2207a820c8e581e15677bdcf6049119954ac9c7f22b1da060910843b3dab03d1c7a483655644a0d7612b4e737af06f5cd4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7505e7d4fc94b5273b127cd8bf74bcd865b540451c3ef7232078221594c2c603511f8ddb82705f0fa68c928d1a214b1b773f5ed670468e2b379db1c717aefa219a94cf6c3a8931d8bef5466345c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6e2b84392c1ff982d12477b68eacdf11d3d734f85f2aaf4ac3c386725527920ea6da310be3e334f4f65ac7195dd2fc36ef56b0d5043278713787beff58648ba02f88c5fa750b8816ef7aa459e26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3494ab9141b734f7632abff510e73c8295f7d428c87f4c50bfd6d518a7caa32102512879845e97dcbae3bc3db6036e223d90dd3f6df4ee3e775aadfa8108a3bc02c1f2a42df69c887d4ded44e42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3e7a89e6c1e0633af6f7f00b2d5a5b0c9881bbc11a50b3463ab9fb5ef2515f5b334e9e3c99a9b801d185f9e6b819c70f66502b05aa80aadfaa4d400ac399f3a5601cbc6f7d50cc82eb3a4b507ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100fdb505301e29161ef8036c48e423ef170b4e4fee93ba4e4101ab7e6e75718209a03e4de5627925f635933bc29eea7679904e31084e82964258daaf280055b6f4f4b055f46a0e6a4513324d371d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b02de6417fc414e060a54315702e9ac7f1e124d0182cd33bc342588995875cec48298dfb66fc227acbd2e6ee72433f38b65f31c41f8d2e2b0326f1f1fa51551f11a33424a5a119b065cb8cf5fa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e1ed2dad07479eccdd59d57f55106501cf8c74b43641bd348afc1d5b72a2495ef290c5bacdbf5bbc0e4f04c11376b12ef37c74dfe96f444c4d671d1abfebc6b11fbeedb594f7fce87a3d049cd91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ebbe0f3c28b64d85469c228684b4001a61a094cd0e56948d5f9e81cfd1e407db65d2bab9e01e540e334ff5536d17339bb2a7b5426ab01a46a3c53e30751c2b490afe1d93488001e56888dde41e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d23432750ace8a555425f56411811e5d9649db5dacfd6906827576c8288a27172c06c76045b765c437a475b0c4197752b67289a0464161ab350a2de4ff1349fe6ca1d6056b4682b5b54319290dc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10902875ee27ae1bba35523ac0c1516f6fc3fbc8986fe8dbea00f54303d253953b948a8469cf109eaf6d527f066d3d12b4e5cf25f723fb29e7380f8aed472bacf47eb262e45512f8c0e071b05fefc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b8d9435000f13eaf2d6ffe01f0088b03043ee89ffa3b9bc9d8a95e8cd5821c48d5065c5102cd74a1e9cf2612bfb23b678389ba2b42248d891a7ec7eeac780b7e96c289dc6e806973bb9156949ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd05aabe15da50283704ea94c7c1238616848f0fa29b2c84c16ea08305153adcf1a1779744cb982a7bb00d9d8c1aa03058d697cfefe2095bddce26bfb08bfa02f01a57c6d6f22054f81cefe39f002;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74d23bb43cedace2496ae699e58d7aca0599ea6a2e563668b9b1ba7b2de661912a06e59714e2345b608472f423348964bc4340f4b4fc9060e8cd6787443a2769de9d83c4efd5fd0f3f17eb3d7d39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0b549bfb6e84f2d8bb21998bd27930d82a8b16709f978fd967451c2ab153a87f6fd7f2a0b811f25037caaf74cc589efe69284743d25913f376f4810e8d1dad90050acc9353c2081bbe3cd71c828;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14005f005c62ee4605ce12771c5b8b7d6fe65bb782787e89e397341d8d64a537804ba000097b49841ae9608b261965377ad33fb257d539edbb3abc0b37f96544d59b3c39760fe4c32a3e1917474b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h665a4b4a7f28a34f63ec65e67335d3023d864d3ad0687c1fe28bbd49142c564020efaa0ed37c057e8bf5d02b721f2d4e4977153c746e018776dacef859cc31b99ed459985135bc20d12d864ea958;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a098f1efa720a82a289363901a6b5ba642f9f70d668f4b3858315e7c0621027993517493881c97b745ad1e476e72543fd8b3ae1170eacbd712ed3dd212119e59fbf9327ddd5ec043834db444dad3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71c0d94d0ec1d5325aadaf747ded93b2521d9248f4e5fdc395cc13acdae4de34806f08833948b145bf614527635827ab6ec7f2e7cc13b80fbd09f7f9b650e0cce272268c83a00e24a112498c66f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71ce065b54a7aaf856deb7f1700b24b41e80462759da4f0336365262b7ac13a10ac48bdb1efa69ab1a97d17a1f4bad207ebfa950fc59addbb2c775b0a09e836a7d1dfcb4a222f0bee71703063d7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h936d6f63b6802727ec65bfee6d138afa25b3d5cc049698191aeb5d2b4e1744c0e37e0f4d02662b93734a006b57d6ff6b591732c60de40001106e5b8deffd7ce09984f26b8a4281de6ad593c35624;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1672cec4b70501d48199abedd74658216c513421cd1f0bf3a5a3e220f06b6bdbf541c0903877068567e05f55d6ccbfa28bf700a5b163daf9880dfdd11bb68e751bf09619c85310dc04daf206039;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc74aa03dd60669de7c32987e1946cc49c65ec14d6f66a447e387f55c3896660c38b503010889ffaf83b16abe5b3dec48bdcee7e838bfe3b9f0d41c28038bb8493f18d650c01b3cdf217eb066fd9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b30ed6359915546787578ced23dcab4c2d76335a8eff19acbe15390fc1acad50755e6e48d3a6a821e587051cf1251f627f3099ee5816e4399cac1210d99760f6de698e3c9c3c75b11fd92ad1893;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10343a68246f147ae3286d33a52eb3b167414833d4112a40a51e4af39707b48425959cd40b37192331fcd7206017c3763c21527a32720c3f9a3867ae8b3e3ae8a7e844495087bdfb428f5f87f440b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36dbec5fe101e307f5be95d15bfabc7d361e4e97a25674d1d6b1248e9113a1976f6b0780e629259b826666bc2c8f5c8141215891bd473600ff398c5726dc018d60ac0bf4441f8ded94bfeb48b7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68c221bb474fb189e842e328d537bc9cfb3e5d08b3aed43f37ad34c41f75de72df7816056a27d32c4d0e6a164bdefbd6fbdd55f443b15db529b6e964200733d841ccc9bf5b6f6981a2a8ebbf993f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa113d6f0fbf8193ea981fce7a57427b068e876cb3c061d709894a9e042ca01692816dcc144ad070af7a77cda09238ca897e03e4cca234fae83376f54d627f22256396796cbb417a4bf1e41d0e90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1714da0510103d6ca537c0273c639d6352bdd5d3c3945882429188c6a845a8da2c08d56368aee685df0e30d884645ac8564d1030a91b4aa254aade669be1748582b1073f8499c2ab2622b2bcc39e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b5de34f2509b28c09e3bf9ed9ab5d73b3c18f58c2547632d02cb6f99343ec5f9014b4424ba1a9cd8696afc5c2f99fcd63486328e3a89b51d041e9f3471fe1d972be7df02c60a92a3bf159eae790;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12eb3752c7f2c3e61f5c365589df0457fd26e04ab1b5b1f5e0ee424a59088caea1f433edf691ea59b735270be7638c44e90a8e03ddee753288b3b529f43abbf41b9c47d2a391bc791d0954de0d8bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ce9297f565b44d837cc3af0c17553acdb49feadc3a958d8fdb5a880217ab0db7dd89fa7327210dbf6774f20bcb2067cf0325f3f337afe4c8d2b5c359b5be547f4a57658e0faacf0e5e76b6d94ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd988b31eaa088f43b279615cbe0be4dfc34c1489883253615b1aa3c3ea4ca95397d51c4b9f09f5ac4d1aff1bfaade1eac30bb0554f3455b509570acaa6cf35e51c05f53d75ee0863eb190289996;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5eba0ee03ff658890b10e936e74950c88747b3bf3c98d195ede3fab8b135ca8214b3a03b1a634e3167a103b2a7b2a24535ecace6137a5ced9e967e2d15e7c4f5568741d347eb36335793097ff607;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f43883b77d8d8f4ae044eb56ebebd4b16e0eeb316fb395d68432601a1ab4ede43b7308ca7f010e24d167ca73cb25e73dca7176a620efcc65121e6d6c3133a27279e1fb6d7a9e7e0468e345cab194;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1675b769845c32effce0c5b2cd575f957feb667c6c438fd397ee205cc4183a45f7006205cbb3a53bb84692f66f2a11255525f76a6e4a0a4e6987301689c33303080963a65dd6831e68bbf46aabbe1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0e73903c6dd9377471475200a4833066790a48af7f508b873a1c2986c85b93525f09c2095d88a67747e10470609a06f52627a1d3bf584bc6a5768f81cbc2d450c5a9057382fb80f47d750755dba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188a63b6581a1f82e4be55c863802a02ee57514249472be77f59db27239dcc46e785c5cfc10dce4808150cab3e0fe8a9ab6187be738e26af9aee452024861f9f4f68a38d8d0f2b17fa0f239b84983;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f88bb160bc5bf16868d2920facb79b8e463b1d0c4949e720c0f8f07c41ee4cc7fa7775ae9855d3cb92f2c499a4839750cf27b13d421321c08e5ab1ba385a7ac97d8a527673053fba7140db5593c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1ef7d5afaa6c8f0ff21dfb4ac9db52f713bae84aa5c2a58c4de6e8bacadd2433ff9c433e489ac43258557ee9f654ca96a1fbc1dcb903a850561f1862640170a852bd22926dcdd7e8f6be4f05b06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb62714c9db1608f1e2e32866cfc335b791acdcef365f2441ffe81dafb6cf875928004cae479590c1a26300754390192b445beffb1d9758edf1732785ed279290a2a96c487d25df2b64279e4f0160;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e18becb6a55b9a12be9958647c0a189603e8af009f2a291be138badf9ddf474263a63720423f56f2577342cb1b76f1fe14383f4d50b777f20f0aadd8ff14fee3a976847c48e866f605246089ece;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7e6eff920c37e85f4795c182d643be63a22d37c7a0c2b13d3d333f7272887cabda76e2d9e9002fc39ad8954922f48e848b47b5f9784af791a34865f9326a268da0942921ae536bf356cc971c9a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d4c6ed0a4ba509d31471f31c58706845649b2ebb076033fd9c84ccb16bedd395ff274c3211b8fd6af68a53dd21638aad709e737c7507555359f104457ceff4e54a9ee6cd681c1584df2181878f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9cad354f960b2d62811d5d6c16b1e459596c16e4a37d5a0481f38bf3bcfe7a3920f99d8d167c57f743da221aac5e0cd0f9ffb983e61cc437db665d80352f2a42c0ea9c0cc93e1efb7464dab9666;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2d8d78b122e20abefce8a256c9fd3d06a81b07def090caa610df1013feea7751537ff0b7fee133adbb290ae67817c1972090b8440ba5afc90cec68bf2c4d170d9b1e89bd2c73cad8cb849d7c403;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fec6479ed159cd757226124b1b403934420f9ac4bcb5dbdb20a916210588898fdb4cc4cc2e893bd6ecc497d475753e796e2ed9709d1e9fac715debe9ea5d2df71cc406703a3d2b435858d2d6994;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf078c079758dbd6097c547f656c26f9030360b970d42a2383e1bd4c0860b08bc4f8a3c65c394f37215edc6d176cd4487694c1e7e194634254123f908d8797b50642c8e8cbcfac57ec20a885f947;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11dc097f9a380fb33da33a0e676cbe9b3c02692d80037a326200113f741dfe349a707cf4178287aae8a773bbcf3fb634bc6ce0a05448849a90de03ad40d607e80e0eef3c7832e4f3b25127b9798bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b479cfa2cafb54269af08528a97df06b6726f6139c113f9c8c64c083b78995d7615319df1be50398241f00144ae31eb39b15895cf1152250688c0afc66cc7170b7c64d3c403074c0cd56ac45686;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h497585e8a7eeab51c54d1311f2541804fd6293024c1ffc8a19ba863a6bf0f104091ead9e5891e41ba2b8e051aac412752dc02b35501427d46ba471876a4d4e91470405bea647dfb0c1188358aac5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1000337fa92e3b74dba700ff6cbdc15a45160f1c7e95d56836018c8c53a8803e41cf2e60e0f93d3fe2bb46e92190f8129ec39cd45d47e4553951cdf4b9a7da3add1c58ff8343d53dfa044320b9d88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4e0df1066cd50f9a99e8f2fd3452b2774c29cd6598b194a94ec4574a8e6c4e7da03e040338e05e494c58c63ef2707c5a2a24847b024e5f8653dd868ca9e8e2e4820dd30066b63bd06cda01a05f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bf041faa3d52484cb70d376d2ac59a838c21ae5cf2a6a6d847cae490843c73ed219ee430fd46051bbe52c267918775dee3127fce9a9b1c282ebfb6709e1aca722d91b142fd4b7260786b24dacf1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187519f8e8ed180cbfb18a2126310aa630c3ec76a6f8b6574709185170a7d1fa8d5ccf89349be96a212642b8061205e89e705627d5c52e32e827a465df60aa3062c8b81edbd5cbbbe1d03172991fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d98b6365c2e15b0afa027277015229a7a5bd5286b7c378cc5928658ab6d0371fea0948768f950e01c2a97bc08d761b37d4f8b649d0733f7338f46eae125619a12a3a03a7e8b84307db1a9bf97eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f94e06b48c9f3846a8a7edf43dd429436c27842ddaa9e9485c2f8d1800645a183347cb9b6b3679f321eb3f30eb6d44219626657ed0959df15b71dd3765827d5f12aaebf464f4b24c93aec347ae27;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5c50aa7fcf5123eb4d1f9def733298827cc38167549df9d34b31b580144e3df6d24e9d1aa3f7f64f52af9006ef19152faaf3a698b19e73914fac7312f169f43f5ad0410fdacacc7557e4981e2eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be36148dbae9224419aa01df651b3870c3c36b22062f6b3e2c440103851fd9900611720efd1f09f48be4e68625faffb57e56e50a6863dc6d5a4c7ae7ceb49f5207cb10be645bf9e6e5adea4399af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef682af14d884ee95be84ff692b719a09d7539792442986e384c63ac0580999c70e0866536e7772d42912ce04c1a54fdefe73fefdfea981e2b56d7ae0f87dbd5179cc35b3ab7eca404070165e743;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8e713d8654a5bc2090d3e5fa70588a4e48514dc06af43a916f1ec3bdd401e383b9de9ee1201285555f7acb6011f12fd7a5f7a01ced3e724c2103d3fe33d5a2bd13505827288e359bce08ce5b19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf46ff8c82f38efd97c266f3b0346c707c14efd7bc7498a1bc6356c117fc61872394851401ee6bbde7c4e3921d31e866ce80b47b803b303a72d01d47dc8c756f4e411bd3c49be5993a2c52f5d973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd278a2b5ccb03ae88a299c7e51cdb562ed7553ae4221d0aefcf199ca10ddec4f5e417e467c8102a06eb1ead7fc86727ecfcd63d275ea01efc75e39243b1eac57c1a34e1736a7e5ab69bcc54f1955;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b4ea508ec03208d717fe745fb0ea512277358d59da046242cb1815b4379848c753e903fd335263c6ff354194f060f03eb4a8e69f59093673d537cecba89fd2efd7ed3eee8927fd34c207a596399;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8256e6f6dc55b6f70defc84c8030e20d09a1cb74ddf0defa32e01f1e0fa40defff7e455fcc7c35731b2116e0cb354697769340d1f363db5914a461b72bcfd9632ecad9e4972a4b9f2262109cfbf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb7cdeb5c2b79fd6946d3c50dcc27c6ed2365cfb5146de448d92618ffdb4a9a9b9f09ce6a471b267670e26f1922a2f9d05a3ae2984e0393cb9b485c658fa044002241f7065c8947ee33d2c98a066;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d5923fb79772ad666f8ed61186cfaf8cc98b82bd8efe49dd778ca4788e3ac9cdf27a39f02dc8e61c6681646fbc21f5f9b780876d58736d5c0aec0560360b8d978d1846960758559306f1e2f4658;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89433962186f5e7e4301bd161272655e6e18783fe69b999ff61d28b9017420383145b0721de015c375cf7b97c12cc9dc0d4a20eec77e8e1081749574bec581c380108338b6bdacf5dffbbf1503eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c985571e2ae2ce6fff659f7f165f4c5da251b6e7a7f7070431a9256eeb68f7f493e686b02420029bcfbd9754ed9612ccd2bfac2a8f8713e165e684e44c1d7e99960bae0eee52a93f8315c8cd8a2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0c38e8753a48b4620958e2f463318921ed1dfecec955cc5b0021952bfad3e5272380900aaa0d400ab4fe19028c4aea9665ccaa92005995e470ce98611e5ff3063656c7e7347dd0d3cac7473edcd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1531f310521055534ba465ca8e91bebe2caab37ef26ca0969ff2a1e2775dc91e0c459535336f42e40bd88b63ffb83decf68e0e7942e3812af83ab8a2724aeb3e13834ad44db916d5999722dbd314d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1cd3c64df2726c3d4590f89be6a9b2c81259cd059a56d9b1e100de3ceea5e19ab260c575aeade1389cd6a6cc89b5810ff111dae5f921c6bf3814aef7b6fe4c2655c218e0a8117c0f2955e3b68ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1180a170fbff657a1ee2ae769e15df5152f280baa916db54c3144f0aed41d8c429dc4afdf2243f957a50c39a8d7761a5c53510aaef32f82acaf85037c0ca36d9e6240827e1cd917e4494b83f93f42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97c04cedff03b13dc6078fe0ba54a8e96ae5326c3ef8bb64cf34a50806160d108a8594e59f2bc35f320b33e991d941dd917ea483c0068412a7aee05f59bd8c3823f8f180b6b97abb4d057a1d0ef4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11080491eead4064d9ede20c9ff1c0bb6402279e8bdbea4cb0e3dabcbc6907d6b0a6a5c0e9778b7725d4e05ad123b95434dce87b12ebaa0a887455cac6232bf97d7be9daea380ad534685800a3a43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc42c161158d8e0d5a796e1b4e854b0a63a1b4ef6be4133303eb6c1d3c4d9ac78f55bfd96ef7e8cd0855d03db4e444c0982c1f6e895555af3baaed45c76fdbf1db5e395926b94b624ce967c8572e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17aad465eaa8797a9dae6c45188954e2385e7dd1f1e6c3689e627f88e6d4b8603b4eef611bfbe257b857694b4c8054e4d5066c9828f70aeb05bb6334b781da81d8eb7ab7d0c04a738be923abd87af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h474aadf53364c7236eb5ff755961f55ea124a6af699e164cec82c8182b7d00184bd0bfa6fd8bdf676104cd167518f0c59b23bf3204e379f1233bebfb5e235182d3b6569c64b934179f06ae1e947d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2afaa351566966b256b45f9e63968c9d1357b97ac7cf352849f25ab883b9d2d2a1bb0dc00a92175b27a39855abc55283152b255ac11542f7a0e72792a3ca410baa61d9693cd038430851ccb751f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h576a610fdb08aed12a8e30a3b3cf170001215c6109e09f36a3c9f8daaa04d0098067871e8a0774726d1795ddce492a72e02efe0a660e803aca5db729067f46ae755fc06c7c944b03c7995d80ff47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h367ca0b95f489cf498bfd82d8fe7f4beaf2b13b0d6ef1e5e9abe718b191a057cead8758716efe905d3cad9f63dd4bd34960046de58bd9937bf217312fe209df58cd738edaf7edeed1fedf1ef2000;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1521c5484be44ed11b82b9214e9734ecde6f56dfe6eeca635d4dd2f28dd9068828ee6821170a5efae14c83fc0670137e1b47327d663ef52124e8d692014bae0fd8dc399e10ca2f3b3b5b8aef7e19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10eb1f0f56d07324cf4aae6ff83ace4de30338f33a150baa318a3a18cc42b0f26b4c397d8091bd00af3ac9bb636cf30a20197090b7a20ea9bcc9980a301f299cfadcdec271a8d74d424bbf9e5b6e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16846c2a707824cca2f7b65398fee0df0ecbc2deb94765c121c45c3e34349112e5d087bc8ca7d8ed14239356e9e8dc540c77d459b4d80f14d44963df76f6fc779bfa52081eb51304440caa1f913ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e19751e54eda64f05608fce29fe0ae8b3d69263fae96469aa321c3baac046835657fcd16cafeebb4d598475af144220947fee7828eab1737dd16e68aa9a1671e6a3b0e2b341ccd1baaa4e55fefb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a98f4bf067e2641515ccc3373657a541ac6e8974e702213b481297c8e172ee1de4e4fdd963702b1cc553f40f54b6cd20edce80c6aaa7b70565ebdd9e912ff88c15a74f646fb74ab472c2547437b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a285f8600aab7dfa1626c43f3b0b067bebc1a56b2cd7f15083cbccaafae5599442a9a5714b644a2045bc84cd8bf689708e387309e8f87e8a16a7fa87a6826ee73d31a3d5b18142af15a0d1470427;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2925ea04ae39b021fe004033daa4403cc206066d5289069fb791cd2789f769681cbb17a27299b6464beb98c19ed57b7a4f676f2b1ba10337076f170ba6df739126d0d64b014ad763dddd06e621d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h304baf0d4c21b5c847cb6254e388587297fe59631708795632c6a7921b093db9f693c8086cb04f87e2fd7a89a42cc6a590f37cc218e061778ae6576c3390a702c0188df471a66ef9176028233307;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5c3fb72b3a1ae4ca159ef81bb344757d84063a45d4e63a5a65a8610c01519588cfe97ecc0e6c682dc4a84a7091f76e19824d98c8cbcb9af8717537399ba314b6b2b9c577767d8cf9de4e9a05729;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181d3cde8cd89418d9cff974681dd393cede46c2bbd4c47b83cb93cd41c973f6eaceebae0e283d1c3ab56c17046ad3f26467b9209096d04579eae242ae30f0f3abafc2ab4694f8ff7014445a9229c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133529f0d500a33226b6eba8e702e6486a45b61a1222fda96a15344e749df7623e93d867ef681db04e2da34b568e8e37ed4013f1f8fc3d51cce0656f7965725981a32e5d7dea89098c62f450cc8fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141b470279127cfbaeab437be43ed17e12dae9b1dcf94e0e35d20a50928db7b394b7ed7267e7a9f485ccf6b03c5474c1cff6e9749983091d2dac3a2840560ce22a9d3e3b3c1d73c3ab4f49fa2031f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ac73e6e000d56da50d7b1697bb7e482e259f04cafaf399d0a3617e0c18a590a140a98fa4e32d8643e1b8593aa5a16eacacb9b6f1c16527da2441e76d6f3747e9e65409329be19ffe36918524d89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9e73f49c014514cf7a60c8b8cd9ad56421ef8701dcf9d11520d8a8172e75c40696b4de06150ab503cd4a55832b9bb63692171bd6afa3cf0f6011d765525a6aa043d5698be0ebb1657e98d8d5409;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb0e94310f931a3dc898bdd4ded8f483b4244148d5d3eba27b4b61bdc924769206df863f74014c6d6a6c3e23bcc919c693e61b2184d276e57fe40460e689b2777124f667cb6bc3ea674103c4649c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e25e0647b06ee92ff871498d10e26dc87f403e409ac977f2fe6bc630c27b983d4dd05aa3d296cd49058cf55e717669b4be597b5859282bb17e728d11df705f9655560c582dd5f8a2ad1ac7f84017;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f01e5e1c886239acf3dd4b206ee5534b4242c12519df2f306eff98d233d962dba59060ff4691f2cd83a8d3f055a147984f655446598330b1a984eb978151f8558208d68da8923f66ecba67e9df61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb4f839268d4abb26eadb49f8566c780d6696ae50fa300f7558fc7b27c863a41791dc31f0a3ec998c21cc01cd919daef55b013a4e4e2b39d1c37177a9ff9c19ce7606ebe990993ea56f67397c7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a30837c3086d6d6fafdfb73f5126f83d8f181f12d65b5be7f36ff6826ed87d09687f893cefc40e1f18d1e7f2420d6b19b7f1203170ab6e176dcbe55c48d8aa1ade3bddae23e60f65fc6e2b1c6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d85c7fdd0fc5fdbd45dbb756384452607872a167df351c86b5f5a689080bae9706f5d80b320f8e7bab5dea0d82ef96903077d973e3dc6a3849cc1ca4c881853abf4e1a35a0e9853a577566638f7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9d51ad63c0f4c9fe6fc6c5c94229190a4a6bb48dd91d85395045cffe18b5a2ec06a39a5489d76dd224f7c9538ecd26689afd7bd737af223467d78ceb151f218ff466969c323ba4d6ee8a7cc292;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad3299c97a00a2953605dc8cbc3b1559f43fd4f0a4807b20db66783876c116a2fca4d1ec7a16265f89f7cd4fae7f66ccdfdbcf4af6bff6bed936addd1e60022d04829ace21859fcb880373b1fb9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4aa7668d94b1a645e12dbe06ed37ab76abd00aae0a13ccde16eadf45e924cbb1b8f2d44123276481b086bc657a1f262a957626e249bcff7115f32cc969fa99054ca2080b43711ace52153db857fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26e502a8c6f1014f6c78c4a36afbb9cb72d5f4355b05c38e9fa4bd29d7d34aeb37773bde8200f475791837b5b338ad41d5605a522bddc64c48c3070c8873cf79e0c429029477b6312206a758b7c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dccd820f25ccccdd7a9f306b3b0e57f85c2df5dd7bc179a090405cdc8294a9c8b77125eb63e630c54a6e94d09b23786edd2c46ccc3b26dbf489b78adefc6a1ec4d62d6e62a86fb364818df70968;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h159ac02f394029f9cd46151d79f1da35ee0e64f7a51e84cff2741c5a1fdd90ab6bc417bde04cabb9b889cb1ebdcdcce565eac934386d735de23fc2c8a34b063ee2e8374640dc7075e59f678079b1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cac03a02949fb4a4e12c4847c0232c981ffb73559dd0e941315700cf8fa3bb4a1f04b8f36c6d63cede71ffa38ba7c9ab531fb8e7c77e12e6706e1c2d06d91b42354ccfe3fbe23775c39dff65960;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h619bfaa20ce393765d3f5846c36d2acd6a4bb5a0e9ab9fb334c33f98c21a364827dc3a651d6a39711f1f5d8bc89110896a93d77c8d049dd0ab35b62eed2b5c31f7fee03735445b65b083a38b4f5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h226eb9a292fbac9432cb0b6e01a3aa3bc9ede68de562dedd2372114b3783e37c828479477099b76bcc5b448a0031136ebb330672fe79ed0a242b9cc19e7afca622794d28ce4bfb08550a603f8436;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16788ea33844623202420fd2856e3ace10428ac53b0951843202b05b66e3062681a7cc12bb238817ded7ca80a601cb7e1256282453f986a280ba0178d850a9638d60a548f3bfe3a0922865aaa4222;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d08a5d9dbcfc85512015c74b02af7b2c383dcc53e1b850fe74c053de39b7c6f7509119e41dbb124737cec95394fa2f30fd73a0071de5157083d6f524ff10c103da9314362eb0467604237b51cff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc95c52230cf3afbe192f86764e3d8ee5d4d490a9d788359e4c17b9ef5ec31b478e859d32b769ff07250ab88523d71208bd7e22561ef74d9f4561ab8c67b59b97728def61c3fd9b8bab4e0a6122c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72cfc6519e84e3e5061ad4def06c08f8596829537649d5a5a2680da62963b4334fc839aaf6a3b878b2e692bb666b255a6836253fc32a00973c3c9350a20cc990dd9b473512adbe3a95bbb426cc8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ff492ac03a27a28621e2b14931876e1f6a1d8d8591de49578f70f0795a700bb592754549ac935372dec724f0f08172a4d34c246866291ad8d01c11b631fa149400f6bf1d441ce2dc6bf8b124c4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109865d285456273fe7d21d724ac22e2aa090b0eab38097036ba8e84ebe349e491338021cfd0e8dc5807851810d701cbde0f6c69a5e316082b510c3830c8f4d1c56ce7b2beb39da3a31b6af2a2bbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1161933cfcc608767380a6ab41fe323572e6955a29307cb0c87dd8e825d80020cae2b495384c8bd1ff3d31bbea62d0bc1e4298f3ee657f62d7d8d41a30016d2c7c853c5452a09939694283207263a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5e674d462691649c32ebf66b2928c0b56b09078c2f62d81320bf43af781eaf1477890ff0e6231d75ad2921e9309d912579ca2646dd71291b8ffd243c3bc62f82edbe7877e9f5cac9ba125d315cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2eaa7e966d448ab2244fa2a4d5627fd3e1f19c5d760ce9f5bf075ab2ad01deca1d1d887678bb31b86b1c1894f27e43d11fa06ec712027369d8685177beae3fd28ba09e4df41f830337343a608159;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf142c2b1b2758950234d0397072c173ece3868d04249baa86b2dc079c72f0e0e34c89c2c0f0da0079c1e312caaf3d2c4a30572da1dca54eeb27ab2b2915e1be0cedcbf2c80dad1810731ba024a5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17efdbb3c5b69a69d77ce2b20e8ad702e0ce49499fb17760e5c465ba8499eecba3fa96e776eef09492f9a5283e27b96373339edc8c6a9b969057f606530f2bf81077dfa12b6d0164d188d20f10dc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1268e042223e1bfee19a72a8a93f78fe391e7902179d362839f0c5347f3627173b48ca6103087df5d605f38b35e5ae9e530132086797f712b079588c3532200b44f0626ae429946a1e62e0c5294cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b0b1a405e4a451050afbd6d7bffc4ba54a392fe897f41eb5bff75e8d96bde990212c91d41f96ac2d0ca66e9c8548635a665eac34a960763e41ae34755f008e81f945aed59523e8d8d907d134f86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1545d59d7cae967007c6e8536692a306ad2107ae65381c078b990d1056f5e8bb132b957d4a68a72f962ccb7b245d3ac2ccc00789ba4f6f1f7d2c9dbc6ec61fabf3b5947e11268828b6522b7a0968f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197c6a5f504e45240ab8bd5aa30af7567bb1d99aaf473d2d8634e8b624a33c6a614fe8e49a51077d3bf5504b4a654c9ed4117df699357671f9dc24bfb06f9a652decac5d350dfb8d8caa52243dbfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h755916c4f285de71416bcd7d54161baa6378a9b09b6e1446b008f5ce15f8cb427df0b5a384f8d86aac2c99676c0c608d97d2a7e232c4b418766ddf211fba38a09b877685ecc457a494ddd3d090c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7984b84d60c75dd7eda562e9aa2a103bc2703b5326be09d79a0a6115da1dc2414d01e1ea9acf2272c9ea7abce0e0d938924e5da7716c7cee44de5c07a2255fdcdbb91c10bf39750f26955992596;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123f8ddfb528589aa58ee74fe44ef620e6630a85bb333e8a9025370aa992db7e0b1b0cb58097f324906028f99ef3e2d37034e069a590198ab8c76d2795338056faefcc09ade4ff2bc474ecf9f57f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h729b4be9948bf2f40dd7ac127a7492d846314133d7d25d7f5e9f639f7b2e4050c384869228c7cc667db5a1539fc977ffbe69482d0878d55ba674dd40d60b98d406311cc8470c1199d505900a506d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha98aa0ff3ed0a4575b1df694e0655f3102ccf40bbe7978ba0960ab3d7086ff314724bcf01084144e5a956e5a509f3392185be5b783c373aeb0fd7037323ea66d0ff4fb640236f35e521bcaf68f51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d446567fdc8d1f0a94b581fe64349ee121a144a16f8e0651deff7e2b9920b3b185343a3966389ba2ace6819b220d5d4cd43641789e2edd3d1ce12715e6a6e1c8a058d898c456f19e368cf0ef97ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6111cb8526cfd97b247057d7213f91acfd28ac97ad287050432623683030c6bff3d0743172e7be2d5dfc6bec62caf85434fb5c018f78fbcff9b71be27fc6dea445e210e201500f4b0fe6d3e5da13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15234c0d778e48b8830312ed0f8be73ba7bf5d2f201be05b071358f3f5aee79eaea17635e89f17fc5d73718fd324890d18cff9987e0e74852d1f013003e945a16c2798858038404448fadacfe04fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec28853abcc901a101fd3dcc006b83e72544518fe17740e6b0171fce19074158e6acbd96c5c4884dde15fb1f48f97e85baee06e36dc4cac8806d82ad6ae202a5b609b659991f551a5ad8eb74bbc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1d84766b0603fd95d7ac1de03cf10e2433b191c6af105ccdd10aa6474bb321aad8d9c355d2f2a4f331ae665d2e12a8f81b0a4d02a1f9827fee8ef33dc4c635b2533ad8841e7b1192f00cfc0aa5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30b1dfcf831ba81b8462f3c1fb2afd3d1508f1e6d93b97e68aeac155560c5625da9d4bfd3036a976636c2e82c646b2dc5cd196196e4d2e57570db164304da426f86a175f6b68f699cf6fafbc9b5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb564ca100f190d95f07f0410dccb726e8de51138bf02306c07f37f6f0ba38a9135ab9398733e67e532fd48997a1be6335b21a7f28fabbc6636b1d5d649a673ca38def75e03e5fd417c736cff00db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe9d882911d1550c18ee113132e24062b7aef76c789c224b2f1835d19a28f7e09457cf967f3373c91f620a7cfd30fd96a696cf665271d8782bf70c5f1e9154acecf7dbb18ca77b4a3c19c53834c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf95196b1d18a7ca09eeb3ede69c43a31c95afc021be64a6ba4b3a0d6d3b40f1d57781d09e1ff53dadb32fb8b7386446863e7edb486609366feabe15cab781e39f358bdaa88dabce65583aad8a6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9d95cb07d122de5cf2ad7ea8512bf36dcc0291a4027f7275c46ce64658d35423b19e8f7273212c224401e95404e1cfa3edd261d7fd38e2f63476eb45b1c567511c6baaeea8317324ae36e9ad7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e97387b261c2d95fa0e2586989171d5d80f68c0023621a766a250ae69d7332b440e84c65bb76a2d706905e9dbc099c1a125afae491fc394937e166e23a24254628ade0ecd15de34f9fdcdaf09b0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h334af4d6fe828dbe8bbfeccbb4049fa0cc463d99adfde3ba36b2a9f1799b1cb2a01ac961bacdc85f9f5aab04a3adb821a8e1da1ca7efe8d6b81ac3245542b70f81058aee81279d7f15082ae34b31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffaac17574537fcde97722e47d43758bac779d492e03cd70660cd5840508eb4f02148386ff2fdefbdcc626999c03037f0a7a134870ca3a0048c518c63cc69a7bb3b14dd563f7d9f412184fa4580e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31288e71cb3aaff174fbed4df376f83312cefba87c75a3a5d3c173ebb8d85e602b7781eef57dfb0df7c99f5ddfddd64d932e9dd983a929c8f572fa058297120bfb0187d1ff3d71b2de87183717b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6adc6dadfa20b92a2cc44c4ce4688443edee648e63d60260fc0b75171193cec0c98643834e92a60d6b7b48125af0292cbc3b7d59a86cfe0f0bf27012919bf589dd2b2f247acec7da9ae8df86e84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18343d8549df9f7517371722666b157a73b0e998a8b28872d35e32a422dcbf178e20576506c6d2bd0daef5757328ba3087748881ef9f5978cd469b272b1555ab5cd192100d04a5e2dc92b2a76a3dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5fd9b922973f36cd580ed7fe1c14d163d64ea904e281a9f276da9f26e0180e33d5e81d290c51a30b3e56c93007447906b2c39f88fe4086a56ad88053729b47781c523c7a33ae69a94ef0bf8b064;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h588006b54ac1c7438cdf52b2d1ed7c65822c2aa8704218ebdd959793be542b213b50b4636650e883fa2254bde33459998f249b6d97627c7605092524f97a076e0ec85cdaa74003c3b1c4f16b051f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f29be12adffa0550951740979b1e652c1f0f523f652d4b930d67b569ac4efeaeeeec99ca90a34d370474a2c1a10a70f20c0cf124293caaff71ff2c1e8bc0fc81e36f449da67a3da9c7260775725;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8f872d27c76a50fdf9284c23d35aa3b119f773ff815c8c13a825a02268b1a9bd52f0ba60c1610cc30696777c23818264eb62a83ab4a71ead7c56b9b78faa8d545c25c3c960849c062ff33448437;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4143ac4af5c4f17577be4ecbd50d90af502dcc38ccd89103c794c853738392dc8175e8848fc9c7a68839146102d55ea6f8f937fd78aba9b4b8f27d8fae9ec8fd4e1084ed9466cfd6b54b7daf999;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c756cd0151a91676fb9e6c1d4d600b1f00d8595ec140cc80c74c20c2988484343f9bcf81ce8a211c78ea289fc9b281b84df80e41fe046e706ed496585d1262814f07fcfcb07597a3ac7cb97fef6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4ab94c5365b2836dc1351ff31c8c9620efbfa155de3410c0f620dd1b277ba893c1efcbdd92272311f41e170ee894fcc507ce2bef64a24afa672a33f4dfd81d1a85b36f03651a2d29bfe69889774;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb88b46ed5726652a3560cb4005a29b9fd50e891ec4d3307954fc9f4c45cb6b6dd629ba4901ef395275a2b4b9ea1f399010466bca3cab8821b8c7df150212bfbfe72deb34c8cc612bfac7870c3768;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda5a69fe07baef8e46d163b8d19293041ff7ae1607cc9e0b6d2a56bf634ebb0125885b5bc7eaef9b856899d8880812b30eecb7014517c71fdf97714fa199c3503e7711f96631b48c4eace8818dc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d99d72f6204ef31f4c6e6d1e946ebc04e0e68a91b8318658a55e69758fbd037b7e82364c61da65c50e0448a6b507160b2be1e340145ab39c735c705ce9e5f6cc32c7cac60c94534c7d29c07911ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h755cc898395b15a8a8ce4b7acfe1f15565a4bbede375f3cb42b695509bf48962f8528addc6034ef624b9e414f69dcccd47de1c0fbbf7c8755423b5b96dcca023eb2f24428b3d0d1a30612e27e1da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd783b35bfb3b0f07eee5dfc2bed111238e5f5d3584801bfc5dc763820f68c5e8ed52c7ef2d9e446488741052867eb46f1c369cc0802a099411c49e65b04cecf3fc5647d07efe7f74398128760944;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf4a893fecf5dee9415fd5e84179cd92582117e839bb3faf877ce2db2fa54ec1e07d8d31f6412a786c7ea8cf08540bfee4c2336ab9668937ce03df3f9864958630c0a339113bcb56af3e16776d09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14cdaf7801ff8448fff11d491fd73387e3980e2b244f134f2736ea8827039a1ffeb803e540401aa843b68f1ba8c05c96f82986276c445f0f1518f9e7a1d17ca5a16bf26ca290184c47f72946a37a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15da3133859baed58e56e28f3c8bdb98f155ba2973dce277b5b764d84634cb381ff258b9755c8f4c21583b18e2c71d2426db6afa1a474efcfc3b08957d0a0c4263de7f9c8c8c3b64769e5e1ab339;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee6921afe9dc290673e1de6c9248fafcab9b81a548d7aea3e7ab36f1d5ab2574ea9cfa94effd6cdf43caae3bbca9537cf798c5bff50b1fc616841cc24bbbea0b52637959efcbf15f072e44485ec1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c37a6c49d9de8142ba8af267e0f243f2054e61bea13d6b83608defc1b5b27fa7b55a793a6a0183763348230309ed2d794817186cfd8d78c41f1fc18aec120e30ec25f9f13b1afeb3a9551ffa1a7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc2275b6c6d63121dda72ac2d7f246df6e07c4ee85a8361ddccea56bdf1df46ae3feaccdf0d33e8888fcf8cb960a1bf9a02e22a0614420c731606d611aabc0a1cfa75f7d787a1143073ca6bd5a8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f456e8af1e8969e57f6a421513b98500aace50226595a76f848092c34ac654b939d6e3958936a3c28ca1d56e95dd192ed4f69076fe39bc1513bfcf43d48aca8072f04e21638d7feae526b1e6bcca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15506964f79241541672cfdfb9b561f3684a12ba8103ee171d15cf2d0401324fe922631a70ea5aba0b78bacbeeb9e85d81994d27836c2c6b9064426ab778fb37c6e9b3220c5c8565c3adccc712c5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134d8735e225da884eb3353539f48569637fde103d0f249fc61e43534e26c8eedc2537775cb05cdb121e25fb5203a479d0740549942cbc5197315f4d3de8e2f9a2403615964ec16435c842a422d4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4d6f599b89378993b4d081ade9982b1ca7d1fd78c5146c058e47301ca804e6e10ebde3fbe9be3391f37a61a87be0970dab1958499eae124ad4d9393fe9e4ebead1e2967795887939e72a630d47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25b725bfd2e18e12783c4ef7f738b91975d83853dbd522a0303ff1da87a218397bddc137d7cbc3d29222ec2112234437d69c3a21809531431b9f482cac37209a14b922693ed63c3b0698fd5d794b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b71b4feb1bdaa741e38e2b64e48a620f8355efb7540ecb54b8ac47b281eb2297b7c6c25ffebba4058dd88ed394af4fe21eda572e24de93776b9fb2efec247e8d32fc367e3d9ebbf49cb9450385b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117344488bc0577519080e0b2db7834bcf47368c8b26ef543e2e7856cb8b0bbcef29b32cc1a7557f4a3adefe029a9b251e2e457dd8bba666546b9f57517b058cc3777e8cb80d9f079408fe53c6a0f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd653277f65342e6dd8932ec849f108c036753f0bb1c08a508a2165324aaeeb2bb39dce6a86852f8633408ed17e30f3c5ef0db0f4e4af3b2bebfa6f4092a11bd15c035775f5c97a3781750187e4b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103d5107cf28ae4e9d5d29c7dae606cee3b5cd48a9bc5bda314f6de2178e30d9608e57f7a1ea9704ba57bbd35dcc2fec264a8fe2e6328884f6b9c413e44b1df018a57f97188d8182f8c4ffb81f869;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25595c9844ea5207391e9db47c203481b8d23f3f62dfffa8f99dcb1f0624e3ad6fd85a785bf6866993b3c30cf70aa4c1f92f943911a391546d3e95d0d7e68e5d6a488f99507f0c050d25aa10220c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5cf1e027e1a0756447de79d9e1435f9facb0bbf03afc5f6139417a41ba897ff5d6e6f56faad0c495c7e5e3b00cd39f266321abfdc17e743c0de924f549fcd489c4a74f5481e75464ad283daff509;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7eaa530fe773355b07e798e4f5d6b9963a3cf00b22734d49210388d4ce818c0d7300d94899549d26fa988e78dc0c981f27b43ec812b427cf23217cd630a1e67d55dfe6b9b4d72b093a30be7f0a91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6043d9de47366df91996ca3a0d0512e9aa40c2876bad8d5f68fa31594b1c40456dd68c54059cf19f26aaa48952573a629332124cc58c1fc98b17345e3ede838b3839f21ec9e7400113197671e1f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf11a2fc3f13d9d015a8a1446fca0346589d7703264d06087ae8000e1a289fa5983aa7b1174da7b457e8a444f284c678f44396e8deedf57f29d1fd1fa2fa60e7e6a4cc1e212f8c0109e31b67d0f7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1963a1fb1d4b4d223975eea6dcf32119e754a5522ffcaed75e12ce16f0c932de0fc71685b28b495755c7a87ce7472cdd29d610d766274b3f9978e09a3986017506d6583cdcaf12a6714944a9fdec2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf1b82548cfcb556b2cb5b4aa795b7794a60fab30e9217134f4113bfbf5951ac100deae6e289c3bd1b567144eb197be6b58ffb048f20fa9a06e6978fcd489e2df394f47a3d5e1400bb1a20a7cb9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3ac3e6c92c1cb4356b6df5b50903828c2a21a424b4f66dc18e59926949132df29ddd6b48ce5b52e2627a5e06760f1bc9a5b36a50581377fa2fd8eec56aee07c2db889429335fec9cb4f2a7f1cc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a41e1dc67691d7df7feb1fc47c139c4b96734736f2d1d0bb70041a1a9a3f4e2020f132f62d3df8ba79464dd00ff1aacbdd7d0615d9ecdac8e77d0719d03d2d140b957519f1ca432ee4500128f737;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha877c0785baa08f920e880eb4d0f0cfe1cb6083781d0f1b682a1c122093dba44875fcbe971c07a9ec61851bc5b3e9b01d949699b68015c9189b9c9e9c6abcee4708af600b4ea9fc6ee0841a1b923;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c2fc7ae9388e4a48cbc781e02ff7569b0a956d6d63b61df469322e84d6bd0128f1c1b508f3ced8594878aee83d433b4e6e1c11f5b23f731edd4ca2c42b624448016e03622c4c921373b83be7973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1557f54b9d34450a32203a7e9cba5861e5fcb1659ec66e33b85f50b8970219695a990acd1dcb9fcf85f43991e18fa309286c6bfac1fbdf71e382e4a023967efae997e6ee52a39c69425613b503529;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha433ee733789ff2ae5875a54ffec3caddaf66478ef91a343681db769c7471727669f821df5cf9e803cc4fe117e3d1e9aad036b2ffd78cd6a3eee7f9dfd9a8f16435d9891b59520490980f80ec384;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181bc941f79e2327ec86f116c3eb006b78ba26b76efc1c4c9554f29e12ad2b90296ae32678081aec96fe4d6d54a8e499c818adaa0e39a76db0ebe9c24b5d58873c6e77e1296b3b9afef8dc9d80b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98d11aeb4d77ed86bf91b0f6ad4195bb63116cb20e4aef9aa976248d8d6db5f033d8d36bfcae16d54332ba7f47062d2ddbcdefdf0a135269aab0cc2234f9d4c0480f33bf89951d12ca1b129f583a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12af3f66d91d17b63661cd14fa18a43fc93fad2fa2acd9fcb5df5de7b4cdf47a8428d624a6cb3b220591a77f2a48f3ee3b3b87f65ef19bd2f7bdea01e17ef743d77da6c55d69088c6d5a0f05fe31b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h596161919cf80721b55cb8aba978b80a2b4451ac75289ceb238e8f9b6f80716d4c7de7afc644d7f04d19db39527b49cece2582a5baeb6301f6425cdb8a7edde87e571404f67dc56c20edb03f5433;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65bb6a57b32c83fb7de278be1f987eb02e5bad54e8ed1aab255dd04e7cc43dd9da3684f3b4a9cf4b5132f363d25197442b5205a0d7b27ac1a2c5adcbbe8e04287b94bc93212347e7087351f65837;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96684965ac0d0e45ff6b2b58e6c49d63d99413b664de9f1c66e357acd075ade1238b0eeb01ebe99f6b69f7b01cddb84fc6b3b52f397abdce3dfbcc64a9db7a38329702e2d3acacb1df4d323241f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1201ba083b575dd4bd6b5f2ae487404ff1b02d7f94d7f5f046a4a69495cc6933d5eb716d47ac4c12c2f2d5af726c21a9c2652216307d149119a382d97ea07f7446de084686183d7f9606805e233e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad82df385b9239a0c2452ca44e3ebe4cafbac4979680288f84dd37deb962a742617210a685b7d9081b448d9c038bf44a0e2586c93fe83d778aefe41fc08a1b85dd4e20776f5d596e7cd5345fbe9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105632cfd4ba6fdc2f7775a04bff25ca5dc9f5dc43e1cdd4a127fcedff94c629feebdfdf9171451257329213da91bc4cb7ddaf1b049b9f0455661e80d8dbddf030ae0d691aaa41fdfa66b0042da0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c28135b9fabc8cf0d367a39c91d07d23fd8d3ec8241012c6793efead213537be98794c836b8b49510b17d7934f98ec2fff96c48ce533ff41c602776b885f23a80b9fdb21ac24da0fc390fc4becec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14122979f7e967d392ac2f8cf53ada89e66e548b95a5a8617fa543a221141716221d4ac1812cdba210c932d4208d074d49c6657e9e040ad55d954c5f83a079d140db5f7c35df62eef3a2c404d24a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9657b05b9a881193eccb6980b9c7aaafaf2b639087fc65c7d842f84e3fea09a5cb6764633cba87dfc38b36c9c3d5aa1d4776dfaf38bd4e3e3f25d7394216ef52d03e85a9461b833a3ff517539900;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b078a3c65f8347d9be046d72eddf0be7ce47aa1062689180e23fbc198ae5cbcde05a73d6f1bde71b1326c69f03c3e45798cdf50868b41a270adb58648c17c1cbad540516c7c793f7201f578a970;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11fb042c33b78c1bd62cfaa3f7232702cf744f573a260eafdeb0da662421d2fd0af91efd4d1d8485c4bb5d9628b3a6217c7cf03f1abc6e5aae1e7f00217d975fef6789336340ce670ae865d917561;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2e7ad60e558eac737d319f357118f5147eada3339d58800d8543a648de291dfbb7fcfc75afba1a21f583dff7f62921181a9be12e9df4fddb0467fddc45083480df2281e418dab1a3f0b7fc4000f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19692ced22b9e1bce3313024e256ce7f049716c5966092eac8edefdbba94e2e45b4ff19b45abf43175e03f65ba438f6b2afd22bdf26ae0c2c6dfbafdd66cc0ad14919fd639377909e8b8b491d10fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12913ff0c28d8205ddc99d4946fdea5daba9bcc337eef1797d7159027f86061644f32679a59004d8c857ac9f7fc6b43c0bf67f2cb7dcba9342941a63d13ec3d8606e735a832a11ec7df3f9c471e5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11caa8c26dd34346c9a251e3d6a139300ff92989d2cec8b9a4a42ee7964e257c8cee0190285276733fcc878eba58a897e642d705bcb48785b3322131387d82d6be8bc9f30c51cb4543c58ad9b73d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf70e73ea74e9099a26e6c8f6969841d59f9d47d47620fdab308a41c95547168155b8c755e3e8e38e30e41dfa4392cdd769252ba8feb26a3d8692fb26d0f01c31267d76a8faeb99e9279cc7a519;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dc51da1bde214e1b421671af055c0b9e90c28de9b3d4b12c2bf6d8096b79ec5d94b8f3bb59833ae489fb5ec462c0030ea166da1d0f5b8a13cbc1b276371aa907601974181da12fdda949995522b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f03b20400a039121961b240d739409b761f73c9fc734280dab30493b8acce5f3a2d16facd23f1b70e5151e2f2a816b603ab7a093c700da96fe68ced8deeaff1bf0ebc2e161c9e8c79afe557f298;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e28e2374da106f8b3e42484b8dd24ad406013c58885d4afb6e81f6da5e359de1c43e3e68807b0584a39c1b7c426aa9972cdce66d33a931d5b25ccef1e7ef536e411d2fdb2139f12886f65286333a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1106e8b9ab31a2e3c1817222680a5cdfad982e3dadd872857c10733d95de278cc13e9aebaed9dab86c8b27b39a6802eb70cc6c8ebf06d457228a259e2c1698b2d993ee95bcfdfde9c8b0371acdbce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h301d39bb64281cd9c3f0a7b390b07ff20618ebd14a117296997921dfd640f371d163f66fd5be034d2336cad75d470388e02840c9103116dc9741c8853e7f80558614883b693cac8dab7f05a9cc4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142c21b4ebc3d993ff68d93a41ddf661b7ece6c01e5fbf51e45f92e858c3f8dc82424eac8161939ff2f7478f04b13e7ca2eba615570c14aba598f9ea940f65102c42940d4c8c32167b28b1375dfbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1e63b5a351338b8287b5132ed7bfc88d3625c901bdb2375e899bd19bce3b4c701afd50ddbeb964e52ac26bb5e0f53de524c54053c9abac5c05d41194461d6771a2cb43315359624707087564015;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f5f6c7630291b6a18292262be1db8becf1fe53e5cffa29926fd0af319aa6d98ce5ebb0aa2d4576bd3777879edde73ad4f8d1f7ccb5d163c2fe2264f78da0a67cb1963b9cc0c63c7507eb8704287;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130e9a0243314820a43951a4d6b4ddfb3744ed07205529cb7551aa49586db00171353cb2a4bdbfab54a437fead38629b9038d984c2bea2f48c7b6cd4fa198d8d4db0d6bd0fe63e4774a8545f54384;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a864cae74272d3d3e90802e7f3b9a7fa3ac53f29c1386d217e67b2f70ad49985839d38be188d32143e5ece1cf4d38116db2440df0189499b2ae07af7fed2241306699775596871c9621d3921cc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc8eaf531a26969cd83275f8aa689006264ee992b235f905bf9bdf007564e00121e5113e4bf493fd964d4efbd5f39f88af95774041fd914f9f319be80bb42e0afab9f1f3211b34588f67e7fe2cdc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ab7e65730ff4d2fa42bfd7fedc6dda6e3243db79be539ddc8d4b58701f567b4a71b158026a8fa7b937a830063e88425a91eaf906f1a809afd71d1857a0a68de4d31d3dc5941726d3e20a2527e1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1677559764b9b8b1d112352b4e22691a3b5abf16d6c545d75e06db88ffff5413fd14a368e86d69e636a66e0de14cd9cf64d68c040c1cc24b014c88cf9769a21a01d7c40f181ce51fb4483afcf48ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42d2c677695a928fa8b296ea5e65ba2da7ddc51c687cbc5f44a4975cb806c6cb14f2a31ac0a0aaffd88270077eab7a3328e5dd87842d8867f9183686cb196d13366083b3e44d481ae33c54314984;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a123a5192c3f3c794b58f6a3ad75b0b389796722f7f8c4574e0a26aa9b6a746dc1ee20c0f6ee46df97d6e6b615af6949b79c561098ea04fe43e3496006cf934dcce2f05fe9d00d91037fc5aae4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1169e85497811924978ca4c9b2601c331407493ff100803a66c1e1d165f3fb732f86fd646da2a3a3792aaac80cffe47848132a9e8e6d7d9bcc03f1cbc287452ffeade6b321b42f5736b55aa414666;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a904e4f2edfce0eb3416c0348514d6065b7be46b0af7a3130515d5e4f13295cab7897639b34d6b06bbb8e7d0326a8bd5bfc1142608652f7af52802b5eae77965fbc829160618c3623fc6da38f322;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61bc9a561f2cd2975903fcb474a7de749d836c833c508331cbc7bc285211e1a0ba851f725d76c2c88e642ba9876a6c34771f63e0cfe707212c82dfa5ad28d26dd2c55f6f593e3c77c4bac030c24c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ef1301b84dd9610cc902edc80ea34c40cf314a0cb8b88279cf863d4eed5901337458435c80f3355d67f3dc93632bc0a1bc764267760fd59ed6b96041ca7ca417e468e74f5fdfc6a4033d7c0de6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff62626ac513c9c30b36404995b8cf2b0e51eaecc9915a2ed4db24c0d1eaf48cb7915c12195ac4e2613a43ed803e3e8cf9acc8c78b655e7b0d1812fc3057342565a9f8d11966bcc46ba8306caf81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9dc5457a7583648f2a770c741fd2f065a906ba8a730fc870d6dfa081c4c9e59d52e28f1eef71e63836aebd9457efc7a4ca106fee52017be499c13be5764d12b64947e74dbf355a11cfbbb29eb5c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1452b4519c3d30750055c33488a22d169ead2a68afa14b7570ab332888cb11482f23af95b53c98a755e583f963df9d74e7a6040e2cb8e1779d9be3604f1ce05452d83d96afcbeb4d906c18b8deb24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4e739d746e10107e1028cea1e142de6d764680b2df5d2ce628e650c7fb3dfdc004215e3d52547a2c48d4fa2f1d7e6145abbc582d49f89f3d1e6069adeb0d2ad0734a3074cd8234eaf5ff9af4603;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e621e5a6fb6e9ef7143fb58c586222847376ed3f057eed5de994e585fbb3b6571fc414b6b7056b4b8a9503340f109faafefea76393c5519eb0e0e18014df7276ed63cf0ab199138f00e5c13c376;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c17e4f7fd331e0cc55451e6dcb569aea803e15cc393d14793335c3803791cfcb16efad2184c3b207e2e8959b8d6e6bf751978bab726bb7e9c5ff51b538f4cde91ffede17223aeb3a3367e23d332b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8d6f8c68dcb1b739ba58a141a88135e2a0579ed91a16d2d7d396741d616fd1e1851f65ae4ecf84848b3be5924440652acefc575d7e4d30231294cf4abb5cb43f688d77a7c07eee0e3b522501d4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb378af736788d628ba78e13d03ecb8ad82f78b3356f38c2df886aaf7d640b6251ee055012aab4e6e9560457b0efc7ed149e5a4ecb01cd1fde0fe01a945827e7743b2f05ee90b697bc2e70d4a5d44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddf26426ba819498712e993b766160fce5b66cb92a42112d2dd954e28c55a5467c2649d361f104364cf432b1e8d9d53bcb3e0b0c9ccda08a9b632d0f2c9e9374dcf755c44967866db965532a6e25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h269c703cc0d232e5030cffec8a30b1b16d571c975eca7d87a3f32f7f1d055d244b3dcd6a70914c80e3082731c0a8be855b49146899011eeb9588d93daffd8921e4577e425b9b0d93ebbc93050092;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddc557acd72ad88a3d98014e01091f8b4e26c26b0e982b10a6279d075648f80f8abcf2f31451d8901f77311804248b89b573b7bff27b7e1b31fef87950b307c96cf4f7421000eed8f898519a2991;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce36e7bf6ec35dc86658f751686b13be7e7f974a992e2af29348bd48971b2784384d1fb3593905073fb2ccf5a273e0451bd874662be4d5a35eddc2160fefcc896b0967503ec4f25395ccb4fe094e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he687048aa81fcc6cc32150cea60e2ddef2d58804e6326479d910db5e84850024d37fb9e75a45fe5dc4dd2eb4152be025343302beea7fc3993cc0c0eccc73a66db0d0f7ab9549d179b891dcd4fcef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165f00d071e203fef1ec2b33322160cf32fac41cc468ac29597a3430b652376af16bf73a7865f3ea524b4f271bb6c7c05583fe43a8fa03cb4d0c1339dcd58dc052eaae23c4ad7833896d6405979c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105d751d6b4b98401b13c95c6453aed30cc64bfa2901465b87917741d67356ef94b25c26164c505e0ffa94b4493fe6beb03b2ebc2ac73d5820af518f909497b6f21d0067d9baf7c123c49101f8c9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9a9453846acf494b7917f6e93216a7ea5a969e3f3b7758d4b58777b8e81ad210eea1435a68223d15a7b0fdf75e7be55060ea06e3324f19bb48d8cf5db329a97dfc8bb565e5e4412b98af120657e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8507c590c8de1de107b1d43feb7c6df325b1cd60d3615845621ea87ee0138476265e4fe5252d91ffc63d82d80792a1aeab482710dbc60c40b7bf2879b502ad58d78e056bebad2e4ef1289fca6290;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h738a740a606ccff4e3e99c13d484ee83f12a93858ca0f671f5a46f602445c2cb7599d1119b970d962fddfe8c9c2b55985a9ce81bc4db803bdfafbc33b28def0a8d4871365504ec6cdae8270a95b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8530d5b2b0e0a005deafd4c322baf0f16a6bb922bf907d462431866c49b3aa27608d3db609683857b31f219f9a09fc6d4741d1261aa82ce7d03b16c4fd360c5e5a3fddbd326c30a0aa8a271897a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ca71acd62cff4b77e80cb81fb104b8d9c6070031280ffe1b3cf92c609c9c63fcb0be01d41db4813cf1ac9cf58d9e2d92fad28b523eb094e6460af4340c987c6d9923ad13e3fb51f2fbd8d69d174;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf811593fb074a956182ce02269603b38cccbf8a1716bfc1999b8cd01ea8c50343f5a3627cdb64244a0f4ee3b4277c3e8116eec47a93455912d2b015e6d6dc21cfe33a709526d489b80450e7f270f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178faf594610ae0f4a28ca2792a10848e026e0cece3afe17e019d9b378a4663dbc8e67cb34c05dbcf3e84b3846d21113af2363444c676cb41806086a5fa1eec88796d9ea643927423d085ec8d0c84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17057893fc662ef2e4f89886db9968434e517e0338f920365c0a75b24289293a1a9ecda34553d1bf11c112d3fcebdc8a178f7451089f7dfca0691e42696ce642683c48e79069fc4764e5acb144cea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d36792c4d5be0991e5d5a425153fcd412b6327f92b6b2f4a6305397bff380f0b040a9a3247dff60855fd5a6831b3fd031cf3f9558281364e7595793b3a3e1810d739050d9ceb6a87460c3d97f40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15990b3cc1957c3c35d23e2dfdefedb6341aab07f7fbd68f911eaae17d3c24c49210902255b8b6a8ddd235deb19052da5666689f3f44bf33a0ee30c8f08d3f776bc251656123834bc3290841bd0fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d86b00773cff16f9843f95abad7147fa3eab9582577c0c69d96e9263d18054d0854bcf36ab4111ac95f5aa5605b3094c3e1c1e65b771b58f3b6fc6f0364d237eee4998c93d15ec34bfada200d31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9baaded98f63e9840a16508368ddd3ef7feeac846153c65c3d885ce9561a2cc7f2b5cb3751bd5fc06dd907fe10ce2da0c029ad5b6231419e5059ce60c8d90c8bb77dc671bf735d94701617a442c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15dc77ae8d56bea3c4636d18dc85dfaab8a73924fec89bcf6ab449b61aea239235fbfa9b649d8aa599d61b0e5fdd6b03017ab0169d7b420d2aa074500dbd10ffe3faa915221b7186e6ec299974834;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha316ef1330d96ba87d6fb4d63aa15c1d329619eec92701aed849af66b6b97e6e553a873c314c70281de8c4daae8680a024fd5f625146222ea2b0120206ae2f1bb479a6eead4b7543df728065e0b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbd447587ab9a006d3e54032268f64d8540c5c01403b9c9d27dd04f33058c12c289a64a8e5b8e0ae07ec3a13a208761eec776d5c0389e1658f2cbf9efa62a0f003c5aff494178caf7191912daf88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe96d7a267f4cfe5813b63a147b8564daf43527e7b11905c1053e09ad171f23c6d9eaee35adb4a9376b107df712b0988e91bccf3be378725514e37d8a056b7cd285db7754603edc123d132c7d286;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55e218f26153d0a5befc95e91ae3c9d21f5112bfbea5cc868d4d6257c6ae94460ee771e3008a42d74423e915f037469d2b05704d6900b72fdc072267f05c05079cfada1ad44328b2093f7b0c4d6a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h933ce62b5e950e70f6ef7885d4cc6c1c7819b457c3e87fba0a8ec27f31bc53b58942464073412072b07807914e937c13d8befcf208b544001dd4c72ad043640cb8045c428c81b713dfcdb2f950bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e9cf0307f33c40df5f6be49a6f7480089531ba4e10c92483a924abbcedb029a82ab49cec16b317becde530563c15a2f7c5f2d6e82185b37ac7c910aa09604110c5ee0a3155822590d2798853e31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6d7a2d8169ff8c545f7f08641a7ae3348b20f364c68ac34930b710a69a3959e2d2172572f5176915008702b5bbfa11000df70578795d0071e8c61855e0230803a068a0a5394ac8bf590bf78563b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1346542466d6601f92e911aae163bd0aebb1b2757b300a70bfe9b83d48dba0f58bcaafa2645a62fe1139bdc0025d3aeab4fa9aa2acf891cbffe6c94180035eaa9cac8ec28956a5cd524bdd27b6b1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2202e49209febe2d96bb0849965aebc5690dbcb90f4c38f704a72bc04d670053e0c76fc6e8004c7042cc1c86990dc71c5654257860ccde7c3c94d0b1ec188b74c80d7ca473c5935c1cfc109f49a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127a29a31e6e8cae9ec77abdf2a90a368819fed0a03afd407386df898ecc649bb7325cb91964ee50d4b047938fc228119dbdd38d00a72c36d878b10bed0042b97ac481b45dc3c879abf8fe281b50f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ca222653fded53b30f4afc3fb6f631f2dae8c7dcf1589baa2be492f31973d0add374b831ef1eb8b5a8108b27697005ff2e59ae9a1fefc399fe576ea101ed1bbbdc646d90a9d3577294db580a341;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26e99d884a5d2c73ee1554bbfce6dd9d3d653f84414eb97c893502c57f506c83b00f3b106f8672bf5be9620407e36c6d5805c1f63238d1adc3ce60c235d21db4a323c00d78ae225b859c8860031c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131c0426c732d647cb5a0f166d9fb909f9c85a2e24242df6414599c8e8a89e697bbf4efc7a2fa3cff90b53357fc2f66e33a6fed6f7ec49fc0192e19eecb698f0dbe604ddc3b4e1fa990440130a7b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hba83aec1290ccdfdf3c747497fdc063479a8bc20033a6c6c2966b9663622b3ce4ea16e865f1cefe24ce04ae3d8c9f3f4ba8a46f6be35446f7a002958607b9a82ae04960b90aa8c5bcad22e28a34b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf76fb9a78894311c5ccc87c0ba981c47fa1bc3fb8c38efac622f1af10fc1977298d73275a03f3c29ab22ecd60e7f2743a9ba18e441ac4da268e8a5b9460c419c57e8aab1c49eb955ed025b3cb373;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faa10de45929bd0331702267134608768f6787483872df2adb4f65935a5134718228827f48484a49332ff4f62aede711aca3788adfbecd937abe78e530c7cff3f5e6891e98398209ca7c3cb4db99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h644102741869ce6a50a34a0f0c387d1cabd9af3ea730b6cc68a2fd1275ed6ee71690515085155316d129bb5919ee48ee82fac5e69a6d2a8cebaad95aed9f347a1fc9184ee21a2984eabf9f90f205;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7582fbdb7f363bda7e32961c31d3eba9f3a1807f7afb3e6dd585c53fcc295cb8bed544459998a97ccb6ffd187a20f834d82b0dd0e8def93f36eb9d9bddc87d7802df0e2083ff3d9e5af2108f85c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12781644a94779ae0fde7801b3103166e99aa8f2791290a0b746f2cdb786957715550ce909f86301b609b8bd0e1cf4dd98d263d2daf049bcd81d77519dbc2123644db420f9cd123c5ae8c8578a4ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157f258a8ad885a37a08c4ecee6be84fec5cef6287fb667cb4480a0f4caa709dc1d2f8ed23fe08bab750bbafe0b16d394610c6a5a93165627713e96cdccb7be128dc4f15e3aeb948fb204f016cb1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a675ac946267998db23f411d2bded5a4277666bdc0cde2a493f58ad34e48ae2d7fbe95329c6c6624f3dbabf439c3ac515fbd984fc419f26c8ec2b4883d0b91ff56e1be490f774c36e637d22d0b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af395d02890db139d3288d04dc9354debdf60d6f45c69c6460739904828cf7f8b9492afb47def225f1284364b8523b35e8b41c711ed8f9bc20d273f7739bdde9b76a80eb6985b630bd2b9a7fa80d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed921e93e251275a0947bc40f85af3cfe1dea421c63dd6ae2019ba83a20be968f2c8365cb77964e5a87de49833dc732e125aebed9419582c08ab40d2676304613e00f42142e20946154b1170968a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f49c3091d59a998aba42992cad964da6839344f60a051a7dd489038f9d0477d371b2751a5e15cf5d1068779ea5555fc90626b26a0f50873d38ab64dc26869f9573ad7016fdb0f16531f4b9df1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha32f50e7ebbcfba3cabb8305af067ef8952f81a341d5be4aa5faa33f07f0d67191f60342e081f17d00f4544a52b10136abf5cafadf3f62143ee027ef4f330f69d016900c86d90f71fb649972b02d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ec1fd602c8b470bba2a556cd1d27b90eda3475dea886e16ef956f335b26d00073bc3b228be2593f80589eb255896e888d59dc82a42fe6eb49b380e47aece1e3c8417122f68e83c00c0b53e67aba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha329d1ccdb80506bd831b0bc7131322dad1bba166e40ae5d8d8b0b7f3bc23b608fea6e5fd5930fe8c3ac7c8ad2e4503e748906aaa26b34fb746d5397b8cef98f75382ecd792a1887954efbb1a841;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb26ab991a6a4fbb0a50e9a8364d5b5a5242aca877f8fd281675726323829ae204111b2009074a48a8c17b3f4048200cf54473483fb9d652154269aeb953d2ac8f97cf3a6d569e3ff0395f97185b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9184679c2ada5ce45251fbe25bb2716090b39ac7de61ba20962ec42e9c376965115a223c7bf692fe2ba77850c1668aa90271d6534f14f38c3286d80ba841634b86387b4b9e251131bb4b37d37128;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18659da6074968d56464c9645bba90011bd4bed0357b390e30fa1e9749ee8dbaf23796763dcb9028ce3408001560e96bc1f466e4c40d34760cbb0608edf245526c7fafd9d1bbb64346e036df3b9b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161d9bdd74b86144da339f5f6424fcbcef25ab19bceb4a5042d89bdce37557580ccd45ed65515cb9da9e5e556bd17ad7f003bf78dac655b520130d0b629db81040e664834c8ad980fc9d6095842d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191aa478fb8ba4e9a2bd48bd93bdfbff3284b3edc0a9912f06ae21054bceef8d5d6ad88bae153c1c175aa335acfba643f052fc1cdbd543e0134fcc92639fdbfbf95a961b6912843f5a6b75234bbe3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13010adf55e9ed55727e58d6a92cc4f17e056d6567532f824e4c4f5c13e2f18f86ee8928c7e9a1210445b698f76aa93b8904ad8e31d9d3e0ff1450511ddb2de7e08a1452121d19e8657e73ecf8bb3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ab43f56e06f43842100293f6201a7f497ce0e16b0cf6c46a71878cfcfb5144ff4165c70f5b91898f254d4678a13f894546ef2180abd3169713ddb5aaa56ca35fefa51d510c7e045248fd32cc948;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3c954b00412783ddcef0c6fae48808be6c3e1be922e0793dacf031a0674cfccd2584225e859981c76779916492ff0493f78760081eb426e0dadf8f36d213d4bdf348755398b46d192a48a7f59ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e69754cc73894ba43ff8946548acd23a5938732ac2dba46c65c1f42e8014d7bb6cd322b987ca705bbc1a965870941a98fb7c07fc9b21eccb393735bcb2c596eee17eaece3ef5c999fe6d85a4053;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b7f2a7776f9d7e8cb88a9770630471ae1212a26f4036a13613619e66b5a9b4279570c25320b158f0116c9e6462461d2f6c0f232adf2abd21390b23181e569b152d1f89ebbedd6678d5812beff03;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f3454967380f6424b0989211b7cd4fe7d1297e68fdb6138021035777cfe303a1ca53ccefa3c2a4ce49d925f84998f42745d5263a9a86da5428256eb5d6c2372ec1f9c196fb574ac7790e3ac8e82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e6a57a94603e4bbd64d1bfab11d396c98fa9fdf607b9f23b1c5d16cfc978666a5f0fe4df761c99e4aab651b10977369063607d732a143cd5a5e476cc0ebf1097c7d5e41be128492294d7a8cd74d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53a78bf2985d462f5af5fb53b93059eac2a15325674a577f9b4be8a128704961052a652dba14170280aad921044dfeb0b925cf471747668b2f35903fd11419cf05a49deddcee6dd22b0b0ecc43e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cafe72be48ed7e8adf585677e4a3884f3fb8b897b6377a241a35389c1df2cda1e32edc5f36aef3dab5b4d95245c8d7b636a2529ec1fb09701b249528a96b8bd7d2b646138e75033e2789788ae1bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1955513064c96a0464e6f2365249d16ddcb8bab20b6079cde06e0408eaa7a19bfc407550f930a4a51fdb4f174c2ae3cfb1b03e1d56b881ea69f3099980c19aa0af7eece183760ee2cf6a7bd36e03e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33576b17a9f12d1a694cbc20cc68a80a5eb42b2c9c2194e208ed7da25eb590c14ed06ee51d9e4c6631ffbcf58b7d0ed336ad23cef76e118b178be641258a3b928ad8e9578020aec22aa37af96e9b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f62d51233106e7aece6aba2fdcabb72d53970a6cdaf228379dc01ae4befab97121b0c48902d4945f5fa07a7727578334038716fdd9d05e95407e495d0ea708417cacfc873de35b30e0300ebc7a5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd1bc504fcc0c690998dc4fba13854b1f89e78f8d224ac1a9c2378507c7d7fa492240d7ab0202b36bf704e51e16b7fe191bb6447b4e3e37081978b6a5061d66b2a058cdb84db7958343ed94d0e2a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103e9d8fbd3d66effe26ff80a458921a42d3f2022cbb4724bc9c4b2dbc6f9d2eaf2e92c688faf6f9cb3c5c7be24a6dcbd0014a6c4dc71675b17362c6f18bc65f0e25e6386a4bb7bad3ca9722fab21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9f685fd39d46652465a67a1628374bbfbc2e186aed56adc3830a984e3a7a554650436e5927268df18a03386f1ff8de705fdbc0a579073a88cf5a2c38e9d138db7aa39141859056f6dee0d638ec9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f3dbb290aed705827f1b4ef504276e23fb6b40fca09988990040b1ff12c271a7951bcbabd1ed7c75c1ef16a316267a9ab3f74ccf794daab98cb04128f4f196ef102655f78b4b19f521f8746ac1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62097bcc73fcd8e7cf80ec86058d325c78375847392c7cc4d63cbeb09e04c2c1a0488ce12e2955246c0f05a6b97180073878374cb2a56ccedc313ca6e4cccb827d817e0fa24f5afe47b1300a6b74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c86e596810b3585a974a33f4c1c4d3fefee325a5e1220ef49a29c0652171b0110e8940886c84928a9cd2d21fa8fd419bf76fd39e43989baa5aa68d0e38bd9ded9ed05b2041b12ea30e903ddcf306;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b273691bf15e6171ad3e07aa584725320cde166cb802e36deb221a607fa9889bd3a6a75a89348876ce91e2083869c182d89e4d58441e063bfe8fc6fb3556c71d19686cf21006e48d2d1675f4f31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1517e524ffe52570e832dfbd1976e3e207bd5ea6185def2bce966eb98cc40f31a05ee3e8db90fb7dbd97ec4074f8e1fcb316abd8f8212716d576ae535be1b07519117e3a75d197d37eb899b5c56d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c0025378e05421ea8b0492c8bcb9e1a9a117d3b74f07f427990cb80ce412af10e1d1da71b6d934e2b44d70fdb9b7098fc403186180220855c84a9b127b5402224c6afeecb62a7159c724efe6ff0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h236eb1a6c95e764cd05680485be34ba0aeb700037336beb5ce0f8e024e535c0e862b5e5404567e2c804b118d0ae1f273fedbc42d8fd11ac6fbcffcb204aca5f1cfc103804d9477af77f3d33cd890;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9fd95af38f8b697f6bf4fcebb6650f4ab3d88811ac8b5399011960e843fa513571f2e5dd1bc94143153f4f9764de6e486f57ee87e51dbd05963f5df8606cef65b0dd4002ca19b065248875b1c20;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2984dea507d3b64e1464ccba01c47f4b0ab17ed0fe1525bb2a57e3eeef89536adcda2fe5dfa5050863f8f77cbe26f5209900ded3863aa8d519ad3e55971fe8544a57098836da63ad71123d9ace1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a73df63b7194c3ed985e5d07245f7fbf41072bb821c07d763f9682707c35f17fb4943d958976eed8d778f312c437cf377fc1f9794290a74d1242ec41493b07facf2330b7ec40494c8ee763422f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179ddc640974f2e984b5f77ec8724c70281cb8341bd2257aa98ceb8bf6b830b06df85cb3610ac5b9702f4082229e3f542efe0fcda41d50411687e0eb026f79c482c7387b9a472db35bc0238c390a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19edfed039e3a90c2f9a62f2bb96b9d174b30287a59b592fc284c406a47a6e4667de2bfb6872ca7a1c56d19fcd9782dacab2dc17625be13c9ac6c0b390a054b43f0be472ab33e16c15d0b4c392b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137f3760c6e59dac3e7dae4bd5605242b8a0ab56f27eb1fd89dd3cd1f3006eb1e2763503c44bf82a9f8e4e1ee4902bd1c8dde818072fa4aeb8493aee39d76f58776c439392d3da97d8a06bd7ca812;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49b508de846f09a69c7526b2e4e12ed795ce395fb90a6e7d3d3ad4a8477477bafb08e12991b4b02dba1db6d90f5fe2cb547e08762bd599174d604fbf7db18072cdaaa3b03a18c95b824724fad31c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191e2880a187c8daa3c083aadc44ea2024a99d621871b13125d30f4759b01b1cb648ccea91c317697d3c041ca2f5f975147d6f2425984758cd3585fa4f40719bc9544096eb842fe2f22bfb21e4af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h412d0f650dc2b91fcad3f31a8bbab8203e6280a810c908d10ffe42d9638ecfe0c1114e9987a0948b5f7d0a80860bec6ac8f715f5b505c7e4bf36d43e449f84efe8828a66f0b22f461f97f8b90183;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e74553210c42abc9bb9619bac0ec2f7d81012c32e437262332739809a24f048b6ee5fd91f82f2184f16e33da69497630f4fe8882c6a71870804c9f7ff345d564d6bf52f6df16353b68ceb58cde01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3d578e04fa47076f4cab1ae67141e13000dad188008e874ff771fba06f1a5ee7e312310613e8a46db16b12b55127cd95b073ba193ff6cbdc6a1bf170120daa7d5cf7f941c7770d0941e13b26a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77dc81264afeb76c7577b1d7025d010483c280aa3d1e919e4716e257d0547cce4db607756b978c1a9448f1a6a226784d0ddcbcb3947c06fb5f56176de99a9d283ef9767172144922aedba3b5babb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d53475e6c7d578c81b65f5b331b434b645638353c92aaa76fe0fc9f3c7fb0959d1f147d0837dea487ec0eac599dc60cc6b1a365e6eada9ced449d9f9cac0b8f6a238f8f29540db3f2720502e95f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ab5cc75417729e97d5a46c99a1907ed7a97a565d1588cd1edd22ea0149ededa185cf3848d2838f68c9ce4722d6a5007e94f982638cbe69ef8223ba5ad5d8e8ceddf9083845fb2b022a7c4554d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb533c0e839a67e6608ec58bde4ce715cd3c2354872de7bfb62730152dcd328d49a1b686bc9404fc9be6b75838d355b6739b2780a9491b97de49935f152dfd18cf2ea2fc0e47380e9f2dd2c565b8e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafe0bb620616ccca291781cd60880b9a01d745fa634e2e359cea418944e9c7592b8840b666d8b6175556cf613b0fa54e80d53138b4200268b08c8f57ac0838ca1e52d7c881513af90df3f368b0b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90f6f39e4d272df1500fa6ef320a24e345144934c19125547a2313adfab95d33493f78b6fa533800c703762e6dd4fada54b55e1418c8bbf9562162ac2affdfc9401870a4680377584858866dcf6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fdd26cda7094407b85de24f23b905a1b3c980435ccf8dbefdc09ddbe33e7632aa778fde4591fb14890edf2cb4de31cc90dd9cbdf3042093f34a70577ebd2d1a135c54917c429f0bf0e414a351fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd531b5b8fcd6bccfbae266038ddcfc1d18d03339e3f2f9c3c124e0aa601e37ab093ae093b1ebe8557c5f95e6bba86a8a73386a55bafe861a766b7c52a3301b4c2b3dc3b8653be3f07e156918636d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c78ebe3a122cb80a9a68bb20598a37e283329ec8e232e0964e8fafbd9a28799dd9b839a18db94657d9a70c20ec9bf6c5de0e7d7d0092e29e8920bcaa4d47b91e050723a56ea3b74345e1a5ed6587;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e659ea98038ad5e4670528202ebc89a87c22c0556ba21e4db36f2fbb9d87c8163c3ab827c58317e9f92f0204bef6ccc8831e346a5a97553f0ad97ae7a87b6633d2e2e2ff6b97dc02efafd5c83a0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d55fabb6c15adf065ff77b29ed0146688fb0319c136f0dd7fea079e5b5e5adeb7cfbf8396b5f7c79d70569be006b9224a0212be839d33932030007331cb598d6f786c485c7d004e70ac4b7a7bb62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149c5a0ef4728d16dff87eeb4996b2cc28bd094ff64239c1d776045ca89c07fbbb28471b35f79d5d7807e72e0949006216801c2d280b537c944026d7ba441826009cf06d0e90b163bfa3014303911;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h934676168134109e5400513d0d45558d6aa8714323e9a3f598343ef5018fc41d10c4d9b557cafddeda7dcc77f3bd80e8fba03c160eced666d7e9e569dd2d6e96f53a59e80454621fe63df65d7c7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38411edc619241181b15a6ad564543249cc50aa257fd552d33a028d09f8420d94e1726109f3cb1f184886d0cfa1a14937acbb0d8a3f540234834f0329c1c29361759cbd09107bf88d3ffc0adf9e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16cfcd9e3d401575e8d5b9d3ffb09b18ae5dee9eceaae444248f10d3faf8f6025d0328de7f549ef3d2e06dbc0dca078969c14a8b74e3aef19c76b726d8ec30bbdb782cdd4c3efd94aafea9256d9c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d19adaf1ec745f880fc3b632cfc216db803e18719decc99d332afa655915ff31a08da51d8fb0d512427815d786679893bf3b9d16ae9f66ab4a01db712b3e1a21b284e061007652a700f31cc3e22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a965b88699041d9b0e9d52170e8d79a57e04ec56a8ec9a6254585f13e68ec3d773ce0372b121c561afb7b15e311ef46f25a3f8a2bbc7905641f03337094b8bea78781fe60927399fed48ceafc89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea30d8216088a774ea5f79a54ec3480fec270365793aed00adccdade31dcf4135e9ab60ef15e81ed8a6b23a7412900ac858944b81d8e5936add792a52d05ed6e02a10cfbbc85f3e70277e67115e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb74ab3afe3c38d09103d265fe7cc2bce28f650e95a2d70cf53efef91ef2a28c05900d0ddbef0a5f77935c2e4c7ff6eadfbf6692d99fcd36e9ab80dd4d84d0a6de476df815bdf62dff8bc279cada;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9629617e32d1bcc824c7f60597f4d7906629dd0a31c17330f660829981235b4a8da8d32220ac5f2362f9711278bde75e2a84594249d8787eb10070f52ea8e9bef4df79b3bf4290cd9d77f8c924d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ff4cab78b31c0b13cfd90dcb3d8c5f4791b6bf21206513d2bad929486e899e87759ef922bac20c5ead922c053599470081a14be74b2e764644c2fc006a75d446cce5ac0828a476a2f94f7408cf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7968607eb3fe0022b790bf33ddbe76a1472a0fe1b29586c2c60fc9c9427cd197070dc8245adc8c0010c7e2cc4f6f2735178a0fdc8058acbd9b742468d46975fa9382518cac7c88d452fb642a58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea76f39c72c7f4810560610d3bd9ecfd81f46bdf72f2d9942da174fdf3caf999f9e28c61eda8c93cf6d03352cdde8b6791d9766ab54a81efc186237df36ac7331016be563837307eedcd51834471;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h301d1e94d9b2e138112f2ceebfc933d46e567c0601712e9afe06ac0ace2095b9ec91e430e94bcc9f0f2d2b2dc8a5592829e04fca8b3f09a50550cf35e908108d39b5b446b88b0637b687280ecd09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102409412842a6a1ba7e058bcc7baf505e6632a94eca240dc72f0878bbd3a44d8a3a5a19e6136c3c9757e77387395770610a25a1b01117beca366f5d04194c26a501a9333c0d2a8e7aa82d50ac7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ab09bf457dfda69937efae001ea8acd93bc1bbc4846aecb515d20a1afaa5a136f4b72e9b5aaaed2a51cc6f1aafd877d407c7eb76781ac1d5b3b19b1aaaf022934d76021ff0c383747de5f383f6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1800651653ec670ac39c31ab0f703a1755cc97fb4871ce8d3519f7b795df723f59b60d0ddbdaf91c456eff006ee720e2fca354f67ad278f3539f468095bc2239ad13edb495186eeb5e2c29a495291;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc319a4e7a753a36b62503aeb991a465fb67ec5f2301f334d9fbf8d6031e541f613f3f510bfcf5aa2f2e60cba36cbc10905b4f0bf5fa13ad89fa11ea36a72243ef963f872c04a7b1d388e4cb1bdff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc57705e11420df8e8fb2a0c5a788c159dc2ac26ff42f5d825226cb948bff4af145769760b05cb83cec5ee20fecddbfb58b9ebc94e6845a5fef78e5eaef7757c867a2fbcc96403c93b326d64f0b85;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h603f1e5e987071581d0fd45817171a0013dfdfa85c17936590864d2f545df33ea5a4069046346acd071e913c41f57ea5b248fdadce881fea999085db925188ebef9505a809f3af4342b880859a52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf120b67ee87b7a6497c1faede43354ba125c411d26825f1c3f8bbfb214f9346257d1c6f947ffc785a5f06b86adfb204c90865db8e7edf1f79c4f0055a3d110e994674bc789a8a85adc373e82b87;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e2959bf8c2cc1a911914e5715bbe4030d132b5b0bb5b0b7a082808be0bfc2df105f64f278f5ea481f44e9b5c15dc3c44c97f540368cac25e0ccc002ba0a2ec09dd0e73299b3c46acc4fec8c46a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c74c0094c1a874ff76a8735587926315f2786cfdc2456492f66b8aaeeb108bd941f78e684729fd9750f64db3cd5751d165de4da7aaf0806d4d5fa7ba6f457a4c0f1ff0bd6c4dc9529036b27d56e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d1545dd31a200d8668cc5ac6a2add0579d12e7a3f6e1ab0cb452608499d63daa1cc6faf149f0b14d2c3ae58349272d05fb191442c4cd8965935015259044ee517ef40741e3bf8fd46627c2dd74a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc84af3c7dd3c7efd5bae1d5e46acaa79dea66beea6279cb5c5fc346890e1b8eeb320c49881e0a53cbb5b9414ab6b8b4dd1e3030487b012d988f967c32c0392c33ebcda032c00a1a96f6e880a9056;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d0f3be732e69fff592f629c9a97f554e30bdcb892f65d9a984add7db028595f05df227dc29910561c2e0d08e7aa65c0882f8bdabff1dacd3a80062e0e75294eec89bf5156175e739def262ee56e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1145cffee83d39a59092721dd6b1da5b170338044f384fb09f8d022a784bb7a75481b1a66a39f894b0b566703b331976498be33f57f8126932d84c4b9b76dfab310b367dc66a18d55c97641094e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178bde85988b68a0615ab0d2a8c1515baddb32b6d69d0045e59b55fed1c719dc6d63aa259fc28f7f1f4c935a1462fc4c3e9b90cfb5eacd5347f297a8497f8d210945f1a389b3263a7980e5ed827ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e9e64e536d75f122e94e2b617df66918d7ae909477d70adf8ce4e4fdb0b06225da28b72bd9183f595eb8a9a699effbc7d208e1506d3979b63748b3564e7d5eff1a793ec58d19e1012a16b3313de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103fdf1010a1481c74c0ad815a80e8adc9c59dfc94246d52fe8b5333a6fa812fa4a7fd38364f4f366e864fafdbdbb0d390d4d8b6b16f8259139b6344477cfcde06ffc31a04fa64d2c70528b20051a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dca3ee96ea6d789a7f44363caf6d357447e4741b3c75a71dcc46fa118b69fc2890bf5a96cde675a5702ba9e1feef148be3876ba30a08e2d515e87fc8d22321e1c9822ed7d821e92a0b7a716cb823;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f17bc1f9142276eb572160aa2e89c683d9c6fa28f5d4835e372e3db5393f011e5d1dd29203f086545b4a6fb2e9f6ab0f8b7fc4230e07b0bea8774f88287fd18e4255b02d4a0cf3cfebc9d9b95f47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h988dba38c8aceae5f998760f6e06bac4c5ca961e339654d00f86c6ee1b36553b1d9a7f7b9060ac8ed7609c51dceac0abb8665c00c72348c91dced1cedfd463f8000f700a842d165d2bcbb1a10c02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8de0dc6b510d37f1e02967eeceba5f0aa3edbd6c401a258d80e348a5d218f30496a727683bc2dd0f52380758524c1cfbedf95fff89fcae6bf95b43f398b713578da3945f900adbd9e74079412d8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe1f83ab50415267e6f882fadb3fcfe320dba857683644ce9b525ecd87b9861825b891262b679eddb2112a18a818b8e27ef1790b2f642a97e676efb7c0dadf52ffd073e38e85ebbc63c1863e36b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adfda4f207714e83aebeddba92cc76d4eccaf96d8603309e89fe264dfa7930c0c44feb33e2a03de90eba556dd36fc54863f29f1cd6abbbf580afad2d0051beddebab07c3f9cd15f7323da2adb9c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h366d91714708120e734c9d81c1fd99893892e57c1967255e6c99dd905ff321b5871bc2490fd01e0a3a0a52c35b07afd59b53172e652df0382c6d9b7c3ca9f7054b0827a67bf5c882d61a4babedfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40d767917844c7fcf67a777bda58c40dea990c63b1fbf32d19b0d39ae7c7d744df2d41959389c25bd9d32cc105459c4c244ad75103a108997c108e37de63fa3a4dd94c6c4908363be67e0760d757;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7be4fc0feec287b47bb34f5819267f994ff90eb1a38f4cff6c2309006f85d10eaf079fb42415891891b47c582d60c1896b3162c100be4f6e0c7ef4ab2d23ec14fef3d73a6471e6ea4b517ed564bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f971813a45de5ed133907e178908ca474629dc6edc341b67d059a6bf4bd5d0e8fe51785c513d996eca63930f85b09bab9693dc12e437c28116ea73eb855e8e87e03314b4e28b28a128ae6916f8dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1379696336110607094e21a17b2ac802d2239a3e1e9d5c62df830aba6d2935d7012316662b419deb1d8a06d39d0d638fd7567d80af260c5d3a783ac14c6832a2e65d2bfa62b3107ded7295358cf2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b52aa9a5dd6241d1c6a1ab4938cf5bebd8d4bef3c68679dce08b612041ccf20afc0afa7ed55ddd081e8d3a870daafbb5df294326da92e556b4ee4dd681afbb97a93a40904a8816871e984fcf986;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7c369995cfdfe6b6d33e80102dd5ed229cd7047172d1730f466a8d1089129ac23e60ec19ce3c76074cb7c251d82d51cd324f7df0c092c724b96b814807915732f8e78985d9de263f25eb3c0f413;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f767de8285f8f9fa04b6b18e2d11f4598cd63a0d9a03756818357b7132114e99396d6ec0245400cc34b59a0862ce7c2f56add85bd2be318b067874199908f61534295bdf51c1138f9a129c6294e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc67a74c73bd50c2d5e05c740dbfda1ecdbcc30f442c377fe383b7373a78e61436bad22e63ddb566f4dc69376df96e013a210a56574aeb203756ebf14336a6595c3b9efac10ba1700bc8874ec6a36;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4605fe3cea1506e439b093019d0c5e5eee70fdfc9c57bffa58bc37ee8c9aae49209be4f40a53f599e96f31ac5af0764e6322cfda5f53debd87d14cdacd456884708161c5e0e74b967605aef2137;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h207f3c0d42bdf39ab1689334ecb02c201caf6d412f27d5e252e6830fb42043a53d57711d475684bef4a54399e761a8758c52b8a90a8066a1e2fa39d907d3838278277cd3cc6de68d831f10774476;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16637c0ac05bca3bfa6fb63718c466cdf4b3ee1cb7199e9378e9f6a26cd6ff2a591a76a88c7259b87e591b0455a8baf4dea67b1e4fc225400fe05233f5b4ea013b6eddafc782043a0a41849e3ca79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66370e4272fdcb270ba4262db9688154dd445e417b9eeade85c09adb17cf3e31c12061ae6c775ef48fb50e3573b1cfcae7d10a6d4967c211d49bb65e5bb52541f36a60e6d2347f71426d44e303ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h371bd0bedebf33489e5df4701cd9ebcec03e66025b9c6d4b77a03005a18927d2b8a9989dccea0dc05c8d1159e46071965356552eb5d05428d07589d382f78d7a05aad20ecd739ef761667995ba67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5b01b60c5f334b23fe54c2de37d513a1f585abc7ebef33e1142311d367df022433e2132d12a5c3f9b40c7b03b86f25f49df4d2eed006f297ffd6855b1d0ff4c897ee0c4a7e6a222c927ee8f846c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135e6cf5d78269ae26693057389bebcfb2ae30e5f713468a15ce091e3da19a7dff6e69e7943a5e6ae437627d9dd0629c8d780e01409f18842513be1fe2a2784d553e7e8c8f1b8ce01cc7e990e3b6c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72a515cbeb36a52a19bafb6a0bde99ddc94d90339876e5e53c0dd87c52bb4e581e1dd132fa244bf78c23f0a509730d0a05a411889e463ec01b75bd170c9aa318691f504aa33ebe87ca0ebd7413c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23cf51a377f814dbb09d29977561d7884023cd4f20ccd6c4cfc4f072ac46874e5c26373367906105d99c34dc19f1bb724af17366e4202e6ede3a0fa94a1fa5a17ff77b6d77649fd606be1b68d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ffc998fa5dddee900df366010b06ee4da56e1ffe5406d2552ff0cc6c5da927e7518335ad421c67bc147b132063181e9106991f83f74095aecf7dd3b40f7f2da25f6a57dfe2f99ffba8a4aff2ff7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12367c744afc0886fba2b1b305e5615928836326c7bf629bc3d905086baac21e0e4ec7d626ee1ba8430f98bdfe89a0b1a45e4ce7cec5335033703a9c416ae85c428370e5c03b40b4b06e80f9166dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33d63006d313a48591a96f3f2e581a967a81ee0da0f601aba88c555fff909e5069a699d881b6c439d39293c10bbbce09a0dff4a0827245e34ae5e3049e2b2901b2d717d2249045c8e78c794a9e70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138dce4b7397f48a4095bc904cf9c950eb3f3bb62f551f12a660205ec02e1e91eab7195fb8ad6a784972ca3808592883637e178c623986b75db65898719eb773376e936ea80b29e3c5103a67a4ad0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf13001acfb8a4f1a61938fd3763a13451901269029146da91dcacc061a121e90a69bec44fefc3ba2c5a6e28be34a07a84eac3dbcc63890ac9d287c367b2cf76bdb72ea5ffa18773ea43327b76862;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a16d211633d9c73e548374c1fecd98891c553d1995e1e38a0d1ac1316a5516f79d9e9508b269fb4bb5837c643860d943ea76b6d0d11f26c890b848e5c8373fae0f1824d4f0f38f616e56339f877;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10822e75a5462a208efb892bb129371bf8728482651bda3e40cddc04c666585d3c95cff884f903f44542772187d39a377fecfdd61c54182a606bad491183d47f1b9b6280bed917cc4dfd34f134ce7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e83f595a29fc1468224c10049373843a992bff649b38f840d094414f71b5e116e3d00039a91504f7e36424d2e13c810207c60146312a0bc36af70aa1ccc0561a2fd05ce292859cdb40fc20779b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h958a0d62fe48756f96fd7858ff6b02981b102e6a33980d0c0f8513a2b7eef1c12f287f363fb1c0b9e9ab71d2a0ced0c452b788fdb7343d8fd0898f9df98b9a9dc1b1e9dc8e4579f4e030beeced8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61e3fed4586f3a863a59ab4ac6e9a0181ab7f1a7e85ce73732cc8bb0242827c216a89d28479eac3c90904630bbf850324d419ac4c1c0f8f4d924dd7b23f3fe11b8885601cff95bb39c2d1350c352;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h939e7c00b61d413f41c687919171f57d6234d42ba63515946a7af4a9f619cc2366a30870d82a8cb285cea1746ec4c87b5206f582d95a371f36cbf06504593be33c9d7138bb9c2b147c16499c1672;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb83b0d59598d040e0166b559c0f4a044f3678fb8cc4cf56ea9dccc55baec081663f6b8b90fb9d99e21b8d509e85c38b088d440285cd897343df28bf833ecd8d669a9c9eb95ccf3ff9d1aa8791f75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc9e721e61ed4ad8728c87eff8c2dd47123a9e2656c94e9c01c4274ad826c79cd40220d19f935f76bfab2b8a80929f3afc4f5db50e458a346f1f62bbe3ed8b5f6b8609be9acd2b14864177b72adb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173eb760f9e3fe9be96aaa75847b2a869d598d873a1ea706574919b34265e6cca7bdecfdb2b39bcc19432bec6b0dc4de86d70f3655f8888fedd3a4e3f96666d420a7b9ef33789e2f6725c2a152785;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1604e935f708ee4be41c370a443443bd04d641705614c656b84cb62781c0c3c900f78b2f7d616f08e5ac3f25a37f29b2fa8f127aabb4dc6e153b251229bdbfd83b880de69bad8e735b333d1331398;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h915abc863e9edd7e73fb8756be7d821e8e04db120ec3c88d39f573f03e71847d2d0bc9a0124ed474319cd4159a1dae0821d6f0c1b88282a3d697cc9fc96dd489782cfcd5b3f94f2282191e00dcf8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c06e805a845329407d701d5cb63b7727acef557c0a17167048906e47d32e0565dbd9defa5f08677152fe346d49b17f361c64d9d2d5a9607122d340fd208e95422a2a00d71063f7f2fc4643b514fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97d9be4d56b7b506cf573a75fa9f0cfe97e3a418c64c6fe1baac9c75b7d004e2b12c0e76a96a77cd8d9a323423720c51b7d57423c27d41ffbe61b2814ca198986efaa1b747968db5804299a461ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b69ccc4fc0194fb681ae4adbaebc3ac237a3f1c4de421a10ed7a3154a4df96e69d043cd0100e7a7156e5f081bf7c9968692e1de2fb7e2fcba91062c5aa42018245223054bbd1cfa115c0e409be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he62048b5b527b19fc012e8ba1de97632c50609548d658f0e7a94886f58c1fe8733de26386efbfad31a78955ab49cf643a5b79584b8b3844482d5a994f7567dfebd563762efc6e7f783fd9c40eacc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda4038aefbe1747a34c36316316c0cf2aa86eb918118f082c719585356c18ee1236383e945dab825611e83ff72b02caa2f898760a60c6162470f49e18d9cc89ce9cebf1bcc257c7ba57caa372750;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6b126cc8acceed5203a69bacd9d4336e1a021590805fa8e6a06baf56a3b351296e0f054dc0479a3bfe920e45497b40dab5a2fa2d05e75f80239da1fdcbdf18acfde390ccf8faca653d391aa949d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha829c01d895c8e71714529e6acc066e2e3297313712d296225ffad9b21c1315ea959e5f61ce56ad24881653237f6319242736b5fb563e4ecddd879fcf5c7d4806e7229f0fb26218e12ad1139f413;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h591c9a66d3b8eb11bb637f0a2af9fcb80bcda79cc2582f7606ff3bc4d5505b32b389d75a99c6e26639a497ded80cdcb1fc26c6637072e1e71d0857767087387c60b0784886de23bceba08058ef69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h257a39a44c7dd665375b0c9d1c19a22639cfc03c2abc52ff40d685bba4cb15745e0d3ddf778c6d98c0e050c250825f26a9100ad3bdfd954e8fe352ecc5ba3c166fc214a148398d27ccf819ef9254;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1988b14ce0944b1571f3147a14fdae5d8f57bc00278d59bb3dd20dead1c87e4f02422b2485e8e8223923ffda57ec659f2a33721c235d68cb8250e2efda41c4786355ff3a9adf6c10f2aaf06d7baeb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd1ec28deecff33b44b0e401c0b1eec0bd574c13b960b50bd943456aaa7fd037edadc4c28e82204f0fde8d92a144222d711177d5371e5252924fc0020ddf2b63cf3e28c0f09c568d747a0d998d2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e80ca7e8da1878db178ee233030e925dd0c89e29f8abe9cae341e7fed403e1fb8bd56f2a2a9bf27959c679b8ca6467330fa1443f963f162a10f591bbfe30140cdbdda2952c508b4f61ca1c32be8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9473a5648220a061f3930f62c5e916241b5316928ca0720e30509d0fb4ae0b250e404ac7d844f206db5de89e187f5bee1f8c14f4856dd3eeaa3379d49821bf3691b58334346d88c01e7df8100329;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca48416dd50eef0102d97627785fc60a073bcae9744890498698df3cabe7f5547179e18371f1ddfe6c601483889bb35bfdf4dd9feee335d10ddb2b9b8a46f1e8a6d1d790e1ad6e1bf145c9f6a2cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4ad48490e2380cda1cb4d444243184a573256244dc1c4ca5a3239ffc203c336ddbd43947bab3b2cd8197562c89db8aba0af423fc8b353b656940b5429dd00f90f94eefded218145164c99164d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a94716e152b7810124b461d9721e713357d70f43eb33131cebc2279235592db8b45daa28812aea459c9a7687f787c1a6b0a4217f887883b30302851e60442dc9fefd252d1bdd5a772b46229032b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc98d6a14892894a2d533c8cfee1d45a15858d914908a66f9dbb3fc1e6a9534b7fe71d4ef0e567632b8e216a9cbf0001ae206a051e93b784d1aef08c621aeff9c6b5ebe33623c0cdc5fb7d4acf4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119adbc8bd849cacb280e94aa7325128550f49f25b930eb7c502377ec5260ce011052971ef9b002ee807aa6737139426826a520ede0bff2e2ccb3504530374041dd3910bec22525ae43da295ac80c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ec49646089eb74dc901ff96f2b51cedeb391a27de7d001101c47ba14bf66b47c813012528c154913b895522d6b0c74e868f097e516bf12851dd62ca32dc3382f063969740b17f16cc36edc85d18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19315090d2c4bf5321ee5bf2f23fd3148087b9ff72ee65e4d08640c655af2c96c5ba8c7f7d235ee2d41364f3a97672278950cdebca45d63572dfb34aed503cf92b575074dd3ec6501b9080f4c4892;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e254d034cebb685ad436ca3f3a369208e1a7a05b364bfac2a862104782cd43991486db1fe172c6e3300daf4408cc9f41f1fd9fd28af2b53a1016caa411dd6fd9ee6438389001b94799cecdbdd44a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1963cea49c956038d2df3589990cd35a2edab35ad998afa263398a1d1ad42cee3ebdd9934cb23ef0c074daa47f1575e5c007b40fd4c5ba654a422e5340c09ae363ddb6d619877e6473a7c2b57a30d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f1937f07c1503cc09d4b121f3a270fff087517e8ec320e1d42ca111dd6f853633d55a63f4fd75456d7d6c220c5181bffc2eb299ed87865f9b5074ec9a8036e43233199257f048c29759043af7f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ea104ea07470dd59f142e6706269d316777ac5cb8997a7819e27571e04bd94ccea31b2fd86d62897ded8626595025a643d778024a80cbce65f4d7933cd0e3d83b8df549e4e483e98f3ac249c670;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17175f9f69a5923fbe187c15818d6410a4b601a46af24d3b029a422f61f459410306b0d05b68f6597940d116424010fc8db32ad9ff0265448a1d3edb7f6f283068827d9254b542d8fb5f8040d3a4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee216d709f2e7a841c37923a082ced364a9ad89c615bbbf7087aa5b1f1a7e1bb1b45ef43221ed084dc5f205e689ad3ac3c807b919b6842a5826416e8572ab36839645830935f26fd26f15804f3b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a42c688acc0c556ca4bc9ff4d5acbb3c42e0d265bd845b9365f824e9dbbb08de2888c9cc4e0e11ae46750b013a16e4b730fa13d421afd42df295fa8f0401317bb1aa53015e244e957b12bc50853;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91a845c4bc2f9af6b11cb41188a5a3afccd6d247167f0e5c65e926cf844ed3d7eed46d3ee79531077dec0de5a4a8fc441df4d3f2af3119ef9e75cf7e1e1fafbd8593e350bc0c6c2484d6aee19402;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db48e068ccf33b841542a59e650eaa93a649cb9a9a249bd0af94aefa62d37a6199f95f72b7f3d793f76a542aad5fefdacb28191621f78e9daaf7839d8c6e0d496b36f0986c8c3259316054e03cfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110b573ff24de1556e158095809c1f853bea84a93c7f8426b1b91cc0bb3bfb0a4756615b442fdb29a1d05dfd90b53e3371f4e6ac1f2bad7c16eb6edc665fd32828e10bec95064373ac1f819651bab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8d88da86950f90ebb4acb94b7bce232ddf1a5637aa11a18ae1a920ab173ec6bf55424929ac41a4b5a472c5731119b1bef80f489e23fa4b7db61f986666b307a19714726c5575c598fb7e37e3810;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6d765c6d4b92efcc7317bf2ef66f64f639abf466326e9c65d6efa851fed4f7ccdc3c0f67f69a28a99becdca10da55f883fa355015fd69a2ec25b1054fa70534ee9fc0a07778d87fc712a7eb0355;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5d24e1a5c8cea39179c7278fc0765bc996a6912a096a98bb08335370bd386320eb079de86607954bbb048a59d6a9bbde1cd3ddca534232a7d1542718f47e866ffa74b2571814d29ef6f1371587;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190a0f9e5dc92810740f0e684d686670f2cebef193e3e8cf3b0eb1f4eccfc7243c87bc6dd2e506e761847aa5c4a3eb14ccaba4e2565ee587705bffbdc6003db52fb8fef304608d6a20ef284fd5633;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he94221ab2b0c6c96fbf183fa712b205715f4b4a66d790fa1dad03be6093ad68c84cd57f392941c43cb3d1d39b2efe08a502a071536be33d7eb025072eadbf5fcb139f9444d1573056ce97257889b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172f3fb7280fc1ecffdd60c83a17e62d55b4de8e6f3ca38ddcccbf9c652691ba7446ae9e1dbb9a80ae97abae8311b969a81f32a1c31b5f256567d9509eb6580dca1ee312c55c26e5162d1e39b9e3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf06928cfbfa61ac0d4edb0850fe5ce82eefa0f4dc06efb146c86983059dd07b38ac12d684440e1cf2aabf12198d541548ec69caa00559abd5f3d407e9e65171fe661edb51b7e7545976cf650c33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf41d2aad3345d062a1b82d1f582c45c37787b37a0b66efb72999393c6acef8b92988b39ddca1d0a4fccdc45ff63a0cfe556f680c27fe65a145d6589100786d3c22837e7e7c214d1ee5f742fbe23e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6e14d6b835819d780a51e359b457f3fb758695015454e320acd55d5ccb5a364325bea07ff20a3a861c9062616e38dc1d00c3be00d012aedb0543e9e9bd88d6f1226bcbca43073471c01e277a64e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fcc689ddc405f007301c9332a3a79322e52d04062f97fdecfdcd124954fc1724f72d5ebf9fd58868e5c2924fc562861821f22b4baf51a269d8123f6dc6647ab17a0a93f7a60bb469ed447d13a39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c22031f6b66f7a64adfd482fed09bba3b986cf0ab19a9781030e765ff6338b8365f79d382007c128ea75e60d9f9c6d0492fccba7d5ac9a4d4c9318ae1d01d4be80f02456ab615c1fd05575b1f663;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf46ddbc0c35d123b8d1c1dda09c8b30170fb5879610ab6fe86abeaa65701557abc21e0042361770c8c4656b4324838cf8df011161500780656874d0d9ba3934f64e7d1dfba15710eebce589af7e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92e10740eb29bf95c19f8e9c296bafc3ca9dc5dba6f2e91fe4cf953d576c8c0bf9a12b746267460a21b28996048772ace653080e899149f5599cbe401dc8102f9868df39351bffe6a34cd5bed473;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16744bec87dab9db805e60d4f8abb177acc0a036ca4ccee59acc8847da42cb195b345c1a5baaa63a5df9a38990909e83b0c11f6ed7572f80a546993755745f0f5b81cbba0a8e96f45c645eee9bda0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c4bb480fb2bc84674f021950ae9c95ea3dc466b5df8b0df173e958b9adf9e92a047ce3b2cb6f7f964fdfa8372f117432a234cf390eda9ae85a0815c5cbf2aa2420fe67c581f68b8f56731407fa2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1190fa1bd81635b3734e5b153cdaee904ed44eed44d667592d83b42eaabe52e383545dcbe953543faee831836d731ea812a3f69f4ce9ee25fed80bca5b624593124fbc38c06bb6001af48ec3f23f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17226ab2766b98d475b9ba772325a151250348637bfc1cdb78f7b41ef2a04022c27ac453b24d67f13191756e361b71633bcb5ab3543df09a0395673aad5a37afc28bf7ad61653a37fdbd8d902b025;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde8cd492438bd3ed35dc4ab1734274bc0bd86caec22f0fb9ead212bc00b53fba7f71e17598cb1741edda57ce310899aaf4a7f291b40db18bea2224af4b4d469b0253f797d55a534a480cc67f8d58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h458f6a1a0cc007d39349c1f1a381c4462dfc97174dbbd8b3e727bc887a54bcad4c10f099285a129705a9748fc266a8499bfb94140c017d730db36de43dc0ac33dae80f7eb82ecdac7de8339d5f22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h949c646e3d8d06899258deecd282c9251571f3f629e5c433c9e480bc06ed50a8ef8a90210a19aabca707212a373f717d25677d381ed14ba9e4aebe59dd1f9c60fe3de413a5199e7c27e8891d65c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h543fc26bc3ae56b9a9bf05ded4f22a49e402a912da3318895113f6da868aa9a6a2e4a3ac0846fb311757aa4811c3eaa216a3087389f3ef51cdee1dd6580a1912761088c0cc3c3b942afdcc9e0104;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1982644834539ecc5cc813fc52b10b6c9f2b16357993daede9b3730f1e901414cebc8799e8e02589cb4b4e2a254ec6280a275cf08a9101f6d2c9053c428728dff9c2c019ffb6a82c2a54984436600;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cdab0deaa680f985203adcc32169881208dff0ee793449a2fb8303273275abd1a90f33cc7e9ba3538c999f9fd123e79e43f2b17415920cde9e5a9d16af39ab12106bb80bfc2b53a63e7585921907;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14904e79b1b9e076cba3e655ecc5e67aebd7e94a5c2ffba81e2e2bec8334d3495925888f4e5f78b0625903927d286dd59c8006b645df60523cd4673fb6751fe1c2aa76e91f44ec514387b57c3100;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb27471eda1aa50d9b61b9132194f006329564d7c5946f02e6e6231975cdac5bf2717dfa194882b18f1b8f16ca51906b547b67bdd64195830b44408859e82ee85f6b698fffdaa44b4f9e8364e47e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d5d09eaa4a66e2595a8be3acfc55b73d86f44d7485df867d46dee954a1c233d4490c172e6e1a3b609db33d36145eb69a0aaa6be47117ba1eae1d24832ce17b4d3755105b77eda3505649b0fc1c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3fa393552403cc6624e19785442ca35ee5de879a1eff6729f228800133d4e6d4a4b6ae7ec0745e426de39ddbea6fe823c5f85c259fc711f20c4a654598613147bb5db2fe8ffc6dcdc7e4058aa94c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f7b4c776b7b1e69ba2e966b4d4121ec70620f2cc578c48080afc106e1f879637b029be96cb0604e2b796a492a653874791929337f562302e3ee3e00a1512da7a678b3b86608e5efd9aedfc06f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1455467c27378c6cfd05f41aa010b1ce6712a2fb898a1f8bd1367afe3e482a437bb5c8b700a7d1886790c217a7033f4859af97d9103acac0c8f978739eeeb9140e9968ccf73f58f15c979633b237d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e2477ef7679253619b3032d0f4b3d9b98d3b01bab2618504ec76bad298aa0ec4283012ac59e9e710369c35f51822d62aaba0eae5d1fb3be9977b0631a56964329c40168a7c188726490fd99b1fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37e01ae9c1515f5859339b11206d6b537351ba65883be939d801b8bace5e59607ebb07a26e21efd497efffd622a8f2383f26aca1acfb07f4784406923bc45974376676a4640d0b028ecdf6ef6709;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a21854359f53a8a7465f2e73596f5e418f17caf02e96ca9bbe1568d827b0c10470eecc6505217344f6cf02475bed45a407a385c6d89f57af71d1dd1c206481f4f583ada3376eb82b8e0036816872;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27f56c662179d5a2645b0ce8c3cb4b477254bf0ff6ef9e446b386a7cda6a1d0b587a67b3bfe56586037603eca466f8f5c308c0439f9923ce022269f85f0f40949a73b692d5b355e00a51fe20b7be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7692b017b491b93bf7250d706a21265b4672808be32700554afe83c221ebb7924fbe3b7d703e946f6613216810bb43602296227629052a4f816458747d7d6da9fc7f9e688aedae040dec4cef8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d07ae137f775576a975865ec8738c13b7f515325f8177c790df0e9e730ac11c34b681f6834de5da50558b21f8b98beb5a54e1aab4d1d491ad4f118d1e944d4a022232478418bab93010620b38504;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe3edcff2672a2a119240a401a796015f0d58be3d06411028f8ee87276e3f7fbb591e37fb8ca268dd84d9c6bc1a0548855088e4e50d517cbd385ed916201badcd1706654807b0e91be960d2995ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1c79ae9dc605ce6ad0c54d2c708e8d807002c0e42ba11d5bf8d8f4d3cd608656758572cfdb899c727ef0a4381aabbc89b8d48f479314749e65c05574661684c31a6b1aa57ca7ef8a8b70a7db5cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167499fdcaf48bd489b4260fd7ce5eb1dea38d95238c5a4a60cee806a8b513ce4a9c40309b7709a77414177701359348a1c7d5e5b02ea92d367ef80ddf3742aed1e30943b07e0a9c8eed6fb686b79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2fbf6bb07809ee94eb8d83a128ac6b819fd9c2fd664fd36916e6552f3e2334100bed4b41475e7b3e8c9e83f6cbac3ca73e9eba27e12700b2795bd6d4e916b36594aab8f6296ecb06ce12217d3bc9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c38df5d530c65fc1581b51dfb1198a558692262ec561d70813e2445b4d85f14e4ce3c8597a924bbef7a41884d4a7bef81a6cd6fa8a8787dbc1422ed886b866070eee364c67207f5550a6fef84cbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea7643443aca2e6ef0f9ae4f03fc8d04b3d67a588119a6c4e2cabb7038d7a6b6fd2957de5191b8b652e78479ffdbae5a6f59501264b855814c3ed1b8b95cc5f75dde033376cb9a0821e16062fc8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he24966014d94ac2f2660358c417e56edf56c06a02d324fc4f6ab8471ed13677c61ace387216d1786948f6f8239c24cea6238a1de0b40b1f050a01b5d183bd3bbf741645c56dd9593b42f3d3efdc0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc54b527393e11898eb61e0550e45c6aba62b8043da6cd81f4429e8a44569db690a977cbafe1d4f7919917c33393831268c95b2aae72c3832da48e0f51907b0c8540412454bf30c3d58a107e09a3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55384cd0f2e239b12cb1f31078f418f25b86a864fda2ab49f561158e63094ab7343c9a9234a60c907bc1bbb2dceeac8227c149dc039dfcb5d0dc6364901494e2038dce5441f44b4d05482606f622;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ab7d8d8c0345f586488747d5d597f14f22f7ccbc87aa616950ee10ef5871e599a8cea0710ad3981a1bf190a43ae68599b96dbb10d46fcee9f3f270c7c27b8fc0ea3c9e9bd705e0ebd68b008a3de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd227b2f943c70c6ba6b02e75fd3be78b50599bc03b031860a5317613abe686797caf54c670fbd2b6e07acad1dfc44847efc311c395d84002b2a9b28f1e75bd2cc2baf191a38c89e07123aaf7e4a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h828e011a62b5d3d4bcb3974e024b3615f2152cb19a2d19195f08d78d6291ec05e3bdf63f93f3d29b754c4ab7161009f970527ce7fa134347320aee452dd64aa9ce552d7770f8eea4ac2aec02cf45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcff03cdcc8499c14ebbe624502a3b1c2c4a62c7f981f84e763be0a7043741aa7e85a5fd40a3f04ee4f76f5d0f67d8508b6a1f0507173aafcb7bb7a14bb1c20d4d892c5960e6c25f7980ec34e6f77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a5dc63817bb64a053c7d7e1c3b92ed32e8afcb76c92c2f1f40073e3ca37fdd775c7726819debc760c5a60c4e29d0ea7cc11a8f5410406fb46d42703a7091b936fdccff7ea4be6689913e15b7fda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc8e4f17a63592bd3bb65b9a9858cc02bb28aa197213e77758bf87252d9af5e9d328958e0860e9eba58e209827f00a77460abb8255a207616fdaba705db9482d3d5b8a6181bcb574e9faa6ba5bf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h394f9dec7f7d2a199b6a17692181ac87a566b5a29b61b65cc01c0a26fe06d3919799180238a51ee6df5f557c5fd99910e3782820d2e1e0af35f4cc5a8ce0b564fd96d5f316671d422e2c35d796dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12490fcc7ab81867e22117d84dabfe406f83a347b6cfd4c08916b991525cfd32b1bde6b361c198c8fe52a2e0786ea614af0c49a260a5dff0949ab173ab469adbdd41a355c09a3d87e71a1028a2bd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db60d5248e613eeb2f0d0bc023452df0046bf4ab528479252993f9ab758c0185c6ba3d5fd79ed54878e5b4f2f7208f2559edd9bce16612178bc29ed2c54e3ae83a0eb25978a6b2c94a12d8fb0c2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2279174a598f37eb87bb23c0ee5ded50512db7ac168bcab19ad39c720466ce4def67bdb9d7dcaa516ba707be2a77ea4a6b1b34b30987f1b5a3f0399eba81a99e4dc808ad5e178b0f7b841a9b3a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5851f829227a9d4900e65cdcfd0551a226dcf5f6c742d43bb55cbd5f4d623baaf6a6993e02ff4b9105dc6eab466d98222ad6fcc5a1ea19779393b62fbd7682a1000860a801bf0162625fce670c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f727ba645801e1421e6d947483db2bec31af71387ab5ac8a6a2fd852dffc2317bb2bf1681716561ecc89cedaebb3790266a712d9dbf5d08cc7859bdbbd99330b658c3854e6baaf7814719927b38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd0110a7bfa721ce8d4fa66798e2f6d828b569376b938b61a708c9b2b2145abaf0b49f504a73c0b6fea9d087ded0668bc56505093d69123431994d313633d516705e1e6b3faf024d861b63568b85;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2f1ffbc50c9f94cfe8bc452cf96b81aec3f75458ccdd1bc6a5aeb84bba86e0460b9dccb3edd8c1259634c8f3e1adb0678475d6ecacde264807a6c47dfa9acc31a8a0cb787154b6f579c9aa2175d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h984723b5074705f2435a257f47b263ce69aefb68a3d98f5cffcbff87d22fbec074b4f4742160669bb644747cf363a48d08ed4c57092ac6bbd3a1d68e200c55903f2053dd8595b1f6cd842008f06c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b530e4d20d8960204a0111e6f91b812e1098f65871ba25383005ed7ccdb2e65126a6f8f16aea62d1cc9cb7ac658b81dc0c74808d32674f45fe4f18f582b43f9c3ad96719b5b872fdbc27265e772;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16349810a213bb633eea96f00c075bef776e87f28242b072445a4f1168b1b995ec34b2f4736604a755479e42cc8bc5110fb5cfd20c2045a6c07a0db58807fd0facf4c7474481acfc369c021677c4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3380dfb5d87785c37456250f06eeb29f596aac1c5b71e7614f62d5074e8dc81a2633140f2788e54b3750ee327149d9ac1112f3ac42e38123c956ba894d8c7f6ab8773d2ac0123fd5d67b652958c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb955b2ad1fe5399a579cc1e74b19dc98b31eabcdb5f0d89804fcc552550e89eba999082b2a2537c01c6121d262275cdb1dfa1c9ee880e2337afdf286c05de1b75aae829f0bddacf65d2dcde80698;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100ddf4ddd227c479925e825123d37f2d41834a7f85e8233d0ab05ddbd515f7c588337e4ce35e70e40383b008d06d4b081e1bb15ffbbca1df1015ef45b77af210f4f2b21f2bcbb908ec34569ad423;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183c47dd299c810e1094eae87765f4cf6a6229c8ca95d100831aae9b5fbdd4b5f79b877a3d3f69d69d7a61650dc1cff1af7a2e8b212cabfc6a0f66a5deadb887e7a3c052c37f578b1090c16b9cf47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h392051bc28dcf3f292f98636ffc38d5b0d470c9a03aabe1bbc89b7697e513b6c06d4111b5f3954f5c55246a0f633e207f0d412ca19428361ca25b8315082e0f9da293eed812190a677935660ebcb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f28e098c054aac99ed64f49922ea8e4c01bb19df8ed9c6618bbaa3e0613017f7d7ed4b3d7b9ba33ac4ae0b5762ada0991bc3d9ce350b9d253cd6874f3d8b5234e2495f7f24de76e2d0aa3860cde;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4e5c10881b24400de76c179c17d5e6b79ddbb89550d47474a6cb24adf0fe8a8bc4d3a6fc4e927f91521418c87e9ff9490f95a1ecd2bc7e7f3eafa2e903633c3c0de93dba4a4b4c87bb0d4e5364c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196eca1c018ca66382baad7acd35a6e0657973eb72506616bb3ab21b17ca9149063079f1d21150378f651f8e9f28a91d7316f1b9577b95c5b1ad77180a1400ca0a57344363f29decdb393659b9f08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc92c367525c2169ac9eb8b17103da8e93cc8554a4f177b6e69ae1d35690a52d986454b73e27f47528f8af1342d7f7a12cf891bc7f9ec00ffc01719ba6986c7d65c9522c78e31f28b09ef630a5419;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0770e52938ecfa4c558682cc83e61cd1a45908448a1504cd4d490a3ca26b5e0a92a8d99c7b21c0a579a21d61f7e70cf2c3c0c690f8e46c222056ff5e3d53b8017f57128c9c66298a0b9c80f6096;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94ca961d154862ea01277eaaf662febdf6cfe272f320a22e228b7b4dcc1b117d87a4af837ca25e94b503a14d390cfe2058a05f14e5b23dad76a0e1026fb0fad65005d4d39e1f7188b7b4deb1f0cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127c9ddb1c643f2fb00b0ece6018a906416f49fdd3bdc9e50cd8f60ae994aad01701afee7bc168797a457a98e0b85b3502c22d7d107fda26f5cbce858f971fee28c77731246314ef7893762ce1b9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h116449ab9482d483d4e5f95c2d6f8008b7c1f8e2b451e27e6e07ef1593362e97b70aa80a7a9f361e2ce5980628094d3298898480e7157b018ac2612fa03ad38cc017c2489a5341cfe03790844d4d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f626d29b2f480a846ec0253d9ae5391ef969758f52b06a2c902f63a083df2a96d0fb601695a78525e32fa1a5e7ad71c938fe6b88e738239383cffd3db0c9ecfaf32608ff5c4ffe6a07dc9afd537;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a87fd6532789577190d3bba90257ec23eedd894c69743a0cf7f1fa4610d891baf8a592fcf4f0b7d1d1833d52831c735307eb74568acdfef4cd43de76cf1bc869d518325667ec801ae88376fd317;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf39bd01b5a0c0cb32280ee8c73c54ebb78a4c35f8a8998551f66554280e84243d0d197c9e1008da4c9b5f53122ad79f658f27502fb1bf08cd54d94cb4f6c76588e5801c10bf11b47448bd1fa575;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe8e27d01abf9fa6ba59d34cb992298b7d00fc5a51254f8aab74156f6c54f9a344c5a52ee1172a037392043f72e15c1d9601d019070d4a033e3b8792d238ba2ea5329d6754ee4148f28e57b17b5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f5b8f0535a1836f9d4ab6a574793101193602b4658e7805d1f6c10d8ca783a0c3bbe74cb125cd6afb13f774c0d3fc0c3d8b1e0c57950c2f3f981fc93345545ee27b9b9082c74cd82fa6453622ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75d4b3a6e7b15cd754484208c620375ba992cb6e02426c711cf7b4b78b4f3558b98ef007ccc1ce4b4211538f5924c3f33b872bba47b2895d687f58f0b36a7f82eea76aa54d519f6056edeac3dc2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7b6da24571c7f65981a9484c99413f3324c073d523e0794d38a805fe72bb9552a33050c2660c4b55a4e73e31e413d36a0dd73a13c7e2ebd745fd7fbc2cfd8334251fa749e07d2b303ce997d5ac3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6c1d3eec90532276bcf77a8f690c8ae0cbe6a9e07522c84dd65aeb5b7f2eb9dfefd1d28bea19933784c204765534be726aa870f50077acee0ae134bb198c141ec5185d3e6bfd7906bb1e45f58fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hecd8159227bc4d52195b9988ab47b1bc6bad8ad678af50fc3ba75e3d5f34f0b0642d596e7e50a7051b49f4070705d4e44cf3d20a2ec4638876f684ceeb9da7b11253d790fa18a33e71a953e817ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe397c64ffd6a4e36c5cf9f8e0666e19fd9ce71ac9bbcb4043dc00a0a4ccb3baaf50a2d381ee2f1b23af988594cf10671eeea2b3158776ecd02702d1ab88612968a475cd45a97115a783b21c20b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89606cdf1660d342418a948160ccb3937b9c1f1fc42ce38ec0064a673736587abbccd754a3fabbd44ec5cfbd98bdc8b4ecfe8e459697c53a96c2f1f872045b20a3d4f8f5cd83c95af8028c5fb4c0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae53ae39be5a74af4fad7055ddeca8430e05f7f852c6d3ce0fa29b91ee028a2e74023c18bf4fdf6182f3e150faaf66e98e10dc33c6992a003231df0bad67f247f8512a2d88a75852cc42d04eaff2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b728ed133fdb4d9ef8f776ea2997530273140c2788b5bd2ae12bda7aa9236183107d46c3dbae270ce4da3d2f22c6b738da343ba48507980561a3a635b7eb2cbed2c27c4a6c511bf4b3f5ddb30cd2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d18d05150fb9446d22657a4d0a11d3e46cf3b7578294dc767d1d395bed1895cf60e89ac3b6d3257c36f0ee79588cf7078c7b5919e4c01933c1e7976c17581876e3eeb2eb9a4a5e53059eee4f51cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h230f8033d95f3a50512ca82a21ad2d31aca59fdbf133e34aed974bd5927c57714e7188f84688c4c50b4529fe954b5c22e199cc64bc422d5ba0de3ef162bfb7bd2b2e0a0340a669580ebddc8cdfbc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b9ce83c44f7645db25c609c0243b27fddc405a4e68c097c2ebed003c962ba5d5b1e62e9bc2b57a0f220a3e14b0a36dc5caedfcd36d2ac65a9d5fafd76f6cb8651da4ec4c6ab20d36341bca25be1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7625fbddb82fea47798f05be5ed94fd6979089a5dc83848ea13978e542634d73d773453873e7344fd48bbca2a8dd510e9af1b183ae5dc432030ae7a0670f26b26b6d0cebfdc6ef9bdb861c1367b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef3ef6adb1e57b7f4daed8ad289e43fb0d6cc07dff42e9bd8dc5319020e1e0a1c30a1f8339c1c7c3b3206d7f5f2c973fe0daacc1361d5d5e94af01ca8ec7b5fe43d417037c109dbbae7f0d02e2d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da48ac3b9eb6b36c52026773d53c7ebbdd5be814ccf029845f93b8483be3456a9ec17b205b0b91e68a591b22934acc9d716149860d6c4f7f5f12cb848c3bb1c6f90af2cb65247ccd978e5dcfb156;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf5b874d8e8c2e565d5aa64acd345f5690b9b1b1040e699c3eea221c0e0e6435b05318c38f40381f8f222a0b82ed73827839a127c457bc2b6c4b7544696902301ebbdc7fc4851b48108f6e830229;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ea9643258db538a3b31879892e8f45b14184e0bf52e272c24154b007650388240b198e8b21a34a77e390d098c2432d74ef0327139607f0d0266bf567e1a79f89ec2eadfc0428a6ad726af9b565d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b642ccab62e869bc45edbda441e223867777e70d941b42f3407fc8bb5ba89483ade06627df2b511b10aa2399766af3eb6f12fe29c4c0650b551ff1fa37aac6b0484ffe0cf7db28df591fda9853b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4493ea87094565912d5b0f8e5a1b7bd2920e1ed2653776e3458b456470d3372817b947aa096d111e7576e8e6541654a68caf2ed367ce2a621603e328479e26691ade4254ad158f362ace1bb3f3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19872701a921a25844f4f2242333bf78a5a88e6fba853b7110fc9d32b12cfdbd5873a5d8f6923c9d6ac5e1529e1e85b4ef39e9a51ca81af914dd20db215709ab7ef0a482ecdef52deecf1375cd665;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1619ced8846685b3e0163f8141a503b803747b86de74ef52be1eb2e7be46bcfd5f40b5679e2190d5ab36ccfff5dada03950020c85313af055bf8f4c4d9401f246e6a8005ed10d1a3ea7424c79fdeb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a1ce811840e243f3d0b5d818b15f9c3ca4acc9c092967411e2caadc2ff9688eb2e0db6f1e3b483440fd78cb4f2024629badc5da96d2002bd7f184a89a7b898e3872a9da5810a397179d65585f72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11927e738d6cf1addeaea053f31ce0ae7036abfa14bc00c651480514f0ce2d9939f67aeb7948842631648866b2e2fc0ee12f42ac80102fb2532ba995ba5e618c19ee5bc3b8c0f2807bc0705ab7fb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h342f882731c5f84b08a92fe5a9f15e986a5dd5128907566b7b1077c4ac429f0f4c16de654bbce0c0478651382a817f59518b24280bfb4c81ec0cf4dd2c6999e24960a9415f12d88ed5c6727a3622;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77ad758e05a30d6d75ce3931a472c1c99bb6a357c23c9ce8f4a7f12d8c3bcfafd9c02b56baf2e761d9afee6d67b028891eadf1af42c5b897c5443b4379b9e385ba1cf22f2c99961c010df93430d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b629516112dd4c6516c52c38298413aa3dbbdae1f8f13ffa5ec6bd59fb35dad1885cce9359560eaa61c42667348e75c5d79859767560abfc09a665bdaddcfa68964d080914356484d978ca960858;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a5f3a6e5ac625fd56260e6decd1c6455d5dd26fedd9a91bf8d2def5a6eb13ee81267201148d62dff5da0bc3bd256d97f66aa1475cf6aaffedc2e8c9b3d1366cc66fc2a4fc39f16dc71576386209;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dc3565ba063dabce2c17b13d961b5e31bc4be065f2b48091bf47589674653ff9f673230d6c13d83d582df2d2796abcf71bd5094612cabd9f40ffb6e5c97cd6d463111405d5ed729b5ba0fad1561;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12381ddaee9e8e90a2eb74b0720e66500f358ff6f83bb349487b13f85db207b78d9747e4b010a220bb8a76efd472927b19064a5f4552383ff8b1bdb24eb9448d65ce0051fa183fc9d929890efdc2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he39b782540dc5078f7db89873cfcc67823fa87f3fd6c62494e9b0d55571d1360e99343f9f8722f5b83df4a7bf7cfabb4874a1d141f41eb913eb91acd58518d61c909b2fcc4eea05c7aff83f2c5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h160ee1eb16062830cf387b27090c76760603ad477ccf80b03ba0029396c4dca09cefa3389153d571fda2751d3ad0a9ed19fe45ee655f91ba9d6c2e206eedc2fe360c69291b0cf89ae0879b0a3b401;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d6ee1b1767aa65d5d8d556909d959e54115fc7943b3bfdc408993ae4311483812141a4f1388cff5986e2e3b578f24af682cf5768ca09b9e9280194d4ed40bc9caeceec8f2b49e2189ec1a563bef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f119e4212fd688a6308b880ec0d75f6ec6c91cf8732d377676141adc47c9860e3a00182a35c642c66dfe89f243cdb32361192dfac3e59503e599d4e084adb77a84520919716b80afad8b6ffec8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f56cf31e56cec8e3b3b87222e519fcbbffaa62bca925cde8d20b36e8d8c8af71b3d45cac3d9828dcea2e9ccd91c0040b04063f508602ae029198fd736c1664c15329995d038d56c47e95565747d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63f91089ad51d3cb216e77a0f9692512ba1dc0c949fb887c695bb8c262752001fe1f91df621ee83a44285a6b6259e436e6ab0d8f1533c74011cdecc83a6ce448b974ab12ca3d8864666af8292058;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7749dff07b1ad833029c60899ce9ee2e7292791ea2f3caf5d0ab2f10ea4afbe5b46faa2587a548170e579e67df83b4d3ac1307cd77aa63a92b35fc52d8a4d47a8c4876dbabf5e38fe7975873d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fc1ad992d713ec9ff4922a9784f93d40d1b2d64de9d209c228de5bb1a923b44a279c8be2ef155f49cbd1e95620a979b944bf88480770cc544092f5392a6d6b73afb4088dbd79e7ca6d730a6b564;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be88f749c0a7b262e3d4cbf175314753e5c37b1f3bdb752cc76bbc0d8d56816cc5b3fab9bd08486671495d02ab3449c6d99d1f3c4b81ff796abf8535887f7b370a4b816178ae757f7342c029a999;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49035507d10157730b2fd5020d558e5994c80476828dde2b0025de49581dfa2889fab74fdfb104b696063f96eb41df34581995b709b85b45bb3abc6fb02596c0a5e237e40cacb8eaea42f3f03e81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68cf09b925b558b6a97d8a87c74d3f50c8e90693092a2a9612fa938943162b9ad6f090cc0ad2ce963f27a319e09fa66dc1f4cc5ea054cecd77ece30c641f0a51d93b8ebf51b9bb62ac572893d760;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbce544c819c8dbe170a4737476e9c39b55e489244223d3552b7149f5c6bf550ca384c8c18d46e7ea61a08724a2d9e90448ae5f48e847dc5d810afde9f1ebbb0b19c64a77328156c42cf0747b3eb1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1540d2a334d0ac58fed0b13b5533a9073a1cf6e152da424792b34ae8e8d7e7e4fd419e496182e8061746a7ab12eb8d2b14bdde22b80c5031205acf75d3055fcf5c7bee2250ad6a8eab96122278d93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164ae037892089a8421c3a0e6ab26682fc0fb4c53fa179acbf451fd67f019e770ed309aa255163e9560b39c57fe4a6f44f7cd0dbe9a1df22f178b679925c0f7385857dde1f354e57c70826fc69030;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c20e3feed28261b318669bc1c7cc5ca41e4c341da2c050438844de40001abab5509916b34cb989cc943060fafbaa7e11fbc300dc5b193272f0552e1818102a151fe876a2ddb1d1e6b797de836c29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171d235b15324b702ed0e9e9847e36f232d5cfe7e0132d5cdea042966089f27be45cd8be81d2d697c494535e2d411191657c82339ff6a434117a5872671ffe888c519e03741573438d4954411ea8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144c7e77a2060334d9286313cb1f3207fb69d5fdc2c1c24bb6f8a155f2e9dee7eedd59d07a848ccd028feeae8dcf2c3ef19bd3e61c0708d3c82525f1d005e3a5d2d5834f7bbf2853099565c271528;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9e7519410af061fee174674cb38b24e46533fff89360c83becf8ddf2ea45bf51af5bb51c20e9738aa55a89b36f1096d6b2da9909589f1b9bcde436ee08151d0aee9e838274bb6cf916189baff0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fecade63d47fa5b61cad8b569604fbe2a8c656b4e3f085c13b83599a992c46ccbf48d0b02042e8872a8233db7a455146c11f72e4391badb5ca4cd805b34e6243996b4d921450305c3f159db17bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha885b3b97d9a31005dcdb3a0f358661bc41036ab31bf5f3f172ba0fc249681f17739bd015f660f56a7243c7870e97a985eadb3b80ff8ef5baf83fd7bd2d76940dc77ad24a6d16d0316b3813360c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3b39ec0478c8d22c41717a71419cbd62a74425b8ab5d235e7fc64aa1f6330f608a3236802bb5126e20761e5fcbe6873fb634df10fcd536dea3153f20d67e923f7b7adb00bfa7ab2705f0072dee3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3f882379465bfd696e594968e3b1938214fd5541c44bc02990b437ec224da6a758b0c5e5bf8da0c155672ac6bc0145986436a18ce1a182139a5ce1a63b6ea92e5de7bc78b26f485dde7591140f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e43c8dac8209f3d033aea9b5c4526d38d7b19b2cf3a686da582308a3ca75eacc813384dadedf2848cdb3f69bada7dd977c01a254958e846b45a3e27c66dc42842ce8d28ac479ae5b5a25723df869;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he80ef3b0c8f0e2531ca1604076dfca1dd259b539d7dedc91fb6fbb36c811221da3a65ccc799e2685ef196cd1f87a6c5e70a0cb80a4a00a2232022e32ce6be421f5d20f19619c5c766ba6e6da8e2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38430113af965d58389264e7bb6ffbba971a7fd98e0198214b4129a7c66c64afffc83d6fd9fbec13665d48eb4f1490533fc0b9c2fa6db2975288e522cfb04e769997c8a918338539cde1e7c768dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ba9827de9114247d73bff896254d90026afd6a4f17ef0ef325a8eacf159c40d36633672c54440d2d123018d520da97a587b3005dfb36ca162251b613a3d3a98f5cc430964d56b2bf3ebc8385b33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf77e67c8b2694b6a9084f7da58f7d3610e2a06d3af1352cd6d9b81ca4c6c4983e5efb658675908ab7710a201dae70604b39d775ec564dea06118afd584cb2b45c8bf20e13c4b181de406c9f4ccd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6695c89ccc46b065222c8c9b16ca62e6003c1551bfe94b0e7f6f5833cfa978ab7952f0b53e303cbdc6ebb953f4941fcbf21f0b78053d6f32535bc0b481d6312d086f519e1e48c202383038ce51c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6af7439596649b843bac7fe7df6d6d9179fde995bb7e310f4e6090ff09de9e355f8da45d9f506b847b62714afb890d2876fb91df85a39da6099208604568fc8b62a81fbfce409fefea77822f2f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c4c216824631e7de9cb14006b898018558e4e120f9c4c008e7302f582f195c42b368f56af4ea2e4518e9ddea3b432f206069368b74f3206b0ae10475c93d75ce253315a40d04977647d043c8e5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd0a181bede4f6912a6e4798c2db5e2e2e7ca9955142bbc41161fc09fd8d95756f2a020ef7b0992edf1d0e0b4703ca7a67a96fe3882b0e18273ba560133fdd6fbe2182f21dffd9458e6dd2ed61eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3da83da60c606c81cbcf206555834b15f236eaa6abf36b3cdc0f7ab3ff77b2583a18552fad8c0740f51b2f2c6bbb778eb67257f83aee576e8a2c0ddde58a4fe3223bc32f3d9b3f43847382c911c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37f592f0df34d2c7079f5f16ca995775f221a0d1d931de690ce3aefd2143bd9213352f1569bfa0fa2583900c6b6eb83d60c5938619066c4de8e4e76834d8ea7387a5e26e965c00a6b13880ae96f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbe7f23c7af8ca46f53ab58f9484c95990fa50f466c51dd27c9ef07a72047a5c121a88b326292724b6925d26bdc99ffa3aa38ef3bb774eae2531051e766777168a95c2fe51846602cd69d79f0ec5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3de3cf214703bb9c4316a57a90d33d973f489e74bac4f972ad263840f6b98f0c766998f2626f7b9cebc6fd789f98fd3a84b06626f5ff6a29c28b30d2fa3a92c5e6e3efe9b271177972db02fc0bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1132bd5ecf6a7dc4d9c7a850356e4c3e2e514d6b85267b1d9063b6274ffcf6b4bb804c0ce35adcd0d25604165fab5e7ff8c68c5a72dc847f14ca6d186d89e06baa1b5b086172e57e49c03482929b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee848dcbd3a41ffe73dfa039a11c71bfb8633befc0e27f0e929d3eaa5bd29592729a7782638b1ddbe8ae08c16232a5667e79e1929ab45e6da2428d9ba62ac9d50416c19627213b19ef9577d12045;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11fe53c0ef823f6e8057cae7c44bb38cdcd46129c2b4a263f6b309299b86e9d5b836f67e2703132d88dc01c86c8f67979cc5993cc78ff7c19f4c7144027ecc116b35b5a5a8f84e1cf24d10012e49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66a2c2982d21c5f4ef9c0f1fc8c9f1a36686b1b3cdea68400d02395a6e9428b93e3ac816ece9af03a44a611e401d001aebe5e6471422a4e85bb64b13ca161fef0e0577fcbde6306f8fd62e3de834;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be9f91723d7f6bd8d77a99043897d79e73bc6b05a5b4f69c82dfb9d19a9274531513b55147de3f0a842c97e61661103a54ad2540e9da1904a8f2cef0931cf7626ca2fc649fd7dfb3a3467bf6c2da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2029bf8f960353b10e4a932482d7a3d080798e3bd4106f8495737ba5cafa71d2373033c4afd23ab9caf4179806dae13c5196d5613ad1a756ba881ecfa138b724b5fc249dbe826bb81d863121615d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127b7285f314af457fee1f8af72f67acd2fd72e4163bd9b560cb4acdaecc43199c92af3e95f983a1d670265b09ccd87b2b2dfcfb597d5d70be09b3d1815c672b4539acfcf7b683df2e0d98f7e06b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4331ca6e9a26f3fcbf66451684a16e069a81c9b06e105fe7f3d86b098a6321654f00a0bc3dfaadad3d51d59df911eab1d28906823c06e5b20fe934cf28ae5a29dc5bf4d828f696b50d6b25cddab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h340893d92fbdf07e1a273f0943c5ba9caafdfa121b0bf09f0ff33bc6e42c3dae11cebfc87efa0623f646373bec0ab1b95aa17682686af6480b818b373be70f0bb69e60c0ab94ebf04eea845f4d09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19682777c01d01ab93803c3d90dd99f34c87d401c9d1d6343ec1629c93d94894b68e5f4a17b8f35ad9558c8f33786b0cfa6b972f98e96bc071d62722eed88e00acacc748412d008cc68d8ffa94136;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a999ef4e8d059971dc17bc15edb9a42dad7e9dd9d705a964ae49a20bfbf3676d0381bb4396589097e795c97d22f96573dff19b945ca46c953082435bb5db3defba64036761291b9b01465c779cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc0f25d7ed8e0a6d6b88e8bf72790ec907727a814f4ad0afea84b71b4d555e72c7e29339289ac7883f55b4ad66ba7f14d1e373b7a943cd39eec3b82ac63c496c28c01d1e12a9e9668d553d11a0b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15de873af6fbedd7a68c24ab5156e9f76998b49e8fe2d41321224d0d8304aac049be6c00de4efba3ed4a57e81f4d3287915f81b27c4c461bd8e4fcddf24324be390140be3028ab827c29e13833def;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1131c402c14377796a702303ac6a335c548922084eef32a361d021dbda6b12fe045e97bdf4c9839dc50ae2303069e4fa0d7114a3780d722afa2a495c60ba64691c858b26d004aca6027b1a47d2fe0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a4f55937d623feb41720a7c1bd7218a1ef59ef0b5791ae63a233de8479571ecd4db762a16f7c6c7679ea457100da463b7aefb572a4b2519114ac43151503e345dcaea94e7b7f9a8154b2b622dba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5460d351d98661baa3cf0c2c7b818b24c2dc7ad0e8003b05fa3605921dec161add9faa53bcbafac39a519df0d11c08bbd34267a0d892732a552f2246d61933dbe9b9e2832b0d7e90813c281c416b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a1cfb5cafb30044390c5bb8e64fe6d69d18e6610b3971132b6d6b440ce4f84a3b7f15f4bb222143e4c7e5c650f313252182e8c4230bc8e5abb4736810e0d83fbbf91f4dfe65e52ab81f6d1f7cb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h357f80c3d5e726735e8e15f78ce7c9badee122a944b2336eb1b416dc0813625bafbeec70d84687dc2be502b5c22ead49c84a5be2789ab23e4875d758e60d31631a07455032f111e0cea690038077;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4753c700518a59780e226308956b8eef4d03506e37d470245d2864f05e8a376354df0d94ee0e574b48ad3fb910fc2026fb202f756abdee45e44525f16db4cb727d77005b47f33ed58ccf6f634b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85b9ce429420cade5c69208d3f2fd8c6ea4737bd0849a31a22a7a4fc9487bb4ae204641543989da2162b2521770743e280a0783cc46c6818c18a5ba8e5c5de10579f6d2d4282c741b59955152d4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a98bc2c186e2158672a6366dbefb66b8d54d0a10019eefb622340fd588ae497c8bc82900093fa05b05ae48d7dc26a952238b84053c379d07088fd33d5e283a0b8b540eca24055128c23aeea5892;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he04d77e67135fbe22887466ca6c2973358ea68ea90c4cfe5e99c70143c2846a292eea18081a02dc6896500ac88e92c3f3c04f75390d4c0415968f1cab919e8b55917098e21645b7786b0e8b71c11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81fe9f1ab723de1193a3c9e2f81c536b93e059343f48e771fb8a382f49d5cfd53452637993ac5a242be6573344cad50da85f8dd650a6cc350061fdab299e1ef813fe552258ea4d957af16c1c229f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8b926822148ed21bda3ea40d7248ca25f82731e49d59b23a3987af55345a772b6e68fc45c6e3913c85a80ef9d59df2e57c5cb7192f337ed64e69f6a4429cdf5c33e365e5a78802239b1813f5ef5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcf5e732273f33620dda7bd411dc855fd32239945d8539deed4ce816424c798ca95a7b0240f728b599c92d04a54130a82f17df5e5a3b3831c78e64276633483e0f0a7f986b2225741def6eea0cf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4db30432f80613ee175046117778ce43f0411fe58408d6d70ff912f7efba7514c91aed202db9cc1212353809d063d9189e1f5ef832b1f38ddffc87cb386c21613066de995843282eed19e5f3dae4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e73dba70eaaa94c185914566b8df3a622f02c5b0db8608b5e0f7baeae559fcec80410329e7d723d1811965bdcc164348329cfa1784b4c332438955661e180af3af060b041aa2a4ac43ee0cae11d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd43e0fbee42e92330025e38ca4e38965f0b65025e6251d781a9fb49657f774509a24d8f5fe53a5494cfd6db67d46f8de16bea47410eb6e408abd8b99f5efab79c38e2697ba7ce435a0fd46b4bb92;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b1b2ac32561dda4ff0888acc3205fe28bc8f0486aab2834ef2180f571ad558f2b3cdd600c40770e5aacc9566c227ce9871c96b430e7b02f7e9dcc04aaabb920a47347829bf8e2579aed60016454;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1660f913470110a4d423812c5c23b6c7aeb3b80b3c039a0a71af8b6f3d1dab39c83001a8d8f2b103d57d746975e4c99c55fe44131fe8163d2c69118346c432c5eadc1823ee31940f883486b05e7fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e86e7b0361ee82d138ac0e03f660a80808fbc45844e61250a225d4187bda54222bb0ead942cd8363577d599c5b331d5f8a1ea9466bae41748c41b9796d355a5d82565ea9db352764dd2266fd032;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he23db37638d2257f809150893c0efd39c69e24c1bd8785e34ce82d4620109bb733d997aa5bdc87efce306f9d45b3f4159efe176122452bb92b0be43187ca3c5ffdb625bc48febaf8e13f13f86661;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e0b6a5f41cd9d9e59345d8045369258780c2de3f40aafedca65ad4da7b3a3fc117b645b2746ca74fb75f1d7eb1f8a181be726aaa0f37616250658bf97c316318faf46cd794b6483e16461198dda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a71b362e212df2f5f4dfc5de9be79c1f17b3fa06bfdcd40e2a27a76923f7302026a3f449c12b33cb33ee9b8faa9b6a6d11abb3fe00a484ce9240e80a0d22934d34a09827f8119c6ba7e3f07a15f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9229f6377c8885e12d39027109b0544f4de839a2dc43034dc0ffdd9c0158b5d83cbb6722707d02cac8c846d99c0fdf92fbdfd6d3e8fdf5589d2aa859cfb6e6160488bf71a2a867edc8a8e6cbb00;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193b103e2faf4b9b8f8e8c7bae9625e0f819aa26992f0ad14cc2ee260bfdb6eb6683ee459c6b11401b88dd43150eecf36caac7a795aef2db66a18fb951fc9d4212448284bb07f5eb2aed825f1f830;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94301621c4763a1b3244769abec171f52f64017066c832269993119fbf9b082f4b3385d0e4777bb8b534c76bcf359745039310648ab5e53e08ee4d376695d0b7567a7774beafb47baf66a92c0249;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c82f858470dece24d1cc5b6434419bf4d50e4fc9f87c644edc3568560ca3c2df4982e293ab2f2c6a37b39065bde03a98b43c4fc0183be232d14a639d9a1f1a4cf086ba853ef5b0694b68fac1430d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec57301307ab4bd5efc6a16164303a5a5a78a6d003728cc0eae458bb0f153f602e381b8268afac43f81c9c0b411764ef897068294695db03920425b143d1714c51a9ff6f15a56941e03d3ec33341;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ffb910c27a21df1174324d27057d55e64b6514ab4b4edf466efa4c5ee5b96a41d5e8911e1621b75be9b329ec7a1902efee4d80f6bfa258d8495d0c18d1bd78875bdf3057b79ae63830220437bf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72513a61354fb9ec5a46a42d1574ccc14cd7a4892188fbabe23398ac3e4db0dffcb8a6a4be401fb3b26f06ec2f74083ce832bf17d7e0395028e63ec8d4b9caab5e5459157f042532918f6c33ad29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26d9cc5f56713d07816366279c5323ecbc449394d6b3932327c7cc81e89ccaba06bd27bfdba82b6ca8b3bb24579d393eb080a6100c28b6183d670ae14ce7f6b191e353eb418398c28448cf980114;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf01142b93ed10d063f4fb537a748f0f9ad2bf450cec490ba861913ad3daa163695759525730ebf6d417d514203092423f5cd8e8df5cdd75351118922fb5c9b7ecbbb0c607a5c4e01eee03f1e048;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3e79cadb3bdf3a2e7f02653429a593cb88a5670b16f54d8b43147e591b6f82c6d966b4ed83a528e370d123793d21e0a8d254807aa89a7fa3f33fe57a2c4cc070a70f1ea7f0fb9732555d5674026;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4cc0106b8d5bf47a0f50992420a33ec97d10121af91a451434503a02c4776ae2cb2c81e7a921a385eb3953fd7184f79365a6ff796715162146739868ee70f31e64a0463f70e429719c35e79445e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3673ce059e38074ff8ad884894389c2e91af9c4e15d67e302b4d9ef637f6478d989f8072b9179dbe60f9dd1e75062045ba85e3f39857b7a7b0e6f97307f9906c1cc77a044ee7ffc6ec809f3cedd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3190868e9be08a3e4ad34b97738c1cdc19619cff9e06f3bd8eaa25f5f2c1706db712f0c370a0778cf0b7ed779b773d5eb6f159bd4a84144cd4938d431e033655c6f22fc4547a03767a3b18277117;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h208072ed6ab030302c1e054798af8e72960090263029b4a651090bc19d2f5a129f695bae7f3732f103e07da7e4939cc83195b283e7c5cda1fac6eb7b57b54d4c8dc3c0047f978ff7494b396e4e5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59d03973f84673b92da2d8503cbbb78f81cf4864d9d99e51841e74e253004a07e0eb869094293e15c04a6fac461c73deb9996dbbd508ebfd0f4663691afa0231d3807d7a999de5c097c6b03fdac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7e640e1cb437d0ca388587d4c4486242657c57c649be43fef17b39afe35bd17a0d0de7f2c7b39642551ca33e58687c6f339efb644d4aca0d2ffacd148ae51af0ce642b884da0d35f346368e6c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64d7a1b6f318c9f4f246914e007c0a99255034544028e09a677c53dfa51fa911d876864995deabe86a48dc8ef598f02ca797fdac89b88009f69ccb3f6a22d940f1550fb2e432287520d1afcdbca1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1542458bb653bb354a64346d45df190416ddfe6023bd1618a5986ca6df4558303d1e5642b5b5cadf8fe037041d064f95d60ae7539927fc2f0875b8626155e4f816c8313892ad30e85b016d7219f09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca7ce61c175ea697a76d72b18c54bac0bcaca5182aa843e83f7d3db8f2746ae7f98e1505af24e42b95e634ba579358d5153945b23aea8412103b28404bb789ea2a99c166428d3acd23c6012dffd9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef33fbdc876b15dcf1aee2cd43ee0234952966eca8174aa652765049523cbe183a3ce728ff8ac58f02d6bd7bf968f038a4921b80b8e23190b4dc6e3df664f1f95e438bcec61d475e2fd9fce9314a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bdf0d2a0b674cf1b6028f7708621664b1a7e95cc2b32fef764d192daea51d4439cf1fc6e32b56afb77478e1af00657786453cb2b237a181a0db63da4e8f784c6826050abc1eb1f2cbca380132ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16bac8299776dae3df63097ebfa48da039a47578e5a8d4f550d159fd83ccb9a1c8f20641b7ffdf094fc0e40ec818c4148e61ccec1577e83373fefd4a8d7629a81e7f8e96c13edec2afb084f5885a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ba209cb63930db2c5a2f2fca55df4fde75c4dcbfbfe75133b68bf138286ff52c290fa29ad87d7c8e9b9ffe102bd708da417ee2ac69fdcca92db940e37e04bf3ae08296fbec8d35cc0b30cf5689f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed4eb210f1d247a16315d9962e727866a13e86006126091df8495f245c38ccbb8dbac792c44cf6e3ae94c1d2ae65288aeaaa9740cb327fba505a8f776935561f2213e861223298791b8ae51e0c18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2aea48875b1d986339b07c2a47296b2c52206a45f38f85c2fbec318864b67362ef0391dc7a337aa60304665cbaf7a735c4ad6f7dce869edab08e92c24d863669bfe096edc5ca4a73830a2eb3ef7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8d9677aca515193bd1143727cca22db96d307e02450aabd2c2b655a24fb0faa7cf00d6c26cad45d438f5a4382f9210c31f6d65fbb56171256009a4911f3b7f72757245eef0de5e0ab6281aa9b2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167c595b27bdb3f904b576793e38011119ee15217fe8a1efb13880b8e822aa5894a80391e4e85bd7f9511e302a88ac4e52fde2b5b319df74b48b4b75cd43d469666daa6db8be786d3696b85872354;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1475206c1d95159bd592ead7fc0d0fa37b0ab8a448b7689af5a05ffea355acc7e4697acecb492cce85069cce3615d710a178afaf92ce8748df2a2f886b6c58480108294d4aee84b9a24c2625d88c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3e3d5fef7f5f7baacf32f9634f71246a3fb599866ad2252b46f3bbd79a8091b91d8fd615476cb851a8013cf7dc02315785bf6effc8402972021c5ecbaafcc8392a14a9e9986559ba244d8f23128;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9de1767eba37f188e8ce964602c04898ec10b8e114288b24554173d88711318d2ff6d39fa5689c5a4bf6d5d94bd0695709eb9c28b3365334d3515ae6350817499b0663d3e1cf3cf57c7467472b74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1316cf1f391b53c5e66933e206ac2dea55775423ccbc76a1aef1f65d3e0e467a7ebbb63b505a2188037d7465e4360a5a9d57fdae148ffd85207973ede17994479f19c1c2027fff7c0fd3236deb5bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d57487162f08d40ee7b8e360ef5a2a3135b6fb6a58ba9a15db3d52975797a56bda0ec6e2f1774291eaa1c095fd0c8ced92e8ed2de4f794f8bda2b0595de40666e6e5fbeb3c0db76ef51ab90ed8ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173460c922d7dde9370e9ca59f72f9be8a684cedc939a56e72df4b7f8724a939936862207096c756d1489d1b8e278c9cc909ab9c7be6f575302a4af5abba748010231594eb7cb97afdbcfba923b75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9f31c27eec45d78685950b3acce7e3c6d3e98d3300965715162eff833db201fc7eeea92c890eedb2f49f19350537379aa4c050224b8ef7de6367f65384eace0aabc0d01dc8f152cd8c6b492c2e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14279296c80777dbc7748dc8f485f438520ae344cfb2e2e7b6f7389bde7bfe19f541302f87a11d86ac1493b3175025c6559dd6a7c0982bc629e16dfcc7fff33b0fa0ad4f06cb876ae19f213f3040b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10639fa637679e27bffccfaf2b0a3b881eb18db1500483900646b82f6235a00fb9b083bc925ae7db6b5b10a8137f8a5f8ee49091402531ede6fed2412151068b2955a47c5ee4fa35682bf03c7797b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178bdd1e2cfe43852bef69d94b3b00c5bd46a3b3e5442b93a8072e53cbce097cb697ad73e5e0740dc2f4393f1080d1a246a43800cc2c0912dfecf7993eee67ebf92e58544505e3681cdc5a776a330;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfee16ef0532fcdef9ea5bc173961a2026ea6c514d8ca5080c8c4e412868da20b07f8104a403c2d44f7494db912db1e0c9843623c6f8e2eeaea1ba34cb5e54aef6ff0102c24404dbda120fe339b11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8afb6533a3b6607bca50530a3e99e32e1ca97b8eb7e7aa6f320bb4e0cd89ca32e7fdac8b30d82b0ccf5f28b48531ffb6de7b45b5232179740dbd76366b9ac0f982bed9459c1b0ab8ee5b6bc2289;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9066bc7342e648ca1b97599d2e9a1ebe06f62301b315bdd3c32219ff9717806ac4553307af4ed83af588bdfc48ba0f6305218c1ad36d1e6ce134fc76e9357a5313ba57547afd9a88a9f7d45d1a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5424358aced233165abf13474de62496671c87c871fc59154574cce7444759910b2f358a6454c7bc3a57b7697ff1ba97aef75b3e64f407133efc5fe00ef0ad2cf31480b15ade38d0ad0efdbc16eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf90583571c313eb7bdf9ec9b1f7718262762001b13bbd412bc15bfc69c92ef02644e3ee4649008fcba9fd2564d78fd8fce38859cef8b73e024e75cfffab97a6b3e49476eed3bdab674c2c99a8955;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c3db4de502df1cce5bb2680926cfcf304f94b057c917b384ff38279f7f91954faac3e856ca8a37384cadf0dae29cd4268727370c4ab1e41dcf676e557a16ed57fa7ed4165a9d62045e48c126c3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13fac30ac806c537ecaa878948b19be3976f8af673457a32a34691960842b28e3840909feabec2a90b22b3aa6fba7fa919b054ada3a6a9dccd90c87a3cef56235ecc8a0300347d6b497250ded2f60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1219270be2a9aaadfa623c072771753377d2c0488ae2983d47b14c6b319711e4f39f87456e431711602ba8ca25c69547ff47280c5f240ebd85f7ac21346ce8b240f692b16a30b7b8d7ccb4d1c3cb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f40f29680b23449f659dbd4a63082e04952b420b70b8799ffc6e664f1b8fa5776afdc2ec0fc374ab5d2a91035d5a1195bfc59717b446fbf6ee3cb5156298ece93393773a30b07d54b478374e0f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6ff754c4c8ef2b65d9c7b98fccc7e3f6448f175d62bdbeab68a7141293c4d507ce65cf570a222d300d2d36039084294d045c84dcab38d44176ade0dfc68b02910743958bf4275b6e9caf11e36a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f4bbbbcebe47233a0cd006e187088e7d2355c51716eca946dd9d70ee54310b82186940e599612b16436980980286b098ce4b644140c3879aa0a88b03085c4e9fb77cbd02440aea17858ff2071;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb617b3b6c5cbfdc8d138ebe382ad265869804cfabdff61f5079184c6a3ed47388473229d786543cd868225b2ea9285b5286a8d8269f1b1b1db1098ed531af2a22b37321ab66407c2e7803a94a330;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce26349da014405045d5e7f41a1af8ac510c3b411c2916b251b0937e2a501bb32ba7d72c62f63d4a2b88a26389d9ebc317fa17d1cb92250b7e8a85ba3de10c06af87379f8582ed7355889118c093;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38db207d78da94749786d3dcf3933987f90c18302c3f2cb6f48e6d224cb2f86575110036972f3b06461000ac795c22729d4d9d53f999ea4049251bd61abeb946609e43697b38113e1708ed4234f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ca8816de85474b5f9286a7af803b1d925f913d2644a6c3dac4fce45853d8f2a4e204f0b7c5aeb9f59602754a4bf5acb5ef3d16e5a94269a1fd224de2a309d02baefb5bea797d1633cc3f3e64cb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7b600f8120a51ceac2df6bcfe08be22bf9721a6f09ec59b9f64dbdc3cf20176dbef32f8674712d293bebd981f0e55d80faecc6e3042da1a4f4c42631006640a8206d0068b5607ba5fc115c2dc5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c37c02879a794d7b714e59141a913ec2e5835a1428e55a480c5e46b7f6eb907c10d4af1efe07f5c54f1b4387d900335e6ea5ad3d0daa1fc3e5534f59c50999531de23c9530b90a5ffc57a663ccb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h233aee6c3de2753fa8b594d8ac03669590f95df194f1895d9fc0657403976acc668db15dea86b40ce55e4a17837b71eef4764e9e362257760316b0ff00bbbf06c4e720be52cf4c94725f6ee01179;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd8038acfff795564ccff20be830889b13d171924fbffa4d330cf1b4e6d26d572702533eb99aa330b493f2d2591554947a8615817308953ff2bbf1d1d942c08a17f741b52afed7eaa89d2e9e3190;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc731a90228b900ca011a61202c41414326336938ca19f6ce4be42599a469a4e2d6a8004cd08ad3c545d9d3bfd1475953b49adbf11e40f6cb672721eccc93605b174003f8e7e92bd67eec1249e27;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ac12cafffd4ecca2711099cb229b02cb553897a02091c20c4bd099e410cd3899542aaafdafd2cafb4879a4a030bd57eb3685a78aa31c44c08266584c600711f64c58c6873d303bb1f8ee06df6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da75bb679d1fbe6220f79149f6daa6ab9c206d13000bb4e7b662c39af7047b7ff0bba95ef107c88b5af59b35b16962e3545baefc8cd8c71ef9930b4458a4657c1450c56535db47a5dca07cbcf24e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h329372b1e6bf0bc406dc8350e9cf60fc0e769f23b908a1050a7248fe273e5f32564d8372c5e893574d45f0081fbd32e8b241aa2913af06fc40c19f4c16b0346fafef4f427a6e27ec92913a37555;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b78a23e32d52619592e434cca5817871ffb01ab410e228c94664e2eb6c0ef53952145b0c8ecae095143740bb26c808d8b9872b26c76bb87bb8ba5fdd897fc7d58b3848c1ede1687811abc0add2bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fca19a94d030d5ca0f727794cb079126006e1547ae45ed910e4ca4c98d3e9888bc625b33e55bb988fe310e4cdfab48fe0be75e3ff0f695523346255f4c37e70dd2020870851239e6ae475e1e673;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167b22a32b74e6e16722fb16fa40fa5fafc12c106b7221ea0502ad69d00b7b842672bd51ef3e9a0e4b3550d289e462c771056a604f2628bff260178a5cd487f7a67f95560ff64b17f93d26dea2ba1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0b6a843b960966f3a255f0c5148ce929b029c0e6d706f379341d6e66f999a49d4c557cc6f42dc7da70aeccdb01892c5a827d5d8b751068eed4f670eee42c36e276ce9a821c5032ffa055fbd8ca6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121f6ced9bafa215b30ebcece91a6a281f16cacb18a13eeb7e24c616c912ca15894c7ffc15fb3f60b6833d4ed46dd6257a4777e2937f2f1b8ea5987a894f4cc93276f6dccddb3077decd27cfe7973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12604687a0d7fa5a1db1f71b737f59df8ac05a9c084de32d0a96b89c94e390ad2346964583af68003510ac6bb9dddf282d6957641273fbaa08a6da794bfbb4cc4cb8d9f218d4a20faac025f0eb0ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c9f7c02b9054a68da0bf05d06c7e83a33b7c530fc79ff09420930922bf1b6c2fa995e4477eaa8d68d531048707ef269773f24bc8180b0f4ba69f36c73cc61da687f4c39ae61d4b4293e60f61acc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1866f21f858db29a9c7ac5c4fb858c050689132e02b968217898959e30867d8c51ab6e4b48d612a23c7b4aa3e39eae6515d5b264238a0a50803f4ed2ae74b602b8ca4317ff4f183d5cb11a85d94ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a8f48895d159d1fdccabb579c6b16fc77d98b573f9b742196ebaed4a9ff36ab9b9a74449f54f659ec631412d4766076386663c193f096eb01c7ec2026dad584c8c1e0fbce036c0610c975a985d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca8310d1f55ff53962ac4d84d494a0f44e4ec6e8ce3982758ee8027ae40ce18f025b2d2d2f6330dc3d0de102db2df06ce53ddad515e65c2c11e15fdee360db0fb21f7ea1599cf11c6fb7f7e7b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ffb7eab30445c2531ea41f81266458058fc8461499b3727d5fab509063697cea8c7b9b358402c26eb5a36c07e7ef6091a6e1b1d8f3d0727473a087fcc813007bea01cc323dd5cf39c4e00d3dc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d012fe65585f3fce14509fc0bdbb2584b12842ecfc8c28fb87a61a69dd37f41714584e866ea726d1e354b92f5827d4d52bcdb0b24a249af0ee7a82883da043539c6433198070a3654f22e5a3da6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde698ab9fec78de41400fbad48270fcf5738411d981ba5bef1d34c429d0aeba7200e794cf69b054006fb7cf0a39a35bced090ba70dbee03afc7d4396ec495bcb394e62eb28221bdde049d08c66c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70fb39b2b48234114113d86ddd3b1dd8e7295fa57262e6bcc5cfee0642394a7016326f37f49a861bbe54b32696f907917920bc86c94149e06ae33e48477e7c56d5b9f020db8366926df74c38b9bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d996bea41a010a6b56525f7fa06d870697a5e36a7373ba9a0faedb5ef35ed95094a46c2b0a6f7a7fc68cfba3402a378b1c1f8726175ba2306b6d9291feece6f00452461db104d2a8ccb424cc1e29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10198643f80f0c4238584f7786c133d19faaeb4e1356a54fa937d7006a8bfa9e7834fd0e59d2b4715eaa9dce2a44b3ff8d7c1639d1a8fb185a368731b3be71c4ddc1ee206e2b17d25d9ead029cc9f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacc2805958420843337044243e7297180cb04d38187eb4d276700042f9bc9248c77ef8681444a6206a76338c33d78de3988b8c9e81aa5ae4917b1bae5fba33a891fcf2a398732db515d04226deee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef314897d0afed6ca1d31f1bf48cce67c6cddb981843da025e0df591cff92fcca4640f6fd09a185f13c66ee5057cbf6310d2e3450ce31b147e19a39b3bb0bd15d56a83f1131db4d6b6ce07e84ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1460b523f79ba3e294cfea3942719d33af7c030cafc445e1977f80bcba4057d980bfc5c6e5b8902496fa943e98fdf08b418e39774f50e6afeb8ee09f76e6dae3c73273ea24b0d92df4d06be1a6f80;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106f03dc0998336163bcb1f2ac8ca437b4bf6a8d391b14cdb9f3cf366e9ef5113b86d07ca2b77607302a2dadf58c9ee45b58eeeee7d9eddb3e7f0b0dddc2c0da84c145eeed1ab2e4e58ede9427561;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d264ea849bcb630c8e072dd3e8fbcec37d282e7d17cc885e76edaa05eb476eb796c670eee8be2a40de49286d9bdb03d7f34444916ff00282beac7c16d68b570616eb7e76d52b4ff364ff6e54ba5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50348bbffb3800110e23d80c37bf69c66fecb800860d7421a212a018ae16e7049c2a868ad2bc4a8d0f378ec48cec979525c150a9322c1d9853a6ac8a8b3620a33908e6005edd337f212d266096be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h398d003d03afecdae25b8cdec18de760bb6a5df96bd06328555209c0f8d15dcbe97006337deabe8961ca3542036dc8fa133754ea2b9afc5f46168e6d8ef33ef5c1e0643d74e695912dc06f9b5961;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45b2ecc4468e9eec06d6f6f1dbd7e7fecf06f012b119466ec731c3192924726b52ddc07343bbdf4de25e05e2469f346f1409b4ba9b9162ca7d8a42ab766d971a24523f7cb4b1134811bed22356bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h275ac053a1381d6e2f3459616b6da71350346bc48ed2a3525f5bf9867572333c646e519774aa732dd9e0ac1f9f097d8b1317837c12c1c41871abfdaf7cc1f5e11326c5a51f9f00e29c1c27f250a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5856e4efc976dc728b7579d45e8f9d877736f58aabc763a11d175ee2d7d3d9f845347969b3841d668537b1b92fdf593c955c3956a6a0ec62b647781c4ac249cde3b51fd3b60d5ec0ee55106a8c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea951306ab26ea11fade9b5b860ad02bcbcc4ae8ab7eb23112f2efedac300233fa06037c7940598d84b1548721247ebb72bc5e51b8193968acef683889e8f0fde7de3df6d0a2e7ea21c69fc317c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96cba1badd02861a7b21b3802e178d30a89f72f0957fe3e04a257b3bf61270ebc06610225614965c7648804236aae05422175b06c5a108a46f5886b5eb8b58d8740a296139e755bd1ad4e38e6a07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17598a0437e9525652012066ff3a5cab76fd8ce597b3ea5c69e0c9ab0fd5e3441387a2135f65cabdf31e998fea9a20dcea338154cfe1fb44aa8c6936b39c90d8ee9acfb3a760b70d1a347112048a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13711d24a8f7f05918f076172e54d69e744982ab300721596b9ae0484c34923cf21ca3e164cba2dc60da8e91f0a6ed20bbe3a48c249aa6ca6c1fb38607750ac2731cee3b9ba6433af0d879f0e05b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118dc4397d5d08905665f495483740ffbedfa1c3208c4eae8bccbcda66fddb6e0b52eaa617f0693a8e3c0dacdba9455ba9cfece3880376d137b4604191d356d00b331383761d955fb0d276e6fd5c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115ca70491067c5742f6ead80ae69244ab9385cdb635c16a197aca78c515bb898c700717ac8745b84470fe86856c6fbc674afa1cdcefecf88cbc819e073561567f2ee4534bcc032eeab9f57934ed4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1abeb18b0f09f671b9eafd44dad78c95363294690894244b6f431945ac5568028d1d07fa4a9191bc157d45118d435099f126740fece9175e6d497272ec337ab6de0f3a71ec4ec29e720f99afb6a70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6b14ffc1f684085ac40473c5cad563ab128ebf3a5f14f5172c1e72388f307c2500368dbb0d2f8ad4c5597982fb706b8cfbdc7cbbf29431c84bd81b7eb1de9d9047973476406531df89c220bdfd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c639c57fd98e173f13165d42618a93805b96d948df39a1f5e8aa89586844068f0676fd4fcf3518f625c87215c9c91a6a656e155519833a6c0ff5a16dddb9a41571ce495a1a5c199e051f5d923fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ce6fdf14705d87ba558786ca0f779e968c607508059ada8032f0c4cc0069c7a156108b3704e5ac60ce7996271bceceaa182327aa041240d56574ff843b3456901c1cee263095d787540d738f70a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf5650bab3e81f85962928416a04d384dbf630a0eb9391009b0383f2b7b8ffa31c5b45a3159f428d47e500530cf56f0cd496e50fb2049fbf5cf77e532c5e8f8340bb300d9b5a0703bf2e74af38f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad41ad72e92ee35797003bf182ec5746cb7aadd863431f0e600131b2b3d7c9f3e53f12cdc4f9a580fc09bc975d28d33233f69566c62918722dc4468e59e90e15f6f545e1d64207a7c14c0cc6055a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1359344e9bf5ad72088cb0b7b4a0fd400959e548cd1c3682f33188b97739b82f679acbd371b3da4cf0e18a0f32b01738406107ea835d8316bcbdf7045fb287c0e5a577d7e06e681de72d29bd9a9fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf32dcde2d5ca9aac612d1507584d8b82c342556cecd710241f8b195a433be3b8cef07a342c1329e9eb58b052a736ddd8909c50bc1ea21cc79fc7ca6e8ab247b87ef56dc2c91437e527b4c817e9d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b50d6370e054f5dcb7178f69477152d6005f56684f509ed911592400449f681a06a05a84edb062c5fb2624a802ee255ac43d14f379c15fa8e3f094b2f079bb0cc55188be2f0e7fb369d5f85d5a82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d4708474c7b8ba364815737004719a97f9b4c1b23d20d5afaeb267618f80ef2cf6110661786af5d5e972b39bda942bbbbc67df3bcd6d04a779641882e76cd502d3bdf9d74106d74bbfb1c854610;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c07c785efe3546eba8c13bb4f5926d575cfa0bee6156babd0730449a65ab431b414f7d18aab3f59660cfa33d6f5ddcc0a9c66af7dbb381afe62eab6503f3b0bbe8ae798db318ffd96b56d0b99251;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2687174f130eacd36810b538d471808277c395bcae99948cf0b1c5d636fcbb1ce8cb51610cb2f639aeb4a536abbe16db602ac0c16686cc7fc3d494c706b6860b3e873e64e91cbec79dbb951a8b41;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121a14014c8c29786fb00f3765987109d3bb46576e8b8e547719d74245d6143752ef18968232cbf2aeeb89ae346c2c254f45ea1e0cf8a4e496af1fef8b5bfd4dbceb27ca666d53ff5edd290473136;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha184663c47ad909671cab2401f43b0f71daa359c6861d49cdeb42f35f1af269abdb85bd17e00de0c2ad4dc0777e53fbb2bbe9dcbcec3a42cc7848cf752e8d644213d2e14e2dcd10f07062321538;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196b5af5bf310cabedd9fbc9f35d79db2edc6979813a34d7743aed0646965976fd753dd6cd1489c851bb0cfef0f3a53e349b7612daa988ca0c4ccf98367b251fe8c489a5dbf5c94b307daba50c1bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c62a4fe0fa260e6b030e499f252bdf13ee0511b33147cbe29e8995eae586a58a0d45a9ea6f802f9a4a7e4605fe3cbb4dfa3d88f073936e534be450d25d3ee0c1280b058b674f10c453fe4b0fe19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11367b18ce5c4e5c883482138150403532ffb2c22dc50d9e1ea117001fa3dcd9336ac035b89a40290e0a251407ff3b003f1256ce7b9d8b2fba03ec55f1a1b527907b49a4f10ba87bd158dc4e83776;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127d63449d947ae32e985b8efbb933dd558bb83605674ab2d5c197e9b5ddd35e1f275468fe58cc9edb84fb8f0db404b8f12c2ae509d44defa7c507ada6d1901da1c5c2afd2f892313b13836a882c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2874b0303ffe6b7277c56edfbf03973c1255cf1c8f7f5290f0231b19c2d61cb8ad19034497d4374f78c841686a6e090af43be493f29bd233cafb6435c07fd6b58c7c47280df8d642380ef4cee23c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1564bab6c5a908d6a4f8334fd2397300a46c72bd5153023ef7c0cd3fa1e5ab1d88d5052eacf624e28620e4bae83d3dae77ab2641f32e006417d8efa4db7feac7dda7c191b24d236d1d8f01b34bc84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2b048475b41e6a4ca703e65d63d2f1ca3801fdc7463cb0c27f0d79cfdb289930070a01c47058023719b08c47aa18dec6f807087cfe7263b302cd337750151aab0d2aee4390a40c8fde9b9310285;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h577bf6b6597b455a238a0d421aa368ec22300c0b7ab2f1ac2f097904e10e0993094419822a42c7a7eb8d063d0c9a94add3620a2dfb4ce13cb163d9ba1d9dd7230637add0f5e08fbbb5c7cef80883;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha009825985d85a8a10e99a5136dbae56b5096f695b7e35f029a5984c51c6a4bbeebc4f02c49b9cc2cde99706666810e69da94664b8d7b9a2151976014bab09839f439c33325468bb1e968185cbf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf1c401ea11b02c8ef0c0d6f5470ea594a28e43353b6482318f4d18459e990736c5331a1b84120740b672d2fcbeb04d3b63d18d0a4efb8862228b4e81e9bb8c9b18b46278f934db7c2eb79d03c568;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d794964e45f7ae872f91874c3b84e766dd4481f468d9b4eb53d206ef6eef1edaf435a484c9d52f065d62b703058338cda3705fbaf249d6dde3a0cc0eaec79a9c779e05712fea4849ce6728477097;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167790d9825c014775c7dfe473dd17c66ee6109c97ab7d6cfc8ac1cea6541b6497e392188808f938cef4f71c1a50c1c0ce7e20b4bdba8d9b2881a52690211595e7d36b950e884b3ef9b347181ec63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8686f8e7f639697cf8a0b58fc106a12394bc73e7759a6562a01c0961c0f8cbd2dcd57a5d9ee57c0245619e0d98b4647a634e452ee968ba13c73d7a01b24ab716637a15b7b1855e055647747fe2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134c91c26b63b842a44d4a70596658ae0cafe47e1ad3ff1436f2507a0e66607a5967e76c51fa810ec2dc74443e08a994c413f7a7bd7ffb16e7b9c8accbbff841e89f4e932fe84855caf6f0071e28c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134db24f94c6eb23e346f094f91d3ec21606f992ac27663efede5089aeb2b052cdb15e04ca93b3046b653b8d9f68024ecf53f19e7122c2d2b7e373b435ea4df2cc2da0793e4aad1f17d33e7ed69f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100d6a49c4290b66cb24486ce71ad7ce6e0f7eea8846d92cf73c9ac129f1db1a8c60b1a89b74e6da294e77ef7b4188d2e6641c9a2e279c26a53979bffd9e5bc1fb3c8de117f988770ae3e0675e101;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc54818f591548140bdadfd76e8c3167d2a3ff095203472aef2947904554ca879331bd7cb484d966345291416c89e4b7a8c042fb290dcd488cd368386eaad1cfb575c545cd5fb1ccc322035f99c1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fafd8c0297a3bf83c0c0cf5f020e6bdacf929f59dc409839eefc63d2a698bd5624c77f4b553fae3eb80c20cb31665c98f9fae1402fd3e97500bcb297d2908046e3d0fa652a25f96c77b440c55463;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6f44f89d95ca3ae5e8496dfd23af6fe8f84f582dbe9896cc790e90306eab8bbadc10b769ea386c4cf62e18d31338bd270d5817b3fc09ba5c2590b19dc5a67a3eaf47051d7a090fc2ffcfb9f27e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36dd01acdcb4958e1c5e09f0075d2bededeb696ee95783baa2d3442705764f78d595702757e67d4b800b91eb4e225d83d3f2dcc3201c549200a68c32f857e308d51e32276b1f13f387bfbfff2247;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h919c50409c7735126681cf36117d9dc485171d085c4355f456809bc07865c74fc196621a9185f76569cdb14ec2e8bd6b0997ad98951fe601e1ee3c3a27a4c7ea4077cb944f58210ef70f126eea0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3106e55f987f2037241f4ab17b00c696a0ee14bc097734deb9f66f026d19860a03a7f6369296e1d661550e0142c1b3310870d1e5fc03d6f8bee003aaac76d945de2833001fdd638df3a011e0077;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9be04a6421e66ef2a97541045525acdbafe55787bbf478091aba35a790c30fdacd352dc52728281be478f26bc6ee668020e56e2b141c02ac0119bfb4c1b399cd9bc7acfa4bc7865f8aa873d7ebd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd132f86844437a8cdb93bb520d8be18079743902248d6f566a12ed269ac2971f467fae2871172bb112291ae2a08a43549944eb4e47192cc83a03a59977beb3b209b9efd5f9a8b7c763cdc728dc8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7aa7eba95e8f9c60e794c2b2573aeccf85d5b750d27471ebb1ca1f2deff701f59e2c615b7a15b97ca9cd07f5a376dd4b95ede2c7622417a32897d109811fbdb894ee1ea278767ac666ba215dafd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1368a984a5e4f083a79d3b4ecbd9c2eb430af20e6972762378229ba02d01d49b5014c7bf0185db0ae1d1c21201ff70357c7a53b833b3383a3ee0c344fee540906dcfafbe6d687410ff377daea06b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fafccf2f05e4b527d3d7a0624908e00a6af813ef51aec8ba68c2251389a025c382c86330cf74368bf5e35cdb15e4df22741561aa494b0384deb15723b7d4a6788ff8325abdaecaa7cb7fc4539f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c81762bbc1c01d338c50b27e2c97d73c00099b3b06b13d339b5581ef2ab5f3cd9e02ff85a0a126c6d71c79abaf2f6361caf509946e680b0609572093779dc6d3b8bb9385527e49cfa5cca804892;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7f1a6510eb48feeb6b683decd5c8b3aa18d0399082e75afc6e2a130b145c949ed95f52683198a545c799c841fed0575645a4ce3b8a5e12693f4ac60339c187f9cf6c24e61deaafc558552c9cfd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2874e34671b1fd7fa942d517fa9384c7b0f1fbb41da0ab7e45fec1dde1173cfa8611197dcfa9a51deb2217473bbde299fba4b4b8c374d32549d88cf95be2515f9b5a201738a52ffe0392e003e2e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3cbc44e0de601188c75e8901f693714c8551b38b865f68398e2094bd15aa269bd475f43b66133f9844be184dcb0c9f766b6efeb852612734c2caf2007d171131a9a43957c1e5b76c91ab2a8a77f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3019143d497e6141c238dedde16c46ab43ab833908775159d54dbc86446d5e0bad7630f3f2a518130a694e8b367036bdff057e8d3c6b831f7268790bb90a2de5d11db564d6460122ccdebe3947c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130f973b8abaea96ac9b7728fc8b30d0e9c2e173d69a9afe07b36cdb526e41d7ed52dde1fdf37081d9df313b9a1c36e5a9de1663ed95821ba02209c94422fb67fb9c3df500462f8690d4d321eab65;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc84fa2e22ad310a7b7b03c09b7e3aed1f25fc82cb89f40c704cd6b17fec53acddb166b3bd4ec1dc67e0897354cc2f697057e81e54cd3d69004c18db30fa9a41d1f8b8953db489f038537e3e89e9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93a9f7a960b68a55947d0080a8036da930c0c5ef5f9f4821298f1de437c9fb45529f4f1ae3c9f571b29632711646cda089fb197ba229bbad6e0d358c2776dd698414dcebf570b488bb7a00ba6cc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dafe68b7d5c50907824adf96689bf96e629a70de532605e4ad15cd09d99f7856e8916a4f88ede2ba88bc29cfb64fce835bc2e49ca075a8b073ac455c4ae504055def180a026cfb433e7cacd37065;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b49d67e457ed8df24b0f869c5b0952f75ff2cc34d126cf87af139d0088b0b6aee4c9742a5f88db394a2d00576927c0869de377d61d807f498479c0ddc133bd3169e1e2b047a5af7a2681982490f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5aa4f66bc7e8505640f819f8d5d4b89b0eae22f74fa049bc87eced0581c225cf96e6a3b75c1b83836457da53094c68607ed2074e163417b66572143cc26151ac8a236dac5aefc19614ced3f37c75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9e68feb9769882702771e55a028ced4d5ebcd54eb8c7b65e317f0bfb09281033c02f09b86c1ddfbbedd787e549d43f39f709fab822bbce7e586581d6407f1cc752f88a836f5ca02510c1e19bcab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef801db4e7302591cee41c3a3d563df8f63eb23d438e2af62d014726187d1153b20410e33de78b328a0fbd079592ea58314600a5b92f2acca81d99458a93195c87bb6615541885da3b8f125025eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17130953ef408ccb06a9989453376e0bdcbee3516316b1d08081c75c6dc3df98a6599aab1a6aa44d600bbd6f74dd685ee0154ded02bb2a0d8686634c0bb3b86e7f35c09321887c0e3a30ed9d927fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd44212f7cb63407f319e690b6d256c12ba19c14e4d8ead5284071a23365c1f31201cd4b7ff69004a6dcc757982992b3bd6a57f1e7d05a227d12f4fc83fd2e11b98930f3a259ab16bae7340c01cda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec4f85570d8bc335e4b280c469eff8b700d14189dafa7de1d22977b43d174e6caa3ae4c828890579f8066a3ba10de30097649514cd0a7bc5bd652c7e2cefa560bbc8c238d4d3d6d336e148d59919;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccc7d4135c270d8776f93f69b7615095025efe36b2721f22d6b7f62cce90922170905711f09391b59a7451efa453ae1590cd11c422fc13eb7b72aabe48253cb4d741886a6aadaf77333196074f55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecdf4cc895dabfe1f3dc23dab19df407d456b19953e35f05450de5a08b21fed330e19f18e4ce1d419fa5167bbbda3171dcaa15b05b0ead304d23c3d4ccdde0497d1885960014a90439f0c6fcf84d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16288d7bb9da396e54f2035157eacb52ed810a8a1da4d9fb8ce582c884e1ec264d51275642c3a931a9464f0e39302dd0414a362bebe3cc0ebcbc5cf0f0c2741ac102697cda28fc0c7af03724a64e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1afd568f634b15d7a450adf872422558a2b81fab422c8b1d1aec6ca0bb3073ba15f474f991b9935c00811d0c65bba54af4d76c25aaac2239057eb1969570bb830c24096ce107009aae3b7f68f0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d822869a2cb378df82319b1ccf5327c0101eb1a934350e838e99222e285435339c10a79b785d27dcc4b8f1ec98748f8a56dea3b0a63078586c4e46e1413dbc8eae4096120fdb8e828f722f1ca03;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfafd5dc85d00afd38b1356815dba136302f7620fe4186b3b6ccdbdee762553d7aa7fdea30f3ff4fa08cc422db63b35330bd0dce1cffc55849b15bf64486246445637d6dac5535b7957ae15478ca7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h737c7f1d7d293643923ddd2490b7c5154be993c93f4a3045f2c42bf2c78ef0cc30261164a2ce32a031b40ff6daff241d11d6841ed720848279a50d5c3b43d28483479dc72711ab406dd83bd3842c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h431bc9cbe5d392ab5f7c3744ffe29180d009c065eae6a34ab5c72ea2e0e819e478caa1ab31a1b772a65e70abdb74fc9acc9ebe6973ec2aeca0ca92534cfd3965ab0ee23dcd9a2d3822a31f846758;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cacdede06c279664bd04c90c4e74e7798be92dbae0202e55f2d96811f464e943c932e4537632329e4db9a7679ec2ea3564a8c032f2839641b5e0daf264dcde81d817f0601f20115dd6c09f1143c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c89d7275c406935203b1f458ab1ccabadc3879809b84b2c13c9d50485db40f22d02f3a34775897a3355c2239e66ac85d5ae6d092f60d3b4e59613e61068c117b2d786baf52e7aa40cae125e16e38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd523b86d97be3279453391d1a040a431a6c47d4beb3635b455a352d3de8fa81a7af1de05fbe18aec0231781c6ef04f9a3717f299d2fd3758baa801ba70213886706ebcdbda54c55cefb69a26fea1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2b4005ee6b16002a4b507e2359468de914fa040fbdd2a476d4e40dbc744dbfbae9608a1d170692b2ad649d22a68991ee4f027b76e7c521175dd4398773616d0e85f0c0fcc8c21ebe66cac731f3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77f88f0a037732707dcb4b66511b9cda97eec6873311ac8014282e46c2fc398e2a97b0093f4589696a70f67702420db4ba1d9e005d0b7362606d6590a8bf6efc3edaaae7189c63cefa5b23ea0bed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e00752f47000b580c99720433d561eedf43534f5bee9783424e1f18c6225b68e9134d8349cbb2369dcd17a35a70f98cb19af5851fd64a8a496698bb6bffcf620a0e5ddb1654b94d33b9b98675a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5a319262efffafd38353c4b4aeef90048cb681d789daaca92f6fbcaedb2809592e5e178cbb2e1057eca296bdadb4929e93b8897e92db6161f178b2f759e642a85957c8ccbd1b46964d4cd3997b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7ece8439cb1352fa5a448244f5c3dde72c790213cc6f764ca097ca8f5b5fdc27878073f94ad6be108ba9ceeb5cf73757c8afd27de830ff5b84e14582bd9bea4628481dbe80861f6df3ef6b2bbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had1b5c5714f4bc64b439fd2615b031822135b2a2e8eb0e82a554e810474dea17c70659378ccd285bf43edf0248dee53243d99997c98399d41be6d2d034f3680fb31604cf4ec77d308e8f93dc7c83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a86c9c46f8585fdfd0f612f2bf6e4e9a6e822619f19b75a380da8cf9d785b4a11c365d06ed54a39804dcaed333b12d3f74c2a0072c39e759a549d2f4f2a83f71c10fd782c662234f6184e00234f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11636e6af28605ae60d2eead99485b1e1a01191cdbb0657cd4566733395e3297dfac8b4d01e6a4e21394c75b3dcfe08b74d529bf3bd9869207fa5533fd52a82f95c9421829ce5114f8bb78fa7e16d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b92a2dbc9f2257c1b680abadaa93693e3f1a9e8c0dd4de5a67658e1ee72439ecf98050105cfba6ef90b6c4ffb56b25b930a655b446fa5786e4ddd7d7f1ced6a4aaadc90e9481cb8331b00c14bb7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f378896848e4a65243abf4de3d9c077e8e2877be54e38f37c5475d28dad15778a3b6455978d696acd9e440ef3dc962e819f3e55f3b92843c5518a649ee392a484081459108cd7ead7f0f4cefd40f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e91c132932b2c6d71da6f427b96b9726aa43b30d4b66c1a155e690f3140fa99dca6b7280eee08561026c0e9a50efce13be24234f306d5852c06bd57061612e524ec317d49b4e5f2fc25931a40a2a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134d405bcb4c4717eedd9bd57686aabe9ddf72a06cd8706db6d10d87660e77a9d14203005b41d30d3bcb9af8775a92c1b58b8a058d1220ad6e98e252543348e70d57d5845ed1146370662462b524;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102eace6f80888d615fc6f8b363716e50336ec3be75402f917bf7a59ec2e1c7a9b3863701a9c1e3750e7d7ab619824345577b122cb0148d5e09a2ad5a8490205407f2445fccab727f06c5b2eab037;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60887aa8ac02437393048f4ddda11347330873030313f77f6047889e1e3baf97a2a49af0e72830e89bdf0a23d2d0506dc78cfb7d82fab4e75c200ab48b2afe9fb1432c10de2b67f25bd360993149;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h630280ea1bc3cfab6d7d3e3468387df90c44d7c9d71184f4374107f3af05ca0a86c1197b86d69e114eeeb3edbc2691bc7156f36500b305ed22c905434568b05e157e8204b1c7d57b0aa9a5c643f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16abd3d357c270ca3d24d03ca46167a04fccff3250352c336a89576d3a7c150e1e0380e29898b2a7139169b6b126406f165e4d4901e6b8f13c099656e70da94639d192a5d19c0f617d99338ba91f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f2ed3b8d80468a97190a1a21a709e851848d8d9c2ed2cd8f56352e658dac2a24351e03a6a923147ec80e1d7c1970979b7285f20acb6fc17ce082860dbfe90c93fc5a8369ca8ad8fb71c23d00ef5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1728e5611d529211035b820e01de965dc4f1f691b75bce79459d6bcc85a66e87085852a97a3bf9149434026a7ded3a11fffad39fa70cfc64a0ebbbac65bcadf248c06e76ac567374607f7645ea574;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h362744fa65ddad3558664267eee5f319f16a8851b6657623d1700cc7bb03d17c05574604670105892d4f18edc2c1ddd3411d58c4d95685365fed088495dbd834068d49a4f7080fad26304af436a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b6a423918895679feeaeb288ff2a4d8e777811d1a3f1a9d5234b9c0c6506c23a1405ad203af9575f0aa4b241470a8680508f6c23fa6fcf29fe4b4a09f26c841edbc6164ea570038714b568f5780;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b93335e4369654f61d77045e4908904ddfe37eade44b038ca7ec939d43692228f59e240eb5986b8c7516153c8e2cd3c0f7f1ea384809f62e649aa6b74848eedc1ed9ffef500ff892d99a0ea2d3fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31cd86bff04933a8d4764b85c80bc961ad83ffcd3672efb207aad8688c4b74e9572913c5200eb175c7940d61cbc67118943b1809fd0460a35e49cd40fec74496adaf21a76996297844ce9011c1d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140452263a2042daac24c8f4c34b0d164f0e50bdb69a1b6261c6e11a06a437adcf72dac7444780f7c4d7b42b13b80ce5dc6c3ba54ab1e5a49132c15ddb1e5ee12a59812c2ffc789dcc845fc8cf89b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44cf96d3df188b42ba73ee7764c41ba193b5ac162650b61de7c9423d5b5395ea156d54c094037a3c373b63b040cb2478e6de3fee4d296e589d73d31ceb0324a311ff604f8b853fd6f155f4684352;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17961cf93aebf40eb12b56830ce187d439ad3882ec41efb15060024c249209603ffa6de3111f5f0d3d2b6729773e52d6dd918c7b3962590f2bdc59de0d7ae51bbbdabd69f79bb3bcb92b550cdfd76;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b13b776a79b4cc546dabb0bc20b1d465a48407dc1f75e1698810e7e38e679cb11a5baf9b50bb74ae07496070af8e2a7828195160053137e5d2b359eaa1f9084ce8b34671291c53b867b8c243f92;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6ac56a1d66663d5d0817dfa0af9948975ac0356df42c8e77d32752eb673481049e6779e6639f4e341de43b32765041b8f982fafb2c45f49102a8790f1af9f921079ef8a3ca554304608c8544f31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9a835f2f78b0cf604ce2d0e78b7b241c996532220e47208d14b4679efdc8c21c319d83b25643fb690b7c0479316299a5a6eebc1e5aa744bafb82f262358b19a9cbd784486e15d0b884c7715ffd7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17401e8fd17904e3b30c6f8fdcb3305c34edca63357ab0219025ca9fbaa6d1bb6aca25e2aec00a9e565092dd75b73ca6f11adf8c8566782436a2d17f5a10b8081c9cde207d18fa07866be13309c15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9616b005005f1d754dc5a87f23a4fad2d2b67ddf3fb62a0970ba3f9ea64f40beedc2225c35df3d7cdfce7fc06d37c254fb7a571c315225c88a80647a612fa3b120fdae5c56d6f98fd9a6367cc6ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf11ed42cebad0bebe4bc17bf62800c76a278c1127e1f453ee496893073613c7ae84098fd3311337858ab488419bcd9dce91dea7a1686df1a4891ba860012318dd589cdc75f330f0193214780a38b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36325bb46da77cc697b9b125eead0269d96a450bb6086a4c6508c1bb84f9be594ba902b5265fbd5120fa6238fb30cc2dd8cade31f13c3aa86b4f5dddde9ade8f295c3d47084e4b61952d52a918c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fb727633f6909b974007d43f1877f51e51c845bc4a70ea0bb550c864e88af76dc7a866dadbd2224900c752365cdf2e0bf3b1a93133103aa9c98bff6891080880e379639e7348f9854b041aaf13b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfb40a79bf0125fdb9dca4f29c4a815dad3d982db319af9dd78c052e24f32a376dfb5f4a6673aec91fed3310fd5d73fb27a7808a2991985cdf4f85ad7813654146215d3b89335d76544656e69fef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83d451ae7bac0227e59bc821772e18ca75ac83b3fd297d7c0e0c7a941359bd14d929def3041384d272fe17328d9273941cc3fc1ef8a23fc41386146f0b42bc1bf9c408a95d506f4f2d52ee501761;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114d0df60090417485c2e7408ce49f384579a0b0aa64233baf2650e2db9d0ab835dfa5b79c28ae53198006fbfa4660895425bb7bc2008eca1bb4940b9afcd38eda7afb488d8edc456a2d1cbf5cbc4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7981711705b7971e73df769fb06f03d354b175743ac47c578eecb08448426080a62a11dbc34349f7e7d3421aef0a896e874f20d3058564e27bae27431e63a7ad44c1ad672e4d087c44da8f41799;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf744314d35185f6a1a5318c4998ed1a29b028d4618f3cae88f795d245c1964c9a77b0d418dba12874743e141d9745bc2294e97c274fe48de1505dd02c18f46b66bfdbd8ad42d706c5f27af5406c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e75d37bd53ce20e321b07a4886130835c1b54f6d82c8c76cccb5812ece927f3553415465b955f23c96f5c39177d3d18582556f357cfdb8cfe0562c7e8ca0dbbbbee7c946b8bb51c0b90a38093c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h989c1a3895a8446079c2e20197181a8b7e14d2bd66872b840b012cec3dfe5ab3eecc69f9d86cf5cbbe1a51ef0992fe2d9c4bedc90291a606e352b65c3e3c2275f6ae0888c7cff468ac6000ad97e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ccf5409f5e9a75e109ffff4cc4ba18b403541d8fb8aaf1644d275ed375528ea3ddc8b41ee411cec307c41c4d7c9a7ca12110339c0c507a25a03c7b0eaebd5dd74635ae0b8c2e282c062e0cdd13a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2305cec38dcd2e54e826dd37f58bc2f50e8d2b62ba6f25b6402845dc5b7d116cce985db85fee494035f9eb34df8ec385d147d2aea598ea1cc3fcba60a37770cd1d60b75b52c6d8952baf600cafc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12bef2f383f832333c8c0b0736baf39e2f956179f8536bb269a4ca2cd911b6230aed0223872b187a0040380f49e0f63e152e24511646eb11a5f3b43114d13740d3ef9e2131c7fbf9d0bd4e429d6ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2b1f1731d90137f1ac1e7b0a9c5697f4fce8ac8cf27efb9ea7a982ffb23339f11d4c4d84b3b58c4ba757be3d977973f076142e667ea940f6a110dce9981de8a2ebaf11864e0d868ca0e9ece1b62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9364966b835de5af0d34380ab05a5ba2e1d7d826f246ab5553cfe4971fe9459eab28c9a8cff69249bc660659a59ce9dc8bc163326878ab7b829c81f9762bd8a8ec7668dca99d2546ebc2b4133150;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h554c98253d1b98fc105fd8b5e29e5fa00c977fbb0d5dff0de34db8f51f40e7873de09f942dca8056274f8cf7ed448948dd4d71dd20347c90195dff37c1bcefeaa751a3c33b63628285acc83157d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cea9eda48d5681ba562482f85832460937ff803ebdaa0ac2c21ab81160e7fa1636c59713d85d1a6fd9d321265c923ce77f95ddfd545c99b25d2e3c0894e80abcc82017ae9425c0050ad9de5eaebd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h673e4e160f6ccfc57248f9620a50456f1fe339d18cdd33e87d14323fa8181d4976a93baad201f2c20691c5dc5f3e2fa5f5c72bf02692077e462525d1c181427922e14be8aa3cba72b098893a0e74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd54460aa1d3406fe1063f70c05f0e485457303cac506d5b38dac6d81cc398273d225fd25f21988fcb513eec44055392bade4e67e1299b431613077a164b38f4fd943b7a160f9ecec70dc63f0df1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16593cd1ac074ec2a619ff9d10c4c86396c6945c15fcb7e24455e78ca37d6b13b30d644bf76cc35fe34afa3b1e7469d9269488c363fcc186fd6b5d87f4aa54428fcf645f33ff7bfbdfd2a375f66f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb0726c1be1dbbf15dba276722304feb7961c438330243e3a37300d57c5febb497c1c2d40e132fa3e449fed91753f5fb272b92ee2245ad1b3614b68655dfcd4d679c74b053a24ebbd5f3e362a8f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bcbfaba43ed7c7ece1804c132186f7463517683ed1da2f33a64d9d8ac5b9cc7a783b160be1183758dcde7099a1af8a2a6f3e3f83601bdccc1f3917c5dee3e84906aeb26eba3398ac720895892a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h646aede590fe2b6c7628f2f408bd2fcfc15b7764d9da5d9511b79b426d1205dfa559bff0ba951d4f03db13460085206a4e870aa00798cd3296f6536691461b2da317ad65c0d0198da40320927ca8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1047c007f73feee04c5827dbb97cb06234c2300144ac432c69bb88b93513942e8b55e15a9ff7d8d5e6ed8397ac23292561eb9ed8e5aae00da66513aeb17c53d9e4e0eab13ed331ab74b28b502b4cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e9e45dd3de6a3f90f6ca76579be2b2d6e9171a148919179be2e17e6df98bdb6acc0c994fbb419616f383eb44ad97f7a36d2b003f152758b4aa86eb0ad22c133c22bdf1ea53d6b3143cc2b3a3fcd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c133c08ed7f0e6cd2c673b37ad95f22f37136f574d6ff1df59e78bf3687ee97b43f0ddc839a3656f71572ffc1f225604b9bcc8588610052ac25149cdef1e7043f88c9bff4da4274d788f1421fd48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc829c695254c5542f63bbebd4d21fffacad0fb7b3ddb9bc25c2280c10690df292a620d7bc18e5ea6195c23b617574eac1177fea75963d59908aed3b44cd3e07d4754b243f14f1df6aa339e5cc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e0a97504238e7237fa9856fd749e7e2fbbd4897c4d0eeab258a897486e84b6038f0c92a0c0c70fe3f40aa1d7272bb38b05a8c24de988224199955f40dabf27190953a0381008a2d6eb45f40e0cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he143b7c6006df84891a85bbbc41a23116e24406a1b5f5dec20c48feec5308d8e60249be2bd2657a1c0dee3f421417486f80e44d0bfa3fb5df796b6e90689c489c5bdcc96e8d36e643e7c03e58ca4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18783bc1069cf0615ce9c9766ed128f95c379dfe198fa3cd3a7acb0eb66cf53b1ec19db397d9ff1487956325688941d86b6d87baa02e19ff5075741e8e37f44694a9d5b0057c0e7b9f38a3fb76c00;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0eeb3f52e64d5c3e97a37ce2d2a06197fa39d1a4a1291d0ffb7e5a745d615a2c6a83691786ed849841822d1c180307fc12aff353799484cd2acd6cdbb4dbfa87b98807da712e76a7163f498712f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163729fa1932eee423e010df53f0b2aaee6fe62ea2b7d0b244bbab8465525f656afbc4bc673a1cc59dcc22ad59f1e81d81eb916d30e47d9d71d28a8b35f3cae654c4224e9d297a96fdf77e0da7603;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5ba3063f18d4f61f2a47e9bb0bb75dbb16bfb344b86e7b6212d3c0d4429e4070076f426b36501ff70b79f5a7811b68dce50000a5257eaadeecb47d778ee574b6bca09e7bc1cf25b5d6cee4d34cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1534994fe7102685d380c1a6b6492eec7b4cf3e77a07da5bc77021848df1b0e8fc958c64fbe44fdb8bf5977760e9fd0bf3a0a775bab1cf3fe1b0106c71e508f7a5fa8bd3b005a2ae1915c14f0ffa2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b5dffed5f11edea16b050be65beafe0d871f0d643035807526617e1d1f3c031ed1b5bff43c55e15643b845d934d4e0fad2b47ce1dafca5d8773060f9491afedc50e76b92a834ca906a283ea070f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8fbd5aa26709b4d5d590916ca4ecb8e5abb406dd681b8f51bec9807095b0a61c3b96fce3b38c2c135a7244739e069960e96c12dca426447c010e60699a06fefd0d2bd53d4ee07e5891d52bc99c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa03d18c2495e1d3d78838f296084e12f4cdb2c997893f33a378a0e9c3371ece6affc0a14dbaf2cfb3126a9169e07fa133351a5d9defcd9f8bbdc3ba69aad47ba9679f6940e92c5b29456fb9dab4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6e560584230bb12ba8a9494779d2a952e110a6fd08d555367c3a64b904794bc209af465d726df7af6ccd71c42e290521ab9b2ac644abe9e1d0bc86b0f78b33769ef77f71d03dde41df214eee392;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8169c5b257f392848a08e308889c1f34ac7e87f0e63ceb334ce47752f4ed7b48b85ebb1d3360daa960d5d825d4ca006438d581d10f286482039bbd79f27b1cec7129d338df0ee7d463914fa450e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1705e30f6cf2194debe8ea977c0fbf3724993821436a374c262beeb26a060712f7d536b021a7d28077b2bb2568c252b9a6fc2038be73568beead6381ce5d749436624474538a2a0ce13d0e47445c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h686bde90e63b8d5911db617df158ccc2cf05465db524adbefa9b9eddd71a804a1153a297c551039e7678edf75fa4933396049aab1d8e39b272c0bf7cfe9f07e306d3da372d41bfe8f107d5872fc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb82d19ab7c937bc2d06ae5a8571e53f058ee104efad5124fb70f6f7a6acbd8281c74dd64fb5c73c8d5dcc847db29aca7bece5a7b4962800e13099ec3c2c3fc8b5a640496b667f683751f549adb53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e250c48ec1d4354d338eebdb5562dd6d3c64d68d3f0b6fcd2a42b90a7e9aeeea99c90e15a124ed02ec01a4a144752bbd74f0b2c7cf1ed2408763bf933076bbc18c53049cf8d855ff42c12393c84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ea1e6d709ef97209f8c677065779b4dc0c9312cbfad3a565ca3692b81be27c6d085e16b0bcc6dddd404cebafc788339550c03a726c4c9a18c6ca6af16f6eaade814f2afe615a318417f955f6ee7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1465e2be45f2e1fbb1beb9532b6072434f47b6fe03841a965b952f03c62dc6bcd43e279b43105676cf6e48e6784d348f418364a23808e8232f50101d5fe66aa2aca83dc7aa98cfc5522554d76ddeb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24483ccc5fb3950f59927d7d1742410cb8c8ebb2840176aca807bf42be4d25026be905a6c0b152e485a775a8332fada7a91b87166c142b0846097b1f9772e0da83bdcd111281465e6ba5245a822;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20186149db7c7a8a4b736ab1e3e518fe78f8bef2094341c3105d840c4c1cbf395db542ee5ee062076df6a3575beaa6bf30a9946a48df52f231e017814f02b1c11b907db33d84245a3ce406e4ca79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf818616aca6edd51fbdb12622f1a4f0f798e144eb9adf08b963e352d74309f92d1daaa1032b0a168d2834d93624a23e9a28d07e4d304136620576483e1a48f51a85006c61d8e5121da3811f0681;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13520d89873cd3f3a5cd4fa3abf05b415cc1a7e905ff1d3b763f7fed1753362741885250e2e776b6415664947c3dd1f3a1c796c3255678bab6c4fd3b493c97825d2fc5bbd4d15e59aa0892378ed5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2249c0ff88d1b4d72592e5f9332918e6311f776a216b69041adc738b0b864c4cff3a35da7e91ab7f1de979d3746aa8c08f2072ca41f8738606a725594aab9d8c7cb6722bcb96fbc9fc111fec8c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ed7578171e46eea30aa700318a3ae5780da22354ea674526925a9eda82626f7566d21a17b422174cfb515d145afb917096b14ad4dc60c2afd14c80f22e3f23b1be4f7a4d80e9c81d12cd5654336;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ebd217ec24dc4adcc88f773a194cf7c7298614ee508e307b3dd73888a8723e30def7314582799f2c218ca239840da2e713ab3c9832254b664e86e364d7b8b1e88acb37a63d8651d3b4b74e99207;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1372a1b471c79bfee5368c945b55436605325c651576e1bf718484ee328e18cc7baa22745c7e51d231a4056a2ce7c30a42bd44a2daa7acc33a102a4d69563c1e4342127f01e12e27820f438d0fac6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b6188b62e11e4fee4bb0b6747667ec0db0e8a8254171dda5f6d945e6c2d24b47600c6df961afb8d9fdbb020e1b923c0405c9eaa52aba84fbe0bb7570d18de19b7b55da0f61b55c6a8b4883e6f8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133e2e491be0ce91c1e2fbbf23c7d8b9915a78efa4a5eea67f0976b3e725e926bf12ca12ad82a208a4b87bffcb60ceecedd766f879043ff96212c9434530148945ad87806d0118deda62e72b5a4dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170ab928c3d3bb632eafb258c3e358c89dbcb6bd8e24a3748ced889c53197b37a650d5d12f8e1e27a7853d93db3a445eeab2ee24d644a4a11188f7337bac67e9da0a8c796316cdcd3486b4e0a1c29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d15aa2aba14149876302721c9571b3f641f3e2c827c2e1cec85ff372ad1fd23e78f8715a970086b2b7e683fa96b4697593a068fa3a1f68e9a235250cccbf34aab6bbeffc3c725f3a230a77d6602b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19019b1811284bfd8282ef21fe17fd48991f71e6ac0dc57c3faae57018ebfaac41b0ba923ccb1319d4706f75b76b7af8bcfd83c2111ab30e75e8ab53edb80603fcff4eca3bd601f8dd23e99939c52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a91e3ff44e461a840ab6c3c9407abe12c8bbe83908179db278c9c5876d601a95d39231384f60fe0940bc89330936c3a4b75d0d553a5803444faa2b0bbb1e68038d26ce01563610359ca9d21c5366;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b3d91b9ba7d79d377573faf2a526ae77695684a34a78e9cb24e4eb4d31553fdb87f42c244725a0f29b9a4f6cfbbfde51f168687fb2f1fce78034c900230caf586a7ae57a4d1a19faa9f4bc62ab7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb804df12e4d9a07f85d8f0ccd04818472371bb23fc25caca492232756dc2a2d6bdd74ec73d0b25687af8e77985bb16ff35dd4e659c1ef69ddd690c3c7a421ee044e27024fb93d2be572c088f3568;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b59e52d0a05a52bbd39c5f0b172ce0398f18057f209ce3399b268c1f00ff9e27a945e675c29e7e8ccd4821888d9a114690d18199b40990504aabe0f01db6f5eea3a7800b7523dc3d62a91557113;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99b876590d2607f0cf9111c8e6d86289d3ff2fea94ae8bbf97e08f60c4e4f8ef14f9e836b6528d3248978dee5c333d0e29fafa6a84b425eb87dd2b2be687a7b5f148713456e809049376f00856eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heffe81d78bfa2c134075f87392aa6a729a5ef6986e2b86de4da1837db12339deb1b1865bdd63ba6a79c7ac9dfe217cd505ffee388ebeade5afb88dee90db58c5318784a57590c067125c8f44915b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8580d021d9eaad1821895ecec599d486b17f053e224dbd8838ab84c87b36c4a96a5946283b933bd74a6c7ca8640587dff68b1610d67dd1a9d0aaa7c91c95bd7492fc243cad3c66c164048850f4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2fd5a1c6e46de707fdef9d7c6feeb7146493eab9ac65ec31210403813e081a777454e43d80d07fdb91361f2ade7d12215a4352677578a3de18388d2af472dcaac5cf469005d27659064730246b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e857552849ff70c7177b39e312e44dd681241c0726e05fcbfc6869ec122fc24a17df38150bce97b58a61657b287d7ee284e6ff9c51962a8b51ed91bcbb5bc03d20c728861ea46477cf727f942cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec06e769923f5e1a4e20d321814041e1aad74638911073cb6127332f56aef1ef4fe078a06490d1be6635c5555c1ab6dd85b98c31c673b5fec3f70ca434b3caa3eadbe2f1480d9192d3fc16dc7b8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b38da71d4b46ebe698181e11c0011a26c240a6caca22a6a1ae50b1d6cf3e301a61753ceb273a7ebc02a8e27bad87c4b5525449ba8fe9b81f073165c5c2a72fcc73eccb7366b0d6b200e872fff498;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98d912c6e82c50d688aa3283e6e0fd046206824aae9c1633209662c8913ab50f335567fb3cb5bc3e48aea777a080b1999717ed657e8b1c28ee1ac626f118955b264732e3ed5b0778f64c7388cbfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ec2b32c5a2fdbabb4d4f051e0d4448ed014ad745175942afcb5c78ffd83780ea1514026da8258c3ab8bb860120096d218fec961a2bd65897ac66d05973e39fccae9a219dfe24a69c06d937b3c21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199300a1b6f289e5eac8983b982b1178e90eea2f594bc3126a5e2028cf59ffd823cb5e7ccf6ad2db30d5c875d522bcf7aa665520f51db1d8b07d29a517f66cf192a59a0df58084c40d3dca1918122;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1badcc5f5596b68ab463ea85a0968a328648a978a3c1e889a42a2f037369524827e3116f310551718fdbeb9e54e8431869d437f62ef8d4eab594516d7f6af0e2f1b9057c0f2be92c00fd26a60b119;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154f795ccd00474a033ab68e4ade1537489aa81e61d2b32761ecbe381bd0db6d9215cc408044871fbcaefb23f72f3f43443e905d1664c9e33137d9ae1f958c0d29e108844e8bb98190d4657854d31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h965e5201f954dffa550b5aaaeed858d615891382b41032b27fe2fdeda1d3a39be371f28c19f82ee1cd1df1056502b1d31607e594e304460f2ecbec1ea14a75ec5cfd316366ee2500ce48e5495db3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3e73a45b940163b8974734a4c643f67f3b1920f23ae1db7f0144ac26c4f22783d9c1ac4e0d232e3498dbc6b46d853774e48ab6a5d1d8895d6069b2aac1ee939f068d39bf40712573312f33166ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d7c30330de3f3f3e981586afd3adc007b32a78d55eafd67141f30f4b47cdc36c5a773734a35b5924a84c0e8d306849dbbd8fbd65604e37ddcc056e7110f380b90276aba0fb73cf6b943411120be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b07eb82745a55883fb9f129eecc2bcb4141824e789dda4fb483b6f5bb826706db2cb35c32473340f75cbb3de7128cf956aa5a19390af40878618bfd39fe5c5499cbe450098bbe6f96e37a0cf8a0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f4d14033e75cb985f7745429c4dfa9d8aecd90e032f5d20a90df1a534d1b6ddad4c5fc79a9ccdb16be279785fe031b2141cd790b762b2c59a29c61155f5d12811972100b6944d7bd0b4f06bc03d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h902fafe2b64c70d05ec910024c9108a9e19bcf4e2ddb5499fbe40d978f428f5ae95fca6351302a1b4f2bd974fe25f100e7c0014ff21b7abf680421a8a4c84fccf78b047aadc62892b780ffded44c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a59d6658baf319197664f42ac2b272f2284a25fe24b3e256c25064587e4be76b8c140cd326256a65d6ea8985208fc46d07c102a286c15a25603450a9fa3a51ee75a6a020d0e5131b072e66018f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129261cc2ea1804c3763fb909b2ad38504baa7b4cea4f39582c0461cc6f2013e82e7696261b94553ff273a7a7502eb008ad5434045e96a7f9fe00eb4fd9b8c32a2ccd83e8e20fc9fcb860935e7f86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b73529a8fcbcb981234c836e1ada29773bd6171e11f7d7502a9220ac7aed179cd422e2859961519c0f317d4da49fabac9e74beaa44e1a68a641c5277a9af50564c005ffe6d7727342a733bb2562;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacd52f0353a7d304b1a1e37fc90c1140c46c17310314bec618b773d1480108a327b6efb046ec94e10d63915cfd6c41e7665e7632e70d0be6d2b8197304d0dcfac2c8bce22788fa9897637f44958a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3c62f9ec90eaef75512b2ae5f3334f0537fe2b2148c90a1d50715fe2150ce7e4ad53838496caae534c8a5143b1ffc803ef48d957669581dc5019f2d3fb03c910bd9a40349c77ae96566b6c1d265;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70c4655beabd94cd5afb9a7afdbb31d3d75c5d7187470f912a682452943d83ca5eb6b1c2b796642749637eae5517a31d11b847f2e02dbfff6065c3356630785b1346349b712969b09dfed4fc5ce2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190809213a50a00bdffd5a82efb085984123a088a2350124b3f8945d4470425424c89c822231562c33d550849badacf5dd7032bfcfd795f05b8c82926c2183f45eb82d0f7b03701550ef41a1b023b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h770fc94bd6412ad1ab08ff66fd84bc02b69e629279c6ffa1760932e8f701f7069a4afd61d29fa495f8a75639216b835838ba3f1c5ea713ca819bf141abcd41f40a0550be74a6f3795af2c75ecd2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a23d400e752ea0bba4c2318960f940b28b6b5e2198578a12eb807ccb806a3bb314989f707acdf068d9923ed66cab811c5fc39373b8e95a48a517236b7464dc4ff2222f31d79e09e293667950ac6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4766fc1d471bb4140ebe044ed1acb09efad0af9d902273ce2dff4b63f8a5853d11929956ed74b05655fd4af3169ffbf6674cf74f4da007c0789cdcfeda667fc51ddd8b1c6ba7600b6ec301620b8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d5a462c704d0c17d959f210d071f6f4761e313c111fb7a76337b725200bdf3a4c29f197e4c85b5cf5014118575423257cbf5aa8f7df9a6d574ddcdaa1cef121c74f0f3d01406ec9577f35904abe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ad37105acc043e5d99afdcf40153971812a14df207ffed5accca327766a5bad3b2fb0a80f7fa9a7346fe8c78e98a8b7f624affd09337314bfe34caf5da4f0185c750e48facb12bf52964b9e322e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13fa6a65fe15b6437cd1c4ac3cf411abe41e2675b9edd37344d41f38a9e4784da1296b919e5a6f737d11cc4c43f84269d976166ae8c20cd32ce6bb8a74bb3492247cbd59142f1732ac211686d0df9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f009d4e3d404b44f0124d9305079601feb6966758f1218d80d7677e772094c5ca905e7e00272a3e566b40dec58e0ad0809ffb6d9ea86a2f2c20a96fe273a81fc219cc5b3ae2b5b47769464ddde9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he73a2919e941df0acfd5c5a8c2b2d3d93497d0b44828062b3d885a6d4921a11428c921510f20e5057bf95c5f5ba1a435dc7ddeeb955e712c47560f247deac5896e43f6a47961ac63bce9e063988e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1294c142ba509d8ebd35f01439c1421b6238359b2bb57ec156d1ce16784d50b38eebf6aaef01d19e2e8ff5ba8f9659d9998fbc786cafe7663810a2e0741ea6e951fc023c83c777f28b725cd4cdde6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2edb525f719468b1005d456d1890ef2d32dcdf28a8d8da5bffbaa976aee7bf443f7a3a46ae78d32f1bd86ab39388157ce18478d8b40292f37a6ddff80e851ca7db36919de2e37890a30668a2783;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d583b6f1fccb6515005a21d6bd72af144e4512a38512b891b699fe930fb3f499e12495300941a93abe3c3c8a6b59087264db3f684cac662d250b1745972a3200db176a1d99f44f285649cda06cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f45e830f9bc5ba4ac61c5695dc61852237526165ff5a8fd60833cd40b474b8d510f18136fd0c1299a8c24921d893898e9ba6306cfe116dff63818f8b441029825aa135e176a625c233f51793527;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h403c1e96508dd08ce02c952af650975f990f1947f2eb82b5c46311a9b88147593d5bfb3e5785bb3d7065566d26693ce858a4e6d359cb3734d98c3c45251f25bbd29a9c24b3cffb7eb67cb105782f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a007997d28ce3baa8107f8898e908150deeb2f2b5d3ae844a119a6eea64363c3e9a6c3a620befdae5abe59f03b356b4c45441974b1354d39f4b00ec0725ed2abca15116036f13dcf31014a62d8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b02c609d3efe6ee23a57524cbe0ac986e639df74e46527ca89dc8390da4730c15bf61477a1db131bdbc5e25738790b845ca97aa310233fe94d5e6aceff036bdf43853a85d43277e51a096f9d7869;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee605101dd558618d5334b41eb965527d5e08b47b0f526a54f09ad701d79ecb6d482f9aed7906ece5bb032fd949f8f2a16976a16c53fadf14cb2fa72407f760074eb32989d365db4a51273f95e59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83a3f5930edc8fed99ffdce9347d013084231ce345d1ee4e5ee10550b1116bd26fced8e87c5e8714b7a49149beed0bcb16774b2e1e8c6291ff763d9be4fd243e4d2bc9ad23f6a30643d336661091;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b055f58d8ff19b7231e32597e38fb831a6aaf62dfa35dc0cf88de6bfd2082e4339a9710395a709392a1b9ce11143f300bca1317b68e2e3cdff3dd2c02d3dfc1d4726affb96d051d2702bfb11b43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104173d753b24b0cb80600dd8b23b933e9fffd74b0dba51e052851e13372fcf1335bbd4123237e34e9c2cfd202607af3128816bfb1069fc7158309abe9dffd9d472dbf89b1bb41f08877667a57e5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7a491ce7d15e2aec3c58b2f5f4c596cd1123cec051160e90f21270406920d2101e4962d4e22b103107ced68e07ce5b81e51fe09857cba8e64bba51046a457919f703139092f0349b2d0e279f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90a0334b78b4be052dbef0b4a54bc10ed463f0907367038a433907a06ad59e0232ee3dd1207f7d2e5d2ef142ac5b844ec414af094a9b97622234f7bae4463694e4d6471bce0dc96e465598182a4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cbc5d332da18159f01b6bcd717cef9632bbc44bfeeda0c0e2484877fef0a09d0f760eef79e3843e4075cc2d9539bf1344496581a3abc82274169d325cc8f1ac35bf8c43051825cb5dff53388065;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14888f8576ac0929551834f7dc50969fd8440b4673a0a3ff282925d8b2f7dc140ba5b7b5d54f7fb9d72a02516b8fc17d332dffb7f5789639e97c75e5f9d58479c1f5e38fb62d50aa8432d88fad667;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6be8ac26d3a934d961b2fba0ec4bce0a1dfd565d4130802d0355f1675befebcc1279a83628fe51e156cb9195d5a52ccd6069318eebf96560e7de4e68875e95b6287eb357304c6cd8d685d38fbbf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fea50a5202888c9feb1b83552a573fbcacccbee1526f27b57f575e128248b830de103152581b9d8e1f9e674f89066b3e18daf47ce574e940715a15c8ef77c26e66b1b0aced771a71a67878e4a24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102514fa58765574daa08d1b76ee75c82705597ed502d6299371d6da6f874bb69115854dc0856ed60928fda67078f33913b4f6281a48df766f0ebc631256c43a7e0df901436d284afd7a8564bf346;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd181d1b76c877ce389948f88ed26c51abc6eae2852d539dea157b345ae792390e141a514ad985a8935702d6ddf4fe1ba666157fb2fb2c1e2cfe79de523176f86c0d2693ded88ceea5971cb56fafc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee8612dd79d5e8beaa8357d8517f2bb251a935568a0b9823b1fccb76cd2d1add82cd441914fb0ff4e3a2ceb567026255e8cc97d94ce0a67b7ba0497b04580665832752ce1298d5c6e3ae900e541b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75d6b4a2b68e887d1221b545a7e7ee71219cdb79e5649b9f781d0dda5a93b3f5c2dad77ca0fa8ccc93383e61c3cfe374e49d9839ac4badfd653853d7eab6186b49b8175c65e14c5c2865a8566e68;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d478101b771c7c50e6fcaab83e9a1e56b371e37800ba2139724d5bb9f6ec0213983c301eaa1f055acb0316cc17638f14d30db4b752b7bbb3479b5052d80da400175ffc706310b83f97e3a633f05a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef72eb58b8787ef9c1d6ce699ac23e3cbfb64d41c07f64c904f952166c6c5ff2f0de142992522e8a3740b7c6721364becea5e5aadd51be20406e1a84d2763adafedb7681dbce7035584434cbf8d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he201f27a9da05f0b408e362e9cecc1427fbe1bcaa95158466fbcfbaff0b5f88daeef86d8cb3029f529206f25e51c98f491a3886e200f59a9d3e1cda589a69960024a0e833a1c26d367a0e2c7c52a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3189cf1d80b2120f2123ab551afc4dcd60d1cf54cfe58562c9105a9f34ce825a6ae3981765dae1411deb216cd3a32886ccee7d2d7cbb3ca84e84093a277a1178e9e84197102cfcacafbe056636b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a80f80554401e64f995df24732fb6725c9f05aef2f49b55718a334d70a05699536fb6725da6e4bc49d93da4e637d5295419c5c07c5645b021547a9b085b0bb9869349b07a6674230847f7091140;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd2136a31c373d2aa66ddf9a28f839388600dd86349077bba084a8a6dcfaec64ebba344c63375b61436d75fecbe5735a7012fc98b2655089f1adfce1e1a9a42b35e435f7d874369e25f43a9eab5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5932d43b39048d4e690ff5343a88f0374f8f2127d591d0228526be5431c82c97d16a10f3b92cd450285765501dc1407d23671aba331424d07cab92fac2bdf135daf58c310b526fd90620297d8a9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1589431b02839816ad18a63dfd82848ee8788f0cda2220b5531b6d93f0910dc7faeaea1f84aa6b971ee60d8731d94752c246fe6be8d4c40b0c65fc350be1768099da1b38c2f58989a3ed77aecb8ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167d5abd2541b048cbf60fcbdca50b66564ab1c1587930c6ae6b238ce2366bb30ae67dc63a959b115b2cdf16e4a6a9ce9997f18b2a88f45ceb55671a47fb81eabd95463953f3ac1ef4528294ad530;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0e7bb6d1ebe5d1503fb897072ca5eb3948a4a468769610059bca521a5dde26b756bf8b6c0d81988178e98accc481c31343797a458f8c7b2fabe49faabfcf0709b9e6509f2934439ec08fa715e2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f742700adead6e88d1a7bce226f28e0425e99aec75498521c542b57b715b97e9ec9e4614b437d3a5440f87ef123b923b54ce888b1b686e23eeb06bc4411ed58947de8348cf856ebf916520a299f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131d7f358c409e85c51e9205594f8ce4a28d97787a325b74c99f62509a79230289b952d1607257cabbe425ade70410ce1598c87c0e50519d845db396b48b712cd1bae117bdf35850383a052d89a8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15174737afbeb1ba387857e73551e55ec7a2efd1fe30f012c2018b7045fad50e6de341612ea3fa8971e07596ce4d1de7246c76c17e533be5ac5e90653c3ffa2753dabfb60e66776fe1551d7f18732;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf710d4df3e3123bcf44340bd46ea00ef2cd447ec3ebd3451cd2e6c334ff03a7bb43c205371402adeaf1f8b5a871c658ca375b4d1355eeaea038bc10ac3ad2a289fddc0a0efd8287493387a06f91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1371d7288ef8d26ddcd64a5688c34d3f9d2e937753f4e65e2800bcba71d595a16219d1dfabcdeb6748c19583d3dfaec537e8f9d3e810c3edd84efaa84a0eb82aeb3eb35353dcc68d9f7e582fc6327;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104d9457af85c072b618e47c38bfa614e5452dc33df3d0f5f710528ebb87edf47e4d26a3dc143f8ce62f44ac7991ef979e60b87f0b3cf99dca4e54d943f099b46ab0f73845a26bcf2c7e8ecbb3694;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c81abc2c2d095963bbeb08c4cc592a9ae0a9ff752cf1c85d254dd147e309ad31adcd08a1569e0afff65203d7321dfb53ffec35bae8942202222d50cf25d75496a26abc0950ea2ab05df78adcaa60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fccba4cfe57b556b0bb6ec7eeed634a31e58e87f36193a24a23b7ad664ad3993a43e4a76edff9a3f579d344b2de59bc3ab36bc5bcc6d985504fe316cc7e8822808a0c8614e63bb998ef803bdb8a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6d06b59086f2747e50cf7e8528c585dcc8316779d06840c4f670984c77980d041983597711e383e6d7ef2998c63ca8eed837114ff0faaa2b0ee289a3b3d15eeccf047883842ae59e6a258adddb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181399bd166fa307006b06ddf5ffdee80e56f78deaaa6c3e12585507b39f1364e3a44feb3449e6b146bc3c4aadfa40c1ce43088d49e8793f72c45ba327605398b02cf1e516efb58b34ed92b150aff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b4ab5c92351b19748a60f0f510555b7643be611f6a58ed76d59605090a011a78749ccd8f49d2788f5f13a84419bfe24bd8158b50413166d3ef79bf7053ced573b28046e3192ff4fd5ab5a145bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8af002a713677b34017baab05312eee935f30f1890110fd565a4b2d9c17c1675edaae9ebf5cc4809e8e6b6d55543e68440b70b4ce72f26da24323a3c3e4dcc8050281ba7cc80505369a174049e2a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cb0787b96b93c127d7788b33585fc2ba0a5dacc8271b0ee590452faa77edb04582bede9a0207d4e5774fa62106e2a1c399aac1b455414ae101b53883714f910885edbc6bac6a1950e1e0b4151ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ff1f32cd5b9ded67e28723827f991de1866559b18720b60fcfbe2507ac6e83b89aec0d41506e6d64547ea5757d4f95c6bca33bd0c9d119942390143c2af12896e3c6e17767fbcc37aa4f7626eef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42c687476e13fc925f74a78f07af950dbd8d4bf01373456ee7e8a22f24ba5b62709ca60bbfbefdf7ea05c5fe333b1c9a5311aa66ce24e85330280d877b51408b6e219f43b445733c1e43d1d11f11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10309cff6208e453444968310a54d9f45ab5fe66c5075cf8c675933efdc7cd90c346fac39bdd2acfe3eaa53b61dd2d4f36f851ae898a0a6336121bd82a5f7f647f6be596c8fc90957574dad9efe75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d126e2b9de301379bd5c6899ae59f3537f290f02da6ce641ad147314eb5d2eeecead6ea6008565d5f5fb5798ee5265fff931bc63cf0f7155a86ceac7af43199fb3b48dc990e75b36b8b01ace5b9a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf4c2bf38de9d10558304c7eff6245333b0f672e04a7bb39e535e38afb72ec0c964bcfda4af4f416ef76218a3778e9f13e880b5602f624e17066097623b0fa7323bf7d80bc6ee081f380153e0ede;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f6d7a64d85fc4b14414b9d115013df0c2e2014d3d414a85b78a8b5bbf52290a274f96d0c6bdfaa418eda6dfb21374d22177225213be5e67446b11ba27e16f75dc76092e553836c4f6f12bb228ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ff3b0c7c5445cdd27fa2debe51be2df66b2608ca9ba1441915f01e689dff14744beb70676b60fcaa7c5cccc2ba8b5982b251bc4241e5794fcdd300196cde41ac6487a3102d7b13ff122c930da45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1e4b5f7c23abf6e5e92edb126165f7258b38555c19de19afe9e3f267d72753c019ecab76da3e0c0b68907c588250c0f5c2bb6ff5c0b4cc56605c955c3df04482a63d63e72ff0463753a7bdeaf10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc51409464211c04c6e8de6fe7b8066ea49c3607890a864649b9bb87d0515fb65ea2362b52779d894c6c1dae608e1c2bab8afde450c1a5def6f4ff493507d8d6408fcdb84915f4a39cbc228bf6169;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15cdd8e5a7f1e80ceb99417f6ae384b7734c1725ab4047d4bdc30a98fe9e3753e0b06e43cdeb6e094653df1308a2beb2732ee96a57297f8e385ee05abbab38691821a0613e5ef6d82ec82df60a39a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hade56ca79d2453bd4032ac88b28e771f47d85a23e3d6fe9f2cea300fd0e799adf87e568052df3508a328a1ebb6923b52eaf9da15dbdbcf771020e409ee6c2507e509246bb5281817d10182ae528d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43e978e02848de874c897c3ba99d1e0879b489afa6228f5c9e5c49e5f4a1d925064e51de78540a9333b353867820fc6c0d13a5943c0e64663a0d3fb901d7da0b16d9a71c06cd805bc9b2cbb0637d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1741cc5c310dbf03559ad3d03316e08f627c7dc9f3da71f20616f4d2f4b662aa837e64d365a331671aa857c493219c3cab6d2fe34cef50dc686611edfacc16f5c6904d461c9aaf123e92a41914a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97a4f2c3efb17a7acea895277680401ac7aa77cd80d2a5d42fca5947866a989fea2d67e62da50a9ab96d03e5a081280c1b477d2a21e3a998f49e5dc0063b681fadefbce28b28184cf6b671951f4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4552e6ff0bc8ceeee8bce4b5c0ff4b9b7e12e5fbcec9258fa75646cc4bb530b3d97f6205846b076a008b2ee5010520aadf87bd3364df9b04ba4cf53ef6725b0798ac28120a00d1b3a487cf9359a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd6240ce50c32259a79ad15f4497b9183cf819b02442cb6c26ca8ab903b68c09bf25ee4f84783de37847e22ab5d9b1a2225236fb5e46af713fc9273e741c1446f063072866e755c7f6fcf76447e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb6a0ad4509f2c177b0d4a7da4e0c6370e6045ae2ff1dc397d77c769d6bc882378832f8187f914b725d9461a5aa9b9418269342120cb7ade45cec42b964d4a657729479e3fde13632cc317840c91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0779ded228fe6be44203eea5b6fe1881afd38eb543b084da1bef0b20b4298e6a7134e340daf9dda79789538abbcda3e6b77a1162bb6bf63a73af4863cbda411ae40977740fdc8929b4300b9dffe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d233b28d7ee145cd428fe02f2a81073cede138fc48128a641271d8674735476110a35273cd651a1effb6ce070fc625d54aba337b3fd56990bf1495d20c4448d6663163393dafdf42045c551484b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1214c58f8996f5c299a6da9812f945025d79b0792987667251d0d2b3722653b0164a44d2d7c30f20a7b7bbd97926d8344d84347be439242b43eaca0d2c3c7f01c41c7cf2e22da7613828d090120d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142cf8533e4221537adc9d7bf12b060e3c04b5120c4fd8885ede897503099122b2ee40c75387833eaea7d092d783cc220b9305d59f4f61a60ee998060c818ac4d79263920adedbc5d22888cbee505;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78b3c2f06b7b780244850366805afe2ceae717305c18198c74e6bab5c3f5ec125d8b3aa8fa4caa6d8e630122cb3058f28a4630599bf5cf6979fcd8768be5a3e8f043d3e0cc2d0f42d8909ffc9177;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e31c604b3c4a6a0fd2966e935ac66148e53b2a4bf0643cf3c4292cee01d99b2b6156fe33d366c95c459385f8de89ec7e645f8a814339d0523b78d3c89d48abbebba12f23b3c66d877337b628ea59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc69dcc1269745839d37b0f47010756b0d1f1088de45bd63f56ff3088d689f0d21d8966dd8b1bd625cd16f721e3916d8883f910740ccda8a39531058aeb1b02580007928889c69c982fc491017171;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60a122e5b1570861c80a76f84ea23d0f08b82f7ca9d36569b1dc22b90df2a47fb71a07657eb4e40f5a50a2506e1f666973b9e47e44c3fd8f16cd604ea10ad81a292ec597f6b88172143e65c1ea6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157372db32ea4f0c46d57c2a7f82948f28dcd9062564fe853926bb4aad8c95e081dc054a060426aef0471a8738c7e9130ce21d031a18deb4de001fda141d458f0be8b3d5f73c23a0ad61ec4acbf20;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c664835e8c3a207ca6819fe8d0d14683ff796bc6bee43a5c56b33d3681e1f5c9d210258dc9b9099b7995c361d89cd3129305aa8963d1a2108e90e93ebac1af7706374728a6096636d474db1042ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e89f8f1c392f4ec3344e57c5c62dbd69cca5eff41d4d5b80573b6113472d868e675881741b338164478cce0420062317661440d9af23df963a9e0990c65e88d03ad7f28dee519dc0e5082640c155;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d8fe1efe6232e2178087b7f4d5b96bd03d2ec196268a267970689631c026cc6400fa4a76ba67a75cf222004c0d093b78f703612e08a1f9dae37e2aa08e2b27b988ab16e543a0ce27dbc1479f52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3490005e7a067e27cd063d6bef7af85e9b3afa2aacbd336f63b9781f41061f5bc5b83b60601c5a88cd6ffd8d12f030dec4c1c6852b2b2db9a1391c2933a3360bf41e74a1e067d6a8f777f1ad47a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173f8e403f99be57884051ecdb099a908bae4cbc01b1fdd18f4b0b44d936276871859ce6d2ff4682f7084506ea43c7e11848f0bb08778dde2b44c27c68a1c30ba60edcbb0137f106354d1b2c7cc91;
        #1
        $finish();
    end
endmodule
