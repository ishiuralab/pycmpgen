module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [16:0] src18;
    reg [15:0] src19;
    reg [14:0] src20;
    reg [13:0] src21;
    reg [12:0] src22;
    reg [11:0] src23;
    reg [10:0] src24;
    reg [9:0] src25;
    reg [8:0] src26;
    reg [7:0] src27;
    reg [6:0] src28;
    reg [5:0] src29;
    reg [4:0] src30;
    reg [3:0] src31;
    reg [2:0] src32;
    reg [1:0] src33;
    reg [0:0] src34;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3])<<31) + ((src32[0] + src32[1] + src32[2])<<32) + ((src33[0] + src33[1])<<33) + ((src34[0])<<34);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44534574bae33693612c00f91c0712e32a724c208441a5ea24abfd7eae40db40ae0b5113d28a52b3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c0a2cae77e38d53da56132be64eb39a83af8b61750de5616f0ba17634c843e75cd00ee489387f783;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10d22d5b3e67275a836ef13eae620042a435ae8020bac29813dc6d15ee9adcf80f47d79ff32a9a923;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90edea32424ae8dd8d3f049ddc3b885bf27675216b4ac79cf5f084c8d4ecefb77e95b0aadef4ac9f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dcf206d25fb750819213384b687cea5351f9835928c70d29b0cc0d0d634aabe9b51123f7ca19b4c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h791e5aee6d70870d9cee2c94c93c0eed34bfe2a5864044264b73ff3309e65ad38cf4a8d96db65a781;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81d2d4b30130f6080d893c3207eab6c1853d2a57e808207ad809c08c401faf8466b1ab29f75c750c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6eb025279fa6e0a3961c3e53ab830d5b74a614e389d712a6a36ed68efc83b928ec5ecdf573bfe69f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc515e5191bb6da99bf86b8351ec0554c141b00eebe87e1caec442391ff044b0d41227ff4e8f606204;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he359077edaf85d9b0dcba511fa8652c2c31b1d3a1188deff8149a2094a153039bad00da5d7ef55a7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h228bb2f405400cf4bc5b87934de75eecde6eb74e4d816d5e2703982564d3471c89ab39fd2fd242000;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ad22bcc5a1238a6ec28c01527992ed31406d1351495cb18d34a3c57b090d7b59a5dd866fe523678d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedfbb55ac6b12eabef516afc357b05980795c1478987d58c89219f58db51502637f91cafc27d5b378;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99ee979c032e285e7f123e4c2db370e77ac440d1c572820c77eb26dda00907b0ff8d32f314ec0205f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b0dd33d956b0cb1b039b265d105150826bb0f380a66db687901c072e27e846bf4dccd32c53245399;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23541e670fbee3a7ece1100dc251e013c6a3b531af21b8c5c876cfdaa856f286c02624a45c9abd2c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd054e33c0b97830f52da4fe938bdba2a6b1ef224f45b961fd64be5ee74743dcb53b5610dbbcf834b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f823d321816653a2a4de36d3c65a3c10602a8af97984327638de57d6c4f63c28f018f949ea710d92;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ac1402d5a19ce08120eb9c368c96c4e7891b9ebe81aa570488942f4a3d889d0846544dc980541317;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1239a45c85fecee0a02974a91e15f7445b6f13be50cab597a3d9c3c9a0ca208c1d115f74f96dcd2bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h220a02add7aee27fda718eae90d1b6a84d04211ac40708092b7d1d0ce262a598393a42870ac50a53b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd0776f1e7e56f655c80cfda7198d7bc4c2127baf92847b41a474c3a0d3f6997b70d5e1bf14cdeea0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2d104ff826c327e903a6d5ae29147eeea99062f6a8d709118c5fdacdeedc4b3b820f6e97a481354e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3168204092cb1ac1f9f0d98dc854e641a0f6cccc8954c0134d61b536ac1134832af64afe08a629133;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac0f74f406c5858f0e4cb7a217d42bf90a2a0259b60d935a6ec76c17c2883b936d507ab28e15b8d54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9370bd88656598940f11d4b564f15040e99b167b40baa862bbf4a3b2c5651bee517de19b2a0a3594;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93c8cebfa9f565b9d6dabe616db41044dc2c5f4512654f8c3f2cd925463b901c7ea3051b3c30122a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedfe44b1aa662cf55cf78970d23d76cdfd6271e735678a805b1df105ad5fc56bdc85d6f64978ec66c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h288a0d29b4c8e4547fd2c1ee9074dcc95c688ceea8f176a817d129f1229f927ab4638292fc3b1b199;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h235e1df7441e6abd52006c6e4a146cee9a331923bc69de2cf9c3f06e268a8cd941049c9463db8224d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81d40cfb1a6a78e05f885354e5a9532c53a18c500462e913b131caffafc2c9242bd24c88b4ef3559;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49cf73b74dd02fcfcbf97ed070049f9cf7e7b6f3ea9d6b11c067a488431bdc21afa554500c4ef184e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60d0bf5a64a690db5df51b190d0d3388dfe1dcc757170f1538dbfd5bef4a5225f19a3dce89a48207d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb24659218f8434f6273930c06df89df5302b3889e5d6edde74c31b1a7ddd179585039273b1a0c8ebc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ea89ee9b9c3e0212ec086086311550e7d8f0ce1f30277772e664a4062a69ff89f31eb289dcc29db9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb59bf05b1b9661346dd933ef2dfc72930f331189a7b01f18c67ca71bdeb5490d06dd9ca05a8558fb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h843cb8df27fb8ac3331abc3b1dc7b9ccc4a3cf49186b290c95d8008318af14686d41626baab98c5fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba0abc3ccbca71c2ef9d6324b2abff5e22094975a7d99bce365e28fccf49e3ac33ee0de40f12cbdce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha588996be411ea47905257984f83071e1eeffe0e5bfb8b98d351116587ff38d793aca1a9c4fb20e77;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1962adaf6efb7b6566fa476a367a958f3736cd44493caac196046d19ee83c1f5beb863271369082f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he16c67bbad2fc743c3c418cf67fbcce42b0fed788e042c0f951a00134b007c3dfcb8ad8762a52376e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4150b8591cf0071dda60a7215ea991c7904c7fa9f6cc1b304d8dcc8952cd6565ba0c6e8870ac57e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97367adc7f564e68193af6d102ca88542654302f43428f7a808745363e3be27eaf2b7796256d69357;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9250ed4d80bc6e20c424f16464de1b122ade3f343d46866d8ac265a53d2fa15e577a36985b0de10c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4889378d463c7e55d0cc8684a97ee42ab5667ea4c5810054d72851482e45645c0b92c4e28edeb906;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85dc3dc48741aaf0c5dd9e1048e8d9a5cb116c0acb65240de00d0e9d323ff77b11ce6d2180946d900;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16e3ee8040912a9a79ff58f8da793bd5288675f86136a42eefab63e2b47e0796873b55086de8026d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8677ce7deafe41bd98c70ab6eea6659e1f0c8ac9f1beb104dbd09cd92586a5aa5fe066170994dee2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd6683c4d7dfb2803b2e19a706e6d69bdd8e61215ad3a5331dad79f73b1af0a5a552a00ada01327a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32a5fc9a794ff0a3f8a47b342bd362163f49a8c978baa63821c9b6f569e7a892589870c6979ad7bfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf710ab5e776e7dd819e58d062e9b0720d3cbdef5b9d93cea97a66781b252c908efae4079f0cbcf77b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3553c0d10870726442559b4aacf8b7f3e0b793ead8a9ba2a19bea912e4c526c1d26b3fb83efedfbbb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha74e77ede12853a2916d50dae3584c0406904a9bedfcd868126ff59b9ea5080df24f584e12854e56b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94037b65a5fb096bb005041e8b6843b91138e35ae697c163dfe72a6ac85ec118070bcee25a6347ab0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88f1247f1db035e0b642e98cfaf7283674fbbd54648b6257fbc13b8d627398c7409671589a58b01e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5155deff874d82ef6d528107737f36a4da555d9c8a0c8f7e170a8213b05290e936e516d4e15dcf2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38d22c49d05515f97891b7655ab48763e7e12fe1ed0c439a9d2753f7b76c6c57323c7a1d810fec2b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dabe4ade02e050b5f3490d302967e7ab7229e28219c83292cf85439923b9986a0d83f62927ced837;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4971c25dd389c89889a0ebe067208f59e1d1d81f205ea728bdcc8698259798378020c70a0c8a3a153;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc40d2ad0dafae6b771686252110e16153432bb94d9e77849b6124f63cf478818089181081d72c1766;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12b2e7f828182b6068a7fcbe1a598cb9f0a7c76437f75124b5fcb1882194b416f49d9f1b975816e1c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha40e4547593fac519da591c9c76f24731ee80a25d7e2523a918ece148c6786d23a8c6c6f487f1fdde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6ada1784d41174ee63a3b63b20c7d59bb1704e7e772bb54d0fdb493d689c6b72a7e309d3823e573d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12bb2d4e4c5b7ed248ed883977e72729912c2941041ef8b7b0c0f63060cb3612298ec35bfa06d0ba5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1452840b3214c8d8d4dcb8ee5d613795f58cf261865840a23995c9328ad3cee82c45ccbe9e1dcbf4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4ecd0660651b888eaf26b6c3935b954655e272dbcd438a61500603c12e8c6a0eb2f75d7cb220e7e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b8f02e16953cef00a676d4740d9f102a18b1180a77ca8d60c5d3969c93a66a761275c121691bc04e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda71af861f58ec7b149e5f853a2aefbf0381af7a03683ef3768ba22f6c7bbcabfca838a487cfdd665;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h232b49ce6e3267d85fb28a14553e83174a1b3a9308957088372ef28bc86409c9f07a7b0101956f2ff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb279a50015539f178b3bc0319e0a6b71ede28c3facc21af81d829ca3e316568155c864ee4a249bb45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2477a499333dda95864102a17d8f7a65532f8d25173100bb50b06a69b8e54b59b19b6548c93467f46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cc663bd7d18f9decb57fcc202c7e103fd118945364fcb6c0aead62fb6af2dc9fdeca25138f7b96e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4996b349a636ff4a94ce481f0867399dbdecfcd0fd3cc1a035a7faefc62b75332beb7d1408b8edb84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59a689a62edc36d4a953337be1b4b584d5df77153edde38860d3aa21c346ee7439db22f1c52ba6232;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ea6935924fdb52e44ea2ff729ab60f9e794b9dc2cafd482bed876f79719634a10db560cd0d1fd5f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf35f9f08f168281ffe7cd07d652077faf207891358ba9280d7a8ffcb154f56018fd26a12efc27d20d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha50a24209204246905dda2a80b62dd065ba87052e0b345c4cb1b5275d37cbb2b7cb613123c178f66e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c7503a6866833b52159a20dbba680d9b0a0609c138e1f6e789432844b38f62e3cabcd1c874a1301f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf162c5b30900ccb902c21640d6af7b869089646ddee7b4ca8b54e5b3d55a3c1221d87ae9dcf118b0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc7a4b79d5744857e7870ab3e2f4af6b4240ac68f49d50d635c86136769ac4f1a30f3b7b5aa364220;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h109e42d3f7dabcd0aa5016188477c07304761d9295064e703195ffd44264506ac95dad66ae307d8bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb74742a9f7388a8855b07c702676cc0a4ef1fa485b51742eec96c0e9973a49ad6c5d9c940145c449f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32514b6e799035004cc6d93123582b7c948741bc43494ba0d5176f370c4682f61ce7f776a83ce7f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd003f32c1349b8730c74fefae829fa90b5a0b7d6d8cef66b6dd1559a880b9b75e25316b0cdfe43e39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7785c417dc0e2aa516299a3decdd155488a9f06d82b6d39687ed9d32892a2fa0d4b5f59048b18468f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h149b2100d48567c4ce1984d723aabd779b56b999a9a740dc2dc708f9d7000c2ce288d14980c2279e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb196944b8849ec7fe42c9be68d19b5d388e8d6da68b2e55532924229f51e6aa7009299c54ebaa8718;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc891b16a009f5c716f16c4170907291420d88f61bcd8210e4ab9e32e7027d9a1b55549739a069a8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc9ee3150502a6a1b9f042f58e71b55834d9b7f2c60dc0ab87e9303bc2431c15d2c6697559fe787de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf09c1548a461e4474023ae4f1aa5e6ca5712883b8ef7d2dd51614e2065f9f1979af980c6548cc4fbb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f67625fb9b23d887c3cb36b840493bb10ee92b83eefcf0008eb14861e48dcb6a0e3f340bf748a640;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e36e77e235c5885021e9213dd03e77af8ce8184ff691d2c17b78423fd7c284e1f3bcd5019d49e5d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32e1b56592ba05593aee4d6f10163c5c62dd1d323f1b845b9ea0e59bc7688533443947b16641b7476;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a20f9f4cbf6b333e3cd2b1e7b905759278c711511154ec3913131223990f6762cc0b0077e006f9b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee2dd68806a1dfcd7344a34f60d655ea6cfdb8bfee38ca81bc964f276f039fb251c74f7660ff6fb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e1c7e35db7bd5325240caf524ba11bb73f4372bf8119302e3b3089fd6b1347478208aa276e7772b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a15d6198f4162cc5f102b9ff2211d6eafd183389b38d0371c4382b093f55189165c89e7a82dda7a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9237f5aafead3ef7aff0226fba9e2cd8ddc47fc151b1a36893bc7ae68ed5f526fcab4285089d7924b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dd721539433e8b1e898dfcb18133892d2b0b11fdfb4f3652337ed883ce86e6714e04dde4f43f360a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9ea28b5e5d4f344b0ccc23ccaad14ae06ea22d64866b40a93698ea2e384fd26960025c32c039690d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49677e56de9fdbd89b58d43bad8e07f8ca42afa8eb4a7fc6d0a6327cc4940417f416684e1ae83241d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76da0e041f5ac47755dbd3892db2b41c674080dfdaf99b012e5eaed310bbab4c9d6317451ae31de74;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffc2c029238c5b903ce8c2e79b0d7af5293bad67c4dcae42aa199ed8a6089ba4011d279a8db8f5cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha040238e8a73dd23c9e31e8278d3640dff31cece202519bc8e328b931839649b0a0e28307343e49a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4081096f1d73b2f42e2e257f4334723e164462f519feb292781881486ea90ce38347f2812265a83dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9f137f23fc8d5cbc554aaf25e1fdd59550e51e5a20e3795ad3a4acafb2a9016f5260739eefb26196;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9af52ccf23c034090257db59d87f072500a5fb3c2e6cdcaaee418b11aba792e723046a2142989a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a219a8a7fcd621c19f7e9627a433f812801142857595b2b06587af5e87d03d7aaf59175d122db0cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6582848febf5c70c9616015a6a13ed4af6934e4bf99f85ce23dc83fa0971d082d45e1feaf170cdcd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d426ae8454ed90bd70af0efe9962976104e34f46060da10173aae2cd2b0d1b9ac9b75b8372cf1c5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39b02b52bcd03231be40595d2024f918fc5cd5c5984b1103ad2f0556ef8811364e190744d14455665;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83464269276ae85c17be10049da61ea7208c77e90c5b8d97ffb9f9eb33e21901b8e98abc84389ddb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ca1a5da73d5bba4d282a8424943f5ec5a374afd0b8eba02ec2d1e2358ef5ee9a9a62c6b1fdcb78d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c26c2cb12a5d548c2a32dd0d2e3e45ea58a347e666df39039a334c6422a2c3f4666cc1056e1a9599;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h405d8e13dcbebcd98ce1c7de1d845d96e8692f9f9a675109787b348736267285c7152b9225eda1cf0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98dd1505dd80ef1bd5515d6a6fa8f3aeb0497ce3f767e0839f9251e888999355cd5270c53fd8210ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habfb938b294b6531b5d6723a77e3434aac642e176e3a2d048c0c00f03a78bc3b04eb197eced6db3be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b4f3595e7b3469aa59ad20c81564aa29e9aa4d4a66f3951ee1a3dfe7477d86b71993aabbdcba17e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2a163251d8e3a7112f9411989bf47855239c1a52ff623cf91d6deb9ad3abe6b097561420e44ab79d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c6160bfe6285b42fbd7cacb8b484071571257ea5e4b1b1bfaacecec331f90b0ad32cc5ea082dfc2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c16d58bf917c4e01a9ec51738b29a11adb0bba9176de827a5766007a43595abaa9708339bd602711;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35901efa2addf394351d90243cbab99a8109261b1573331508386b713a0cbb938a2cb9c110b569ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7df6e900bae586e77cf5f941b7960b151348f520eca6ee09758767f12e36b70f3e8cc54d2b4efec54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7389eca905d37191e1a082fd45d4df50e98b532994af72b6b5b2d6c166c5ca2c5ffa8f7e3c1141d6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1df249fd23f319717ada8c3f3b8d287cc29b1e3615571e6eee37ee0415dd27aef86d3b294436fc326;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dd37d320890cfb03444ef4e34fe32a90be34f41621da15d8139e765d43765ccbb8fc4ef85cb40bc9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f30f0971f38824aff938e0737cc7cef5d01a8a298ef46e2db9144c602612fac8dc30bc9c8d2959c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba43e6b70b598c25f0c0464bb7b3d6d94b85290ff9a1b410cd8170e9db9a3800eecbef768007fcc95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8e7873506e249b5271eacfbf4c1558beacb2349e16d121688921698f1b1449a4c632c4d9651759bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a53ea539c70fdcebfa7949ed3eb1e3362479eff8329a8fdf27e7f8b3d06f52b24f92b155cbda7749;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1372d5102e4bacb83c436f5061cd68ce6687cb117b76f6fc680d41b2c1484169bbf7c9c8f9924ad0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bc8a5f345d2131f19d73dfa3286b4eb95074982d7c608406cc2c9246de8ac699221e3b87393ee1d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf2e2d14eed55679e77eb4606b41d96797e14fb197c51579d31f57f3bd6b60910aa43cc412bb6a2f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46dc52a4d18f6ffd41febe28bd91e1dbe269b9a2ba6198b930be24d08b86017dd4789db3f49adb993;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcab0e7a448a8c706991fb19c12e919d8de5d2bde35f373a82c18b602070c87e663683be836fec332d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cb4f5ae009b5b621fb3f19acf464adf98d10d8a8837a5489a3318ea8fe8516fac9763067e311887e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcef63a7ff145c392347ad9ff7d8c2dd0c1872598ec69b9a98a4b5568e9da127d0cf568c064ec90691;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he914b57ef2a2c0babc7044283fbe850818e9592cacd4c3948d55266db195547c068414df6c0c0e4aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3072275aeff176fa445ad1fca58273f2b78e830ac638b475b8889034fed44a36159bda5aa7e51cc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7013748e7c6e3fffbda08681aeaea2be766ad016981c3e760fb97e5c371db24590e10a36747bc1a73;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb3502d855dbeaa6b868c8b14aa3ac75925ba346cd48ba2d4c3de84bbd9f0e47256f8b8446dd4f97a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd268e5463e94825d340548adab25a0cb0076c4c27f578a6579ee5f45251c3c764e7c06ced1d7a9848;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0c19c88c9375a6b39bd364b4ba553dde1ef5788a92da85979b75ffcde857f0e958b979387d252f9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe98507a596fdb9ac4e9ccda19bbe593404aad6892a804b12d353812961de656ceaad54a5a5f0c50b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c3c7e9ab34a5777e1844ccc20534284333c5263501d3ac45cf5a1b8e4d1a39b1c904d85fdc226eed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3756f3653acca5bd745cd67b4a16fa7a0b5ae27bc566b5874c6ba326e67def4bee701419c451754c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b77c763e01a6f940ee4f583a3c37689b11ab4d4cfcd21bf2ef8a3b63df9c5c5e5d344c44c06a5731;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf63cb84284e9483d2d12f2dfab61470cca898c1f5db7cf2f38fdf0137910614df420215dd96e72307;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdce38df90c97b4fe52f6f42e164dc36b72fa0dea3aea31c94575d29fc7a4e4ee43a04a863a5ea4f84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73aa048edefc792c4b73438cacc72c526178df820224a0296543cecda09c484545f89c99f1bf90792;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h488fdaa11470a5e0d530b67782db2d8add88e7778ff61f2aad1cacb7a0e35567564d25a95323227e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38c8802d73e959556a3c21cc77d5ce37195550092e5931cd5358e2526747287dce0660217cca4f263;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5deaa3ab82e102d4f1f7eccb778627352c840eda24a1360679b0f927b14d6cd4a71796d0e39cbd48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ea7e1e994af15382976e50db05fa426437552fc59a9175f0e12d303a05339e7559f84df9ccd90eaa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba7fdfe2864f2b76653b233dd0a51db7723a612c5477e22350baa7e0ae1a3a53ee96e2b2e7191e099;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf40badeecd299b810377e7f2c3a5c8973fdc24fdeab1fad98d6c99e71288bff486c6d65be15569243;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h177fb68d216e8037692cfcea6eb2dd31a77c228c72ae193b410667c26f61c76c8b17ddacc5ee2e848;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3be395fcdf580318a29087ee5a6344ab279b2d8ac2c91cc5db67f12f4faf72bd297d13071cc985db7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a7b5a32d831414c05d24b7c2a103165238fbeeb5ab19ff607b0bd59851fad95cf3d0964b9efdfb82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h476eca0de1244f251503ba5bc31045d81a6e29674b2c4d8b84c48194a97dc46f81108ec4f30d5c1af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61ec906f6233212b1dc355e33160496d19693088cd203eda37b589c5d2cd7ec261c91ef63f978b014;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h255bb4f0d2fc5e606a07da2c134eb8463d7b26138ccdb7f065b7ba0cadfc7a3bcafb5385ed7d73468;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9984c7dc7d8e155b68673079405ea4bedbb6a831e2b920c294063c1afc9ee8159a050bf26008a5c06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10712c69ce4c01ec419ef93ce62b36686c8102e7a8d2926a5ffacea63c30eb33d2949658d6bc4374f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf301370e12d2e54e1a5c9568675c7afe1ca5d8387130417c29c8a5cae1d58fdeb3216a0893d0fc26e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bcfdc5ad755d717041d0b411bcbb6cc4821405ebe045305dd8b39f1865a394bccce529da7aec8cb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f3b653eae4ec72d3e2d202ec3040ac09deef0adb384b43e4e670945c30259d2ba9110e3f54ed5ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6493ca0ef1df1e4c3219b967994d09bde38d644c2151c23472d525bf47c2ce3c3979a9ab64a16743;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5916ebb8407a0d7afb4e32e660977d5fa0dda6266069757c3e6eab3370a78e65611e3707d79e25e43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29cd28188ef31455b48b6abd2fdec85799928d364a41853ef5b2dd082d960c65fa3babe4fa23cc591;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h136a717b3d265d7bd65e936b1f9a89584e40adb34539d3b6d07cf86eda1a52389f003af85f5c45e00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24c31fa78051f15761eff5d89486ca37baa39a571006de5c14c5db5e231da652821a229a4c1f18923;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25ae006f469441390211a61fd79467691e8fbc98446e83fbf83e91f0f2ef05d4e2e0b5407a284099f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff23c6a3f17a78bd158221bbcbaac3f3ffbf8695716ac886fe35653f24b0253b3226afa607c9adad6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6da14a8558a7c851644229549dd2901a26cd159ed3167c00ee24175c54ffb10778b1d337572b059e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccbb15bd738497ac7599e756399e8e0e80b0f7db66eddb4a80b93e6f837f5f3992b5667806ee93144;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5f9e75b961a2c97ec35512cbd3f2fcec3dc2adc35dd617ca2fe0844b23d665ee74360b767c4ce0b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12deb8aee0a9a9e46bec069d2ee70052248d3420932aed15e1f47f46f52fece01487cc158981b585b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfe92ce97a52ee3f6bcfa61faf46f16743531bd4dfae9bc9e23af76e57434a8473e066747e8b994e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b67e4c2d47e850013bae6165e3f724af020b3a99bccf31d52b46a1bc3c80340db24ad2977de41d82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb997c1e431ce0653c08ec8ffe722ebb590969df6ba7aea65c63b5892c2af203863509941c913b0fc6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30daf879fbb9a15a5477c0afa28ec9de88ff5fe269ea58d06dfec5e54c1076121c6e7432710269035;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19816c4cb9dd6ac04cdd1d70f4b725357c2a1cdf906715e7ef1f61b46781680303a2b771f6ce303e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85c3f3c4fafa132bde79d135e0181480e4c7cf2de83d66d66e1d0faa17a2ffa0f7dc06a6ce7e3297b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h890f3f78666257c2e231e127e62b8c11ba57e966deb64863881d4a3cdb83de4b40b02035936385b2d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b3b6ff0d11973ba00bca5895ac36cbfeff6ce622c031fa655eedd0e90497ab6a5be818ad5a693b4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h176f5a72cd2c5cf9ea46180b213a6c190f831c4e00e70cf36f13a51113f5213064fc48c96f7dc2154;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfa401f370f9a81525f600fb4fe710079f56d79daa5efca0bbc0a081fb8ed93ca3cf6dad53a858398;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc6a3050ac4c447c1f1274dcdda9f18d4a22b5c7e3e9e7d4cc81a24e14da0631671e169893ff48412;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h617e102eb6739c9c28e2df4a13c0b624f35a0b647831081bb4667776b30eefb3051ea82812fa41da1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83e2d2443af1e2cc34c639ee4a8da00eea6638564dc9bcb703eed98fda99acfeab5ccb9efd62a12e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc537d8aacae22773533ed70d60db15370a8d8fcdcab80981cf20f67c7c3f40e9a9c1fece1af934f37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc82427404c2686a61fcfaf40552628792128e3854c7e66383653eb8dc90089e78523dc263ff453437;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b05d86116251af1367ff9d04ac0afd42b3e36ab8417016e510b3f6ea9c33dde4774cffe29a551679;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fe2f31bd75da45d067bb6418651ad6aabcb83e2b5c2f8773608226a334b8ff581616127dbf5e2f60;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1ddb70755ef08c060ae9b4732431e0b9424d642a959e1d926d7fd322a51a388379a6bd8dc959c7cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91e64c5ffdf6b52eab9775256fff8f52b674d1c320c797892954a7387f51a1660e42a2bb43130faab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b21c83bf65d413a3e45db9781fb70710829dbdd5af6cbe8b67b52548040c5136bae7cb2251c3f40b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cf2b732b82a5ef564b4518c629f9a57a8992125132a10a8efb8de8aace178ab5a1f5aded57bb4ac0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5f186198b8d0a02fdc9f3debf57fb3b5474d7cb928392a79e99c425f4e440f0f95ab94ac37a4b62e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86748945c7b61e3ab601ade11d1633bb1980dacf23dabeb7001d6bc49896ac2143c3071e7ed979c37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55b2af52c6b9db08739a1d65bad892c0c1216312da26faebf205a0909e0a0a826ecafc0c9aa00a635;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h147751c80176546f4cbaa04c703c8ebbee57edf969f4f6fe87c0722cc95b78fb04bf79fccdce89460;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h258c1c701e32c9fc38750a44f2817321346e2ce404a2fda0ec5b2206c86b710394f8aae3f713c5180;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h988300eaa68a287dbc939e70e592fd1e4c9949b0770ff37c4bc24fe6394bce563378c34e3c24474d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d39a6392e7bb6c6c3f65225f22bc7540fd43da7b1c72be93e0eadcd52e294318ee768ef6bdfecfaa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3b319a54d229c16a219667c3c86e7ae545c9a2ab82cff735483d8649358520ac71b9b87585c3e383;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaaa874e495ab6792b60e6892ef8714fddb65b9f3b6ebeaa52bc9773e8c086e7a3da4309ee7dffd8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3635f13969044817f14d55d764ce2aff5946f0c0d0f6ddd6b36df346849fbf6aae723d65fe84be8a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd296ab1a741623ac2fe10dad481c51821dc8b7eddcf98c379d51ccf9757e4b5ec9d822848c9edb5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2a6c8c55813b746267588a32277fa229a8a1a9f9261388bd6e530da005ff702d0be5887ee857d6de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h340bc8fc2bbc7c727f2b4c9a2295f885b13037ffdc04000c0db28e5accbd1cce84f5bce0577db99b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27b1905f050f3102c68e0696285fde3ec528e8896d78f426a98056abb823813ea21fcf3e17c291c87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h629c72214290c9586e49c30a15d368653fe718749043d6398ec8f7f95ac39cb2de486f222cab68b8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb887b1f38600368937519c18964604e2c5d36a7003a625ff8c9e7cb4d28fa0d824c0b5951eb5da08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9fa44ac49a25a013894fdeb19bf90ecc800e2a7b604ae1449e0d56660917cacdcbc6952499369aa8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h925f1e9114ea36e8420bcb0e822786f3cd6ac054716fd574596c004bdc92de45d566ca28305c5994b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84b5afc5a197613432bb4d71e8da04d095d65fc4352a1659657c476ec4e58fa69590cd5a686942edf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd73687a20f512920b869d00ae18476d772e5732569ef33ff3c1ef0700a338da38078a511fe4f869fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42a7f71d8747deee3bcd8c5bc49ee4eee512e686f5b2d748577946690257c778bf91609b546611fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f9e82991791ada7ba88179de4a2c6a740b50e4f6b4e1febbfbc07fa891af3df159ceaa4951dcb81c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdb7e6f2bd5f57fcc4e36df49aae33f669fd2c9771a73d2bd5b675839781b7808b338147023efae31;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c6baa5b52ddfd7401522062188cc8a4a5d00832230ece27a8fb36c9442d763c36965a2e2205ff56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h698686f9443496be043a7e22a8c5713917d655150577718bd89550c9edcb3d86eb4e48fc1acee41b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb4fb339b201dbf2e5db87725b14a04b91ffa0f1f8dedd8dfb1dd886837812be2d3da75d70b4b2e69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3263ebb3586077079ae8377a20fcf4992bc2d09d7d495098c1e28af92a6bb43d203595e8a643f53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4c45157ef336ee58c1118c8253aa73b7ea623c46fa9122b325dff38868b17acc7b51142076d8986;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe024ee1d5145cbf71c9e6103197d1a93f0c4a3127a64cf3397304aac9dead0fc6c991d2f67631603;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h736fb5a2551fc8ee891042202386f5dc3e8294d3c4ea8eaac4da252512e7c67910a3c4a998010c2e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec564f91e074796a46da13bb57ba55bc32898b7ee991cfa6caa55a83c82a855166bb0ed2b16afbe9e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4d93f56c8aff7a1a2debf4ac921abf47f60166afd17f0ea2684a172422ac33643c62f937b5360c69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5d3db6ab44b1331da387b370a9450d90851ae80fa0f07ba3457d99b00b7f546a2455f2436872f06e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef4cce3e84472e5fa124d202934ba36d89066cfa8b094a17fd70da780f31496ae77d7be45c14c983c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7291495d4623c2f3f3b2e6a8f894ce01f7d93082ba5b3745fc45cf9a2fc3a81cfa4674a58d722a45b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b4783355d4cb2f74196ceeedec5502e90e5984707b663fcc9589e24b3f5be5f77b6089f3d1f0af0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8f72a2887a504261fab18884dafe8b5af0f85318800b373116b84a210bbd10f081bbaec0de22b64d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h556fb136fb810ab071404c257e48fd917f973586bac57e8e6aa4d2f6165a17d99a853fba3faa2d656;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12fe82717142a72c9550e405905b3e61078eecade2b6414215bb4821b234400330d428ff3bcf22ff8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h317fd211e8c8a200967cfb95e874851f8e110a53dccdb671caf43c002f2fdccf489190738667e44d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h228f9c9c5d81ee963395332ce6aac8abfec7d6c47fb0db668a1cceee2df15c90f5fd035fcb51af72f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha76d8af60cd69a3df09c98993d3b3deab056bbd2f6e12c926c510a4869ab472b2f6f1c59f74386247;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h829df4c6f2904950dd81d3656a4c9916470cef4dd839369efd7165cb0df5f3ddb1e686b59743bd734;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4e5d2289e545bc4c1e081f0b1d16b37705d9d30dd7e1cae3468d32f3b720580e7e719d8015fbde90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc833c4b05918aa8ec22d6cd6fd5510f7210a85313dfa00a9f85a993c4cee4f9e3a50c72c941a4cf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6882b76ace2cd8cf191c1fd4f2aa146982910c289310c5a31c4bf888f984b7df7b77c832510ad8cd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6bdacee143c72f1af2dada6af3bdb01b5f011dabcb5ed12643b7521dfd94ce314ee5a5d7bf5e732b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb403ab57a5597e231469bbdb24b18c5d9ebe700c4e0dfda4f8e002c4ee401e89cf58abec6ea157abd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff70e51b2c7a92f732601d97aefd0c5effe100fd992fe96b6b5e9e42d5159849803ca985c093885a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff45bdac7dced45780b2b88f5653026ef2351d2349907ce537429752373bddd7d4ac0d9bbfdf1cebb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h372373d5088dd9626286184a8dde120e4fb67b2b5542ba5cd09c6108fcc1a8387e696f1adb5a7fa0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40f33f0bd4fa9425c711b87255e151b87654530d95e747198cb11101c828f5042c64e5c66ee9580c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c9f4b9b69c6fcc8218b8e2df40c8662e4c26249bbf1a8e7fb3f5f8324df2eafc731e9785318d665d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1a7a636df9ef88c72f3e0f8ec1ac5497db54fcd395f07d5e76cb2bbcdbf67a5d69e8cf8dfa6b24da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54c018e8b0b70d25d16f865ec1e4a595c9b962b6effd7e7af05e3e87dae16a9772d8dfcec5c6ef74b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8741e706c0e4fade414d512c34e243db88891131e4fa92b0c1d96101d6ef31946dc0197dac2f8f1fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf115189b33513a25f973053aa70ab4c0b046e324bed8b442ab78eedbaca9626799e41e4de9c1342c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h397f27d2a912e9c2e3e6710a816493f3691fd22e7b001ee5a1af75d70294c64e2df1b97f597719b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc13da02938e2140a57cbedb1838909bbf8ce3e7902a3f4fd4f3ca0c6c233bfdbc683780cde03db0cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h643330180671ce99046273c6eb78493cabb875c1934242741928277227eb02aa502073e64922874f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaa8561bacc31293f4a0b769d8bb4d57620c62423428de857ae13065d6188d443bda7f44373f5cc1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e36db2560801eca3946771dce2577b015e0395476919fa8fb2a86c58de3a8aebd12f290096b6c63c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbafd8dde3e11e078e812f4c36733634c5d22136f321d745f6f5d7d79d50c280048c97e1605f84a5bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dafc04a9751fff6c524f732ab63a37b0a245f5043654375d346e618c87abc3a52f10273f7db71f35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1ce226769a32c40d57cd504f1b1214b56671b8ebb4cb2fd9c99439fb9663d8115f31b5448bcfd4e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88e592c81e8f8c54bd8180279cf68f887481dd21f4fc73f0544833b67eb3d74cef15522562e4e79a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d750553ae4cee0a640972389db883eab2474fd38bf7cd08e7a4fb5bd57e6256ea8eaacc62f3e6dd1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf27f1403e9c6e0a25f56b8b89b9a44b70b685556e0bab4c614315ab168ad89c430365f31cd20a1505;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d3c4bb760b0597860f43f7943145fc7474b5b1955683df6eb5a2389dbfae886eea28b87ecb104e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d183277a6e9e8c14e1428680d6d43f26d19fa76dfab8f7a8d221fdb515f5c7063b90181e04d590f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a189919004a056cb2d069ee85118296bb601317eb562d058f920bfe3a2b83fc12c8d4b2c9e887918;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e2786219bd644709c673cd1717afff81c9e4fc0b44ffbb6dd11583b1c8889b971b3b73883cfee101;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9e9f7a6cf6829ff6f14a0a214e1dfec71e7d54b221fb0f2177500618da7e75ae4bf3fedf214c4a6b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6989e22e3de66238c97de7fbab3114d056e021846666942386ddf5a954acb4476ec0660041c833889;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h423ebc1770ee38cb7507a83872a61a0475ecc03d1953b83614bf27abcf9df2c30fa7020729da7a841;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae42301c1639d3584b7a162541fe66b473a6790f8c93dee7d6bef190205456453b09c04b9778449be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6a4f631c077785f4d9b3fcaa83e13f51e3cd660e2935f42d3fa1f5e14e08cd5f8bd8c950fb0a9092;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heed28ec3b83198470252d30c0d324dc562b11b2735e183bbfdc304106d999c84a3f011a3c49f512b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f5f528a817f55daecf1d8d2bac996e4d1c577d7f5229786009441570ae24984a461e2f86c8d929ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he22242666c93fa15c90a48d10a4eb3d961e293243d14ee228fe5b10cfc83f36e725ad669fa307bf7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbca73613247a9a693c375de8ba9bd75ba4182bf1ef79807568eef7f75cecc2e0c0eb169533c77735;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf64fb020fd395698bf8e83a3a503393f77872f7ccf55afa00acdcda6c9607243cb04d934dc2750256;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aecc88712bacce53f768ae4097c3f7be51218c2d29d0566a9af32ede41d813f83c6d83005f2fd937;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff208dbfebe04fac3051d2c73a7e7a4d435e1237db49f0f57994b61e40aa510ea2e751475493f904;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2e5178fe8fdda039d4dc42f8d460a7e62b11c83bf71d4fb0ff2312275f85d27fce1409fb269fd356;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd0a13a16c5d53ed0878c2b9aed029932b1d69128356593c3873cef639ee4ed1b13c16a3f36a36e94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa8775f26b9b17148f6cd4299b349fb01fe38642efcb258cdea027217839d5ed4335ba2a16286d1b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9f401c3ff9017fcf79d216c24237cb71fb807f3b18661666bae8c19800f809bff096c78d2fae5b54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16c2253c80e548ce8e1627b3475364ae3eb196f81c4275cf5f09599507763bc3f3c439bde24e19e07;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78ab92323e280d6055364db67a0adc3247aa6b4c3cbb64747f4fa46c626fb7ed0682056f4343df479;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac2fefbb6df2a71efa12d5ab4d2118ee532384dfbf64df59fb5c1bf5a51d821c1241922342fc9ea1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdec8d361607380dd516db44db08e476274a468897f62150b92b3a7866883797b7c8759fbd8d6af6c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf58b751a521962be15c2820e011b478155499ffcffcf286f7fbb9f9bc626dc8fde9e9df10e2d20eeb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fca42b3a0d3c63e53222aa6f2a592f8a21664f299fc02e6aef27e252301534b5fecb55f1cf606e72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f0738116747ab5082fa3efd46a9dba05a857f8e68f6d7229d5ec1bae75764f70d947740b97d51a8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7479804a3347b9dfb31402fd5aa2db0d2beb3d566e2dae336aab46ee6e4129ef1664308700c210d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e7370818602353993c4a8df0b08b5e4742c9b3b4a0ff10190fea7b4a788a33ea97a93203fe4ccf13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfba3a3df9b216815dc009a55128a5e2c95a13d3771da6b73db7857560365522b4b752e7ba70c25d8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc080bae38c37c67050555cb5014888e8b7c12ead82b7349b270c0b18dac270cd9971413df4ef1d6f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff38238ddab3f1fff0bb5f3e92fe98c7ce08cfbd9ad893b3700993e14910a50d4a8b578863fb8a1e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40fae32c02e714be7c470a797c6a12cbf73da89606f3f71967e18bbdb507e131d5bb8a7f060eb259c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33d22b20b1d7d60fd3d033cf2930a43881b70e732d4857c2494d6fdf8a4dd53b8ff91c42d1abb931;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbadaf84163d500354a5fde733b66dc035a8584646d16aa3a31e1289d3273478033719fbbb9fd04ca2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31b637eb734952d8f83e4394127b7c0e6131b4660fee18bc5ba500f121917e03255a4f8bca78612c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9257816a67ffa44729270b390806824b61197ef0c2879ffd7ec41b76e971e51738a690ce3209439c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h226f2f4f61f778c9d91618d423241425fe68074de1ca089f38dd54f4c86d2ca3e5e7072d595b71b27;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h920f028358cfe31d32c084019815f2839718d6a24165715aed29b0e42cd1dd97f2919b7081ed2201;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heade2b0820a0430cb1f58256aa6cf49fb9939404e2006ad50542ba8c5e9728824c92f4e55ee4e9345;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4512bb79814e1afd0a5306e0bcb33021a96858eb60985e7538ec6d29adb073c7dbd051b872ba9f845;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea9879755c2651cb689710876fa804eec59fed1e9ef306c9319eb1c3b9e4bec8f2f7221637948c500;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha21fe73d249a990668c81baefcfed147dfcce661e78f030ff435201aceed14e51f3a0f0d56a0bdffb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a590d448272222d247844791f709b7b905c50fc825b87319ddfecd754ab3ce583f771aca3631248d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7092c19ca7591298b99a1c5824c1b1d95e8d0e6a0df5ff6914d41cf990843ee6da9fbf810d05bdd94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a73f849d5b03a929f8c92cb7b05cc5b28289d440ec37731a1eba729a5f505e28a5f02e7ebbbbb3f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc10a68d83cd028a09566ce0c1c19311284a691f511b21ed3c314160fb0fee603d86e9d0a99dcc6878;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4b765ce62b0a0bb12329f62ed253938f23b9205edbadf1a760710a680e5afc9f6a007b7226661273;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf60be6c2a212757bd723d22e27307829e448768f75c062cbdba189f4b2a7893a184d32cf7601e4780;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4598adcef328c4f8e2cc298150ea432c372c327946954e119f856d5e09ff967d6cb446e9593d4af3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h963a7a2cbbec0920aee3cc08ad007fb127ae0f95d8d1868a966b1a27905afa1430031df361b63d615;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f57562d25ca0f7ecd2b11dd9cb0f4e3ad7f7663374d192733a45408c7324f27bd6a9e3485a3b73e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51ca18f1a2674d7a9eb70fb973eb9e84c45c1198431144000690e2061ce4101282f236e9781c02e08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94ee5c40f209afa3c26c61de09f9a5fa109e3a834ad69b620025601244233c7cfebe890d408abbfb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27602104bea9827f618ef30a99f2c231727561215f0ed6609c2391eba247faf031497ef05af8d43bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16ace62b8329f93f6faa027584e58123ebcf418f74902f5ec71110747b4ae9526577779d3a449ffbf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h780ff435a34a2769db67ffd599e64e1e88b1af4ed5ca917044f5c89ccbc4074b849428b8e91eb70af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d0de6550c52fdfd5291b22a012723ed2e8603678f196a16088265bace60c1c56075c4b0ca3492def;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bd92a1734ca82f9b55bfa65fecc261a8e0d2be4ad2d0d2902e7aefcf054af8c36f72ccb05fded17d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4eb32538d28b976d30377392d37ffce69c41d5fab1a02ff12da4c1af6590b9d8941754707a79a8818;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a4d7fac9da184d5597ff1c5a60186416fd2736effecdc0942a934627764ff6f70117170841ca7e12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41afa7dd403d83780613d025ed84f7fdf26d6a5d2ad9989f6707ee067e58c977a03487c30524130dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a4fba945bc154c465560ea936713769c30fbb58ae129daed0764374d08164b9d5cf4f3f36f18229f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe57ff9a5abf130ac26890de99b9033b4908f26a24308e317c00ca8651bd873eaf34e1766e03f0c34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd730f89599f70f752fc7ed37bbf27ae44dd863ad51c926e2c5352ec63eab360fc1fe1d76df3c5b970;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c08148819b3fdd3fc14f4d3c90097f33ec3dda1cbf0ba0a0433bcbb5bdf86b3467acfad5b04c44e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8a1839de08051199746914dff17c627ed01fd01a8a03f2e2fc43c2474ad7b09686c36315900d1c44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8064f92cc558d584bd98b44835c45e642fdd347310dc2613326dbf8906d98000bd2a84ab5e4051583;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11cc06ed42eadb20112b976869d846d5b41ea4be125eb5326ce0ff85caa28c0a9fcf98fdd04387037;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8395ecd0bd89eb037dcb94344ae644d4c3433802a492e546e1e9b66b39b5a13238a02c08a7aa88561;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h145c529c7d75609cc282f1b67d936f7279de819f611169cd087eff28dca7cd5797c6075e69fd4c560;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ca8f5ca3b833938a7ddb7b68daa015b201f84687dcebda85599c6f51929e6f27403035899cd209e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc661e5a605ab1764790015b8ebf8039361d49c2d86aea842c97eef79d6bf063784d99598481b1d85e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84cfe71b2c754f40dc9d1b8458ba4fb134ce29e5f92663b6ad0b21a2f579fd88813add3732448f1db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h870c6a02567507e8fb975571266992d6e50e58e4758ff698bfd99753121f3aab06bf970f13c9080bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f4044e5fa9c9ee27164ca66657a09e54df77a75326db72c3a77ed10abe088e088f9334f5bfebd7c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb46c01f69d2407f17f3074e92edaf64fda0d8567b9466d1ce751e3874a13258257c425bbede4472a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dadc3be0bc3938107b70ef8d52257be4cc01ebabb9750a6834615fe23e9e05a8c108bf4bb6725b66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h101d028287df92687230cdd3edc6f129a5454f1bb96618d9f6f3b16eddf65440f495461c5e2a1bc2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea8e548f5181f0d29deba28bf6446c20a879d4f3832a030213d47173864ace41621aa7c8951e8ad9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b012ee2b3c4af0a7c210d25f5bef57caf46c187d425b4e95b4f72c3418bd997d88a0709755979a92;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53774bd7de5ce596cd3e6d733591edd83e9906f60b6f1f9cbd5139d309a06e9c7200adc5de0ce8e1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb92b2d1534438a3ee6ecd469811b3a1bae4db4d4b31ce7096518d299dd7f727c349470c24b7128b34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54f9982c8d7c3a4359f3bd544c0aca73e0d89151e274a0c5aefd9e7b095c9c8a9943dc6e556690333;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h499bb57d13065f3db52c5465b017b7ad1585592e19272973c030c87ee0580abb658cd1e690dd8857f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a1901b448f9286de16a2490447e0a8869d7d32e5eaca41c73468f137b01af03d68c90f3f88b93b96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c566481a2d5957e70a43d70c97fe3feeb6b52e2d27a53a48fb0b7ac46bdf46f2d9ace34104452ec0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he848f751f8c9e01794357f45da44620d6cea6a0bdff2b6d94c0f73c988ccbd73b6e13e882c28d1ae4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89a24639db512ca901342c8da0ee6f615174470ac44ecde033be95ce24cc96b3540c5aa36e9476a13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59f1a6e6f57d4a1bd8f01f5cff946fa8706f5b36cd9774bc73f60ed85d3883bfb3796720884bb2e4c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceedc08869d27088f7eae5c4cb0386405a00066125a5d54aa35e7f4369684901a231a63533e80ef4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b2cfcbb2faea3d387af270c0f8f9ee0766e925ff6f6f434146f927d61d3d1e92a3ad7fe8eb081e04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dd5fe977efde2962e7a00920b71b1446e1389427800f3aa0d228d83585931b090ffe48f53f3408a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15e29cac919de5028146d589341ea56efd8a64c66999833c8936cef9ec156b10bd756458ce97ca4e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d10b4d8db902c441eff5f3b26c6978418e7451595761cb9e28f7274f9b96ad9f4cebaeaba5b94062;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18a786898934f601a2576775ab815b066751f9b3ece718ca54ca1f44358051775664839e533fb48d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f885cead6b6b3d2c0876778fbb051c6f85c517046b5c87ca4af094f2225a545caff9529f2f81e2a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9b746bc4809ac60def0f539b7d08777e44da2c115b3a59af71290e0777c403ffaea8dc92ccd9438c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a2d17774bb5d3aee482181e22ff5c5069b208e3a21a39fe004ad7c5b44dd8a002a1bcf06f636a37f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7b7a72aa22f2a419759575d31b16bcd919a62a72ebc85e9dcaa12e646db9c2d0e6cb6aa38766c492;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he146580342e75e34829a356ded40e45bee7a6f7645fec47081327e4628064f0b31e9366f21d5fd3ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bfdf7068773d5b27d7778c5435096ff168af96c76ff4deac8bdffaa5f0100815927c9d52e257d491;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h714fe16d58662c7c6bddf98a259089f0ea96e1196971dd7cbebff42a44b954801b3461e9544692fad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h811190ce35f1b3ae88cb265e6a30ceb3078953c605c8fc867689b194d344c67fd890b06555d5bc6fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5905e756e0fde638aa99a9cca09155a5b67ae5ebd508d494f789fdb274ffc3773c66d6aa4062ce91c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h500bb319ced34bb459d7d707edca6aa438a6361052ba52b2f33570a9610f26b600082110b70758db6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6e01e05be35747e328675837623e2e5b0944f3786a05b20c8d59bf6815dc3e29e38e92cea93b9cdc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29c8f3bc6d51853a050c09df3afec27afc3cbf69260e018d33dd235aaa9d50b4f9e10d306a20de4eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fef542699a537989ed9083ba2bdd25e041c59d39682cea459f86fbda997f6f25228c8b087f83f6dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2716f2ba20b84b6f1b5bb4aac361965ae1e529eff361dfb0ac49fc8644758174d3c91dc458e697625;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b81855af08760cf1cb74d1802825a3576c864d1205b1f76b762e1d3e83b8fd9880beed11d70c921;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfcfb49f2d70967c9923d285795d239178776f50e35a6a5f9e1364433182c60620e45ce642baf2f34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82683aa2b576601cb458dfde486f4763605bc8746ff60daed0e1ef44be5d1349c6227832789e5aa67;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h194e15cf9c04bdde8f646beec57a18dc4bc5c0ed965ca3284539b70e85d1b4cdf6dd8cd2c418bfa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c6eda108a6f2122445ff7318e08869c39da2f1231d253e266d7ba24239f0bb277b617de8bd16c0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9367440e60271d624fc116ee036fd0de7055611a9d375b5c71c65e866ecd9ff151308ebee3c83f5d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca40f6bf55ef750c0770ddbd379a451ef940eb952a1cc84e6a1341ce659c43373e0e38eefaf45a8c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3459a541ff2191dfbaec8f015aee72b00927a771524ded187ebe89e2088a599dff2ae1cb8f2a2c25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73e3ea6f2813bf36a1b62797255c0784d79bdd2114207a354f4d6558c5c8e595c604374441a913153;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7302a7c33d80a7eaf93454ae182db956ab18c4f8c805ac80a2cbdf5a4b99f89f03573393cb8686059;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3b9c1fc607817c6770f4a0e23cf4b55c943b7b4bd9362cb208cd7911eade96a816dab515ecd8333c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd48ea678ba724e97697065c2ee628c594c0d438791e60be1fc92a9cc41140c16069f7c4b776f079b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7250a0a50537d640ac5eba8952fa7768c4e1a5d24522213c3123308fa86a2f8a6976df96ad565636a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8103d49293d1bfae3185dce0e9d38c79bc99e8ccc453461fe4c8d1077a40383085f5677d6bacb5f12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e032187888acf67d09650fc435e82eee60c8c412e3633653f9e848402761877ab575898fb065c802;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba5a6ec2f44f2de68269181fdd4bef47a9b91b2ba022e2b3fba2b88555e0669a8c3b9db93212fcf6f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ae0a6d6ccf0d2ebd60a8c9cc34e52475d9e3d5c8b17ddbe125130cab6b8f691dae925f5eaabf15ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc899337eeb50eced4d76468c78c26f1e336749065f6a6569713934972867da88a9bbe293d5cd9f9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84377d04e83ecca808cd6d8e6dc2d4bb5302cd978b9cde792ef83889527a8aa3bb327128235dbfe13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb49e25809c5c22562fbee0b23f812ed5d791ecf3709e757b5e06121b98f38cbab8b2599c7ca78ca7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98a1deda775aabcf6bdc21ae2fdeb28e17a126585fe11102d9c902443e72d6f180be6931dcecf5c19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8154c4e0211b77eaa92e266a3fec9fe8800148242dbc1bac6e9cfdc022f73eba63ab8f01db2aa9488;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2a7565188e7897b91c0dc3882fdeb1855d96515d2198a95da2027be8a9f6de0a74453e2923b96993;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae192a2f4f1b65cff10af0197dd40d6456fda361c5efddd5e2628b6c918fac719c7184ca1720bceee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9841f186682df56c15c666fd85cb5e4c667a1ecd93055ad745494f15852d717ad9ab4deb7f53a3ad2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3883755703c666becd784d9b8cb51d731c9fb6e6ed7d813bbe3184085a9ddf2c04c4adfe671fd12bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2323cd2bacae177032dec1c67178804f8bd5a5c8948035ce63bb84961b4fd4ac8c5b9931c3a9d6a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcecae317b5c7e7121532636674918c3848ed4c267f70cefd134b25d62d29b558fc87864254aa82b04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443307e1bf6c21cbe21d398cf2738aa83bd4e6294edc2df67b29e373fc8d1a7f122a690f1862764d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18077f58751217a06b4b85ef51d94c81efda86cf73f24dbd8585168a3eacd06a6bfc6412f7a0302da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa925ba269f3acd0530a548251da9e43d4f1f81bb86a3c12db4782018e18d214d15d906378b43afd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f32c0e75e24f8299ba74a4e9ab86ad1eb0b9cae4cfd61eb729fd88639c7d5862f5733cf613aa33aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51c2bd5f576a236739896c6624a71d95cbb4a384e8d812dd00c75c962e319b8cece29fa6ff7abd985;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30f877219ad45b171f78619247f5fee26345102f87d48091a0dc6e87f82dba689290e4581968a8b81;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ca1f63467f31e6e448211a4659172b88a9be8307228fbeab5181ac3b2cd0769d0f6ff26b2443ee94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1880236a40d1df586b7b30476c265ab753c616ecb8a4f67cfdd2a5871cbb265a97acb7d108f5e95e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb8fe45e3d157c5b360cd644868f4dd211ba3f46c270f88c3705eb12a24da497d023cf48bfa2b047a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84edc7c23da5052e46da2b58e22ee267a4cf4a56890eb951030d8704c2158bad82bbfcaa0551ce562;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h582e07f474669c68cd1639f5415cb2b634ddb99114cccc3a4b92a51ece7e02c740dc9eaa417828ba2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59ef5d6bacc2c1da579d532036607cad1540e36ad6e5add3a18e2a68af568620f17e2cadc27825758;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7ada654e4197e2338c3f264abea66a0e7acfbfbc6eb8744d72296430870d8e6264c206df92726e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd67a9760219a9f6545b758345fe98ba66fdc60b806951f817bfb89e1c1c07310296be25924716a1a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67a17f90d6c608ecb9fe42869548c7fb49a4ce7d82ac7d2778a3fcdbaf4f13b206c742ffe8af9af5a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28036aebaec183019573657250e405a975c8db341a109dfd20447b950c785335b8bde4dab47f406a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2b46c6cb36429129d98777117eb1ddba0c5091ad4bc52e99677ef7a5c1c2eadfd3d4f10ce6132cf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h519ba60cffd7f56abcfaaec8a5ee8c1c7ecb03a23c6192410c398b13aaf3afb875110dc9fada1ab9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27ba0e2aa89dcc7d7745ba0b06aa4f83b06ca7414389b5962776834614080ba2423e28efcd2d53982;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cc3f1788e54ca8c866d24138d05e68fee764710144792cefd5c10d3fc96e61bccd144ca4076eedd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b4a43c43991cf6476612cec26012233b3cac9249fd0c6ce48e98a528bbd434d0724c8dfb73ed1b8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc009d7689e807eb73f09dbde3f66d2a763a09d8e43d5ec26afac0a9df2ac597e21d48979aaedc5b53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde75bf52d9f9002842d3501b61806691b63051b0945b4adb0763b50a5a55c5635c452ac5a91cf3d00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3b350fbebf5e4f9c25d5ade849a7fecbc34255ae6a41f4ae61b3d50fb4a95f02f90b41cce5b520ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d4d20bbba86a4e8c1c449dc7a113aa3ff5fb6001bc133f54eebfb749cbdfa2dbe4803c69f6fde595;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc11e00172a5f435fe0a8b793f84491017413b62a346b008864d650e6cce3af9f4e27929109cafdf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd27339371285390be52f15da7662bf1ff426d6453d8f023eb47fd216fe0e2668c5d8257234c09b63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h473d9746e44144779cdd285b56ed5d7d29bfa0e2768fc32471af105be2d32c2a4b6c552d150bf0184;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3599d03a8350754bd230899250a404fad8a479b7d7c0068705335cfc288a81b48e3c8f4e914d071d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9acd8e1c7a7201dd1565886e1547c8e70b08761cab1d00f754bf3b608b72c3789d4730f7bee4ac940;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h792531439925fc0e20f931d7f783c6c81a8949e3ed435804aa28570571bb8049cae87739e4faeb83b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97cf170bb587df053bd6c9750aa277e122896317ea6813c78e8818f92edf0bf97cd55638d12f9f260;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d6bcb5293d88edfcc91da6b9c6e513727014455982f284af228255efb4d6b1e81aca0871319b303b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65622fd63d52934adbdcd7342442b21c9f5c688a64ab92a4748a66cc6a65b49f146ec321b4328af9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacf908f15d9ab6f6f2df53729158206a69981248f8fb68593d0ff282c04cd7f78bcf94c9258360d51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heeff15588f19adcac229303770dbf5d5c85b3819f94536da04590c866bfa4a7c88b5c710ab8029fa6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97e2f9d272e90e1c89dfe94a9102d1cc97a153398b26947f9ba4a98d523e83ccbeaa93eb168cef96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha09ea85777ff765e3dad44f0e19730537a737e71c2a19f3e8f6a305c288320277268d7f2e68785a6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd503d4e2c871f0fcfb0b3764ab4e26b2d3283492c4aa0816373f7c512b6f889a3c68b4e60ab001b0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cd6d6261b65f1462d8d3f6947407f3963857df8fbfc63c2cf85c96b7c35ff984b39c0044bdcc39dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h824b449be0df3790162be167d446a78f1f9d805d9a73f9a30fa489acdc152376bc85dd1a4e57b747c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86f1031f1a19f8d5f80e4e5e9376e256af9807d9924f1b542269108894a2cd1e6f53bb370a4e4db65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f9ffda367eba73c3ae3c69bd7f7387e597c39f89eb59760b4257c98bf6e1579fe747eb674218f021;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38a8c444f9df9b1075d1f2c5bc5a3ed2af8ff216bebd3b82552b14c6f5c11adc59f32b42186edcf29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7df437202c1148b8a5ea3378367d8d43aa6df1adad038e53cf1b19c469ecfe6cc5734c854d350175;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61826e07f664eca6c3094a6a6f54055d3d83bc07da60826281abc85d6395376f64bbbffce740cddb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h434f717e157909dbd41f2dc1b42e17cb0911c12dce23059afb403454ae30562db875a7966e6c79323;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h470ee98e9482d4e7677d797132c06078d671aea4bc2576142782b0745e4341ee91179a62571d736b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4afed8706289ca89aff2edbb3be517a82ecedbe879967947b2376e1836d2ca869ffd2ba11f36464;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h712d16cabcbe1a92fa134641d4244028bff773ed2efe96a0f912bdec96ed9857e76f40f5f62396b40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e1de6e1c3d0c0757f7db6d917aebbcf7d404320c8604efc55b7e7ca62be264ec7aadd7b7a0a04540;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h882ada80e7d034b6ee01c81ff00d7c562ab6a04b694cebc4e1c660dcc172b8eee46829cfe025c52c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa0028e35e4424d4d9c5a0b91b9f78886762437d50e8a999a7e9a1ad53614107662fc53291c09b831;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbdbcb1383fd2551e667e57f26d92e5d195d9069fa1e6883e87e9848f8635f775f1a42311c8a3b8c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4298f129602b91acbd8a681f7e28840982d53f82e5935840fce2738b86dc5053af04a979b2117caee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h176342b8bbed7eb465866236f311517c022a9669b7023700ffb233618d572400dff0a44fd95eb6a32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha60684582e6719ca3f57f8a45fc290e7c1c51f1553e0b4e37aa2e6261a6a8700df9fd91b216c59a82;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc441d76d4238d4b64dc2b1012b7e5fb19fdb6a8f074bfb852570e6b50e910e06493c05a0ca7586842;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9849a2a85fc19f97b41c2978ca748125cb7ac07386d2843d236c7bf3b67666ca7942c4f120f53a636;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58f125820763e4dbda9285c6d1ce6773f0e267f9e848f07075297a2344e59623a6588954126cd4ddd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd28c5ebd9442344787e99bc215c0532c3e2141ac45c31285882abcb4e1195bab350759749a163f7b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he80cff039c005aafe9c06de3ce19b27dce6dd99dfa994151e4a88eb49ab0426016191760412e7e158;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1fd5bd5d74a0abb756ec7b4c91e3d4352a5b3bd2f91487dadea7900431580f87e5858b8a4dbcc7e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fed59f54650daebe6c2d4da03d3c69b7e68c47c379b4a4db4579fb17bf17997022b754ffb9e41fa9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc117618da02ce64a6f0d574d8a2c848439a6774033f3b528a9e04b5d1e03a29aab2f630bed715cd22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h497b54ee7ad133d913a589807266c044760da423679070869f7ad7bf982f83cd84ed975106c3cc421;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f6354ee416909926c9b354e057cee7f89654a75530700b7fff7cd2ce95e1d7e8e18e222d75ca499c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79ac7af6322f09a81eae4d38d64fb673ffe982dc8ebd3af7d5844c2b53603272f411d841a00078c54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9445b1d951338fd9cca8b83959535bba1c9d77eda847bdfba60367f539984cfb724f3aee7afefb50;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18ddb64fccf3b1400734c60121eff8e9d2fced147c7a19df4089b847b97f205edc8ca4b06fd3f8e5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h621315c3279d71c0afe483ef9b885d3cce2fc12c7245fea3bb68f95cd5eddca4be162b6a31e0bde64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h709709f1f49fb6a10cedb8e70b780244f7ad3e79a9f91936e346830a26e7d18792d82c81ab800fe53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha04a308263d77bef27f235f33276b03e8ae4777e76d11cfcf30a23eac89d1fdb0eb65ea4240b01650;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10434e43c57b70939c9b4e1bdc3c2db0ecb7ee4d758143286638a67f3ba8c6f1d7c9859c01bf59429;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf117810bd8f885dbc4a2407c5afaf2597e9f5727568397e7abafe5011980e0a9875e2623314c2fffe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fc1d17527911b7ad0526d2e0a818101bcb563ef01a75b40142780f2107a77afb5d3dd531d588410c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63783317942bc5b529d30f2301821a1ecf7f37816ac283b7959e59ffeb5654e70019288ed683b1e21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd63c90d1d7b3af4a62a58aa81fcec7ec9007ebda2ac63caabddc84e3c7424bc87d5f9d6de52983b1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h355ac8c24dc79e4703f08be5f267ea7668298b97938a4bb723685b74eb262042786b5e84e9252408b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6edf896a1be932efbe37d07d3f22d342fb70be9f595d1c1b8e8406d0ce21c5257455dabe2398f1285;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1ec4b1e7514621d14f2c26cedb4b3b91794846b6be60436f32949c495b0957a6676938fa7042274d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b23ad544e997a441e5e81c9956759249e8f75f217aa627278cde1f0e48a801a7e7840e22880f2581;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haec33a06862c20f30288bf0bcd8b70bbfda35f9f13bd4646dcec1592974c3fcef55f752873adee442;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h507696e44b0987a1b873b51a26c6a1a703c12c404b4763423837feb9b86f6f8ed5113af6259648864;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf61a9e98d59c887a3787cc9010ef9b7c93c2e9980b332223c81e72ac6f93af147264f9e8590a91d3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d2985eb6dc54e378e76c48de1c4d66e9c74633c92500f5978e2d27d7c13808c00520d9ce3a6150ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb13be991ffde6d9dca396da7235c9a18eb60ca64d762da52787950b01ed128d32319fe56b309abea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca3c45b7e85eea47d8fc105bb3eba8125b837e9ea1eb449ea965ba0a5eb942bd1f30fb8c3aa1daa53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc90bae6e67effd3d780c4d3729947c984d5a14d03687f757b697a08b8e31c73e9ac27752823e68298;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h533c4259ab69187420f3e79fe1c226a04b5ec71653b24c2c0d642f6e4d52e63c70b3308a6baf69893;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddc692858270ff32de9351ef564fa2205cd37581449f760da32bb47c33c88dd2594f53630fef7e057;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fb96a8f2c476c4917080f1be853174ada6a4466ef05161c1e6af4238f00b14b6f0702b6129490320;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf084ce6075e98111a7520771732f587d96a75b464b26bb4659adee098ac58ea4e80aef1271e52f4a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heccc040ab22b90a26d286e4d632d93e49ea84679d8c9b1dd9a8a3dc25e45ff11be7d707dfea0e6b96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11f646bf9a36e91ea1e2c4574451481fd9179e17f2aebb43dfce69baa7d3f870297cf1cd0a335858;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4ed06d94604d774db2730e3f75666a110e963e2cb9a2a7255e104ac648b565b430d25641c61679da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87ac5737a242d49a5c8229ccf00cd881ac694b3b81d3684667540a7c87b1cc8b4297885514e109c7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf13a796af2b7d3548918addba62b5a3a36367b09ea605776ee468b63f8ada8797207ebb4aa8ef12c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he57c95591e95f6d4097402cae3f75b61c2c67e7cb2397215772863dacb01979b9a5117b653f1ac7a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9ddd75130c92754a78443c89caa461c2a537ff3866e5bb10d72b8186be40998013930defca1f2692;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65d1e9b7fa435c718a0a51cfae1dada761b45e12b53cb43c3d2127956cc92f5ae995af36d38fa8674;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78b48b10035c3e008f9169d13feae9da4d6dd5bd9a8a00128c41eaf193115f29457629bea087261d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h612b5d6f011a8f92f97c8135ca686e842995e3057316c93bc63d68cbe751ac69a96d77f7a88f89508;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51e37746a49388a7e7aed3f39ef91ab0140b03a02658f99515461a834c80deed55a0ca1b216439975;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42f96a46a44047172ccf330e61c86c1e2216042e2d646f6e6ac9143a2fa8e5ded169bc072e232385c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77db2d88e77fb18dfbec61008607ed4421e78689d33481fc25ccd28255e150fd260ab023960544198;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ef885636b641fba9ea4f3e29abd6ca794fa59cfeea36f4be2810e051ccff7c6dacbad6464c22875f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30dbec90a77ead2da9f5983ee9063995814682a856d801a79fb10a4dcaffb46717d3ddedc2e50f786;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86372d4682db0956aea9c2a222fd611f6994de63b05b7e8af980ea355b0d3a4f1e57160cb90cd16c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha604ea90ec8a7decdff02fce8f1a888ef31fa768f77edc4034488a9a4180dcf84895ce21c8c6cf1ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0d33d32be49888d814104c848871bc61cdeb7d8a831cc6ba8385e8e7257c4df9a72fde8f7cc47c0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae21a16b792cc682422323d290fdcc94c5c70210077abb3d9cd775c31dac43b2f56eed3fe982c070e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d93cec5b15beb645cdd8eb9f861ec22a89418e96dd746b9a68d450a2dbad021ad5a5deabe612dc6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4d70bdeb9854f2fb29ef8b757f7282ba00e006cc069f7e422c438f8e3aeed7056be2eb1239856a55;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a6e97fe6c1c2767aeeaea6b03bf3a6eeb269f1cf78e2767ece19a99d95232647cdb7e6e57aef19c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78351a37b33e9a5f5d2c13052c7288902991b1614a8325797197433c0e6d37c2654452a3e42670c89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb82a779700757f7e72feec1325fd45af954ee98e6289f654317fb188dc87339aa0b0525d11ede08f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bf09e9d43f770b97639240a3445b31123f3c684dd7f13c6e97e74c8507d748255e2d4f85fac88249;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdec150b63875a6317855a19db6b3c60c4523270acc78de7e1b55dcbf63b2bf8c5203eb77d1e82e1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h160050928ad902a00bc93301cd63a529701eb1eaa61430a4e18f44fd28a06a337b41321a19ede88b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c256aea3490b95da6b3c684afedb1b0398be9b6dd667b7e0bc0255f0217db95a639702fa4a59764e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h728ba18627aa701cacdfe95d4f2b534923be4735aa6b962b0bbe7d3678dd878c150f91a5dca4b6f1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habdab613659179b29bc8648ac5aa3fada51a831ea9d367d6ff54a0a7469a8995cdd8bdc5b4952d330;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec65720ef2c92cdad36def5e25a6f9c78b7ea997ae53224ba63b5bac372a7323a068e83eac5d0330b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86a012b260ec3c62d413ce790825f2c0518a57e16e3b00aa1ca28b701661235e6fab4102fcd06738e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80d05bc7ee1a4f30b3fe710b10bdffdb7b4bda17fca384ba758f13085f1f2b4e909106344c3e80ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5497ae92efb4c757901cb3aba7dbc0767637c6e823be59fbec294ca8c1c2d67735fa9405e9dc69de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ff28f95914de920a8ce7ffaa84e56df0dea4a06663811c3b9d639879470d3f3aa969ebff5c2fb301;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33b8aa9672ecc9ca8e279702bae0574e1eac5b56dbe03e8294815c429e7f02fd4b44657af738bc2a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcba3fd70d49ebbe508519ff232487899d2a8481d14b9fc7e5d99d7980cd9f262c863e05dd3679a6f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ed1f1342968e81fb22a2a639e1011c724442707efd257b4f25ac931d1b1a44dd1b7c62bd6f2dd231;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd66ee1cbf6b45b89dbd85a5f04383d6915e2488a495ee9d0c34ef5656482e360f403d84d33d97b18b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f7963a55becacdf860ccbc4e335a8ac5a631120d7d84901158927bbcc9217fad54a5ab89e147802e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e48d3f9151f586f6cf473bd66fc965a575920d5321161753acc29942e19f964023de173422e433dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76fd459d9bde7c69b5e22d9f2230f699a6d40881edeacd2f865e090de626cb9042fa0aa290cb4285e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he24639d4a44a44e9a0766b6024ea6248476ce538da4e019cb23e9a5048d26a5d65db738c10dfaf9e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc487d31c1f4fdae9391674b0e8fd440cd3556ce4ba5db4864bc3880f3164a99cab3a958c7a648fb05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca5e96315f46b4d256873084b2d338e800c848063abef450b31806a9e1ec813f70fa0e06d24b87cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f11ffb7c6200c5d3d79d4d880bf1eab9ffbd72ea5a0e1d3588174c77d30580cfe288da10eeb790c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fde18cd4beeb9acbce5d1e9e1a503b17d564574ba48eddcf4e08ffff78c040142d5df66d334389ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88bf435086ec3cf60b13c4521562eb4d020e26a01b535ef43f9d3bb49f1a93ca2099dc3717fc055b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f5486d531124cf50b044db336334105de3dc9ea9da4886b62be35864bb73a41eddf4ddc2b14439ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7be55a2bee5b4fa7fa219b2a5a7a276b1fe50b0095682acaeb4497c71d037df31fbfb55347a37fbd9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbfc1c4ebe8017ab7be1c94e5edf43dd7b9228b95704d0a71cc604d15383c0f680873166447cfee1c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee2ba9b53495fb411d7a1b02d4c1611296c9cd81d80e3cca3b3476c19425dc16e40ab4257c571e3e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7236035b86858b93c52e62dc9e60c48e78261dd8d53efff6b10bed341b6a74372e823c0e51f7d0198;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce3f7a8fd4504d0c2bb31dabe998743991ce12922997bac455e7c115c8c1a8cab1f673c16b905c691;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30471a6a22bc7156f3b062efd5f38235192312b7d8f45e343c59afd453164fcfad1efec9ad5f0ec3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc7cb6c657da0dd0a6b63a892bec00825f3a0861b1ef5f4e25832c6459ccc99b659551f7e4d45a382;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f288b4af1bdbe0b741515878aa18e416ae6b432ef3e4bc105e9853e6ed72ca28c67b1b001a084c18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb839d89b1096529f9e5ea1592231fdae6d4f49565afea7b42a3914eb28ed3713fe5433b77cd57b770;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h560616715dd1c066167f620ac310eb6d16e8b531b2b5b6fb641ce556989c391c13dda82cbdc7973af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8315fdde638c73b05eea3aa999203fc01220fd70c656f298319793b1015d786fce89f73ff8ce6b88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h450d7a59a265293e8979dcc31d329a3e550a87a632825824ce5460a4aabc97f4c1bf559673c49cc12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefc36aac62192182b860e1d25b4719321c44fa5f57dfa7719e7fa7e7a6e83bbf3f135d5fe6788c3be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb56ecf833704340308c3732867c7913c9e4522dce09927e16a0b503eadfe00cae13240848b983ac04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89a7e35b1c8c603a0f57c3b8073e6dba86e3351ad339999e160103419c63f1ed93ef7e543a922f4c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17620ba7a876dbb92ef844bbce73574e0f0fd83345e47f27678cf6ab433cf51f2ac6b68f86b1a0f57;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb82ffb0079e5e95cefae8fc70e7202d36d43be795aa8a99a4839eec9716d02a1fcec3c6c2aaf45dda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33061ee1f3503afe2b9d65efddc8da11e59ada9f3fe4ed77cabae840b6335858db7b1540c56d1e060;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4e7da101c93ea2b8f9ca625ae453387b7d38ce1cd65b1272992c5a7fabef2c22e57964151ec0c13c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a32e0247e35b2589347a7623be582ca0d1c22621fcdd1ca61683ebac0b5c4074d74e572420e2c156;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2512ecdfda4e44ca6bc323abdf3732ddc016eac4cd1b8a0e8039266e7915e9d477d76e6367bba6328;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec171c8a03f9e17528fe363d315e7eaf20867e552040ac9067563bde7b8ee711a9653e9c0efd41140;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64b628d837ee3f4946069a58ec232f2bde1df4c2cca3659463ef6e5063777e5d2372b1ad17161924c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8191b48e7efaaeb40992595c254793089ee0e21ad0163c645062e612d4f3f2e59ba59c855c2d2c820;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c035aeb77444ccb5c3032dde487f4a89479170327c6a567e89fb5a938377dd4eff5006a35400142;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c7fb6c4163d0cbac046423b56d458e40b31204190023e1294193f234adfae0ac1e3dbd703949c16e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h864e1e6eacc8e262571f25a81f0de158ad1bb5a2a44d63af41bdb75476c150d17fae6ccb1ce67320a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf86fb56441e2bb338f6d91c914b2b17c597469183da31d7fcf26ae46cb9e59da7def1a9dcb9ea0068;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf676fea677a24c3b0c2c53b9e6612c36d42c00dd3256727fc89df3d542e6c217fe2508f56763c3699;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13e64536c993b3d1aa1265707b08c3ecbc02bd9ed0fb0171ea43e83e369d02bd6251d9c4054c52c2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he04245e4c069bca7fa4a135289c88c88452985c8cd05f8a5a2d4068f677adac61971e224c2e5355af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c333e81420d36e660684e85a3e7b7cfa71c68b6a4557fbb56fac40276596fb1cbecbc80f43a4ff79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18c66f98886d6c406ec5056b64ce01edb879b50f914f230ef8c75710ae53f4db9c54972cb081f47c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf73e7c31a0ed77b57217ca27a4b4675b7d53abc292e48994dde963e47c8dcfa05f06335ebd30194f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88a5f88b09d7adc964cb519ccde497f5c53120d2b8339dc4f5fcbe25b5005f25d3b653b6a7a3ff4e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9454cc307352d9e45d1d40c79daa2e6a052350496e09df3093bd95e10dcf9e74f328390a5e84040d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d35bab9c388073af9b9b19130c58c9343375146a5a84b2291e0310436dc8425852c99d210a70a056;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc3de7d9905653c8de5dfeb3a907e57948c149d8cad9c6f312c492a5d1d37774474906e9e2cd72ced;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e1c0d11b07932a6ed46248eddd066ed3e55a31c14d2420846df69f0e4c3c15fe46ea69384de103d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fc67260d0c060deac16ae94967c436690d3a394123c2df6bb0f6271aed1b43116fb8c3e6543af8cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c5f7f99bc5075307779d1282435a06c69b1b732236f2e6bea5e55b2a9cfac8e444830ffe5469535a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b88fae097d4d7588b937dd11b7856f8decfb588ef4b8c30ae640cf798fd8d2fbb511d23ea03b1767;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3f21a59a5de4238d55cc22d11020229adb140bb80944ea2aefd7f59a65768011289c9f3b7fad3cde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34005c3dd6337d9a982b940ffb8ebae66c90f7d8cf58e51116414b7419eb73da6a700d58f53d85f2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53ffe92ad1b0d8aefd169ba36c003a83d9d07c9b8eb351c8b8a0badf1919315ece9a1e53bc7f8dd9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h303246dd43e878118d63968b8d988996f8a0c98f08f34412bfb4265755ec8d81c6669da3bd74637bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha602cd3cfd23158e10cae3fb56121eb1c71bc04233eaa60a9c5629e13511791f455ec1a6d76f830ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcfdff885e4ee03d966c6fa35038a1c92db10020f5fd6273bc563e80dedd5d4a8d89ffd6aab6fb3f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3034b51ca1e673d7e5805ba997d978b1456299713a6dd5fe953231ae985d3b62a26dd3e6101c42ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ab3e424e555eb7d134e96581db5ef2d613f3c5ac15da07a3707c6f68a661256b9e5266f57bb22191;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha57ac4e853fa027a5572c890efe372374ade8d6267664e2409453d034ea27d41e8589aa90a205ab07;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0346339bd20deea376f235b2c5d324b03657bf2a0f8df43901479631ff9c2bb59140a06af1ee1137;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc337f107eaa840dd069dd2797ea4d9fd954a38679fdc3ab41b735ec5bc5f7f24ebfa2a496b0370535;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h933bc007e5ba8b8c56b65d6b003370d7960e3bb6e1c24d496610badb61ecb361379d2c18a53134c62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb4c7abdd96d67b4e1dbc2e2b7875ad7a3d05614e83eaa4d9d01344cc0f1db05331469d56a33a4220;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffa6651dfc347356a529718f5b6d05fa35803d0c8ae6a6ddf7d3cd6df86bd18a22b51ebb252941dc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb58c6b8cebcb8852d14045cb1f25beee25d134c072e4099544d7f0c7dbaff74b2809623c9ba9a308;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b34252f33ff1577ecc9a349fc2155d4aa56e13f3b8e6e16bbe2b723f90db33bbb900ff4f139fda3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4ef6d5c493cc1ec1c90d8b6c4ff253761dbfe6091d4d42b63a103a59556a00e231a87c0740776a4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23903050ad845b5b40d5f69cc50c340622b4db2ce150b7e693e0a77e6226fb0645646167ad6e8be40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h938162b2d1b0fbdfddc57dbee989b23124ad2eafc396b395b3f11572efb6bc697244145a1bce5fc47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d73eb65478eed6cc8975f74ff527944cf4de790626370d4189578a507b61c56b5dbb720a6253c57d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95c5db2eac974f7bb6c49a3e4422ef4672bb50f61aee467113ce1c8b4d93034e6aa692e1a3167c8af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb01603b9a176f768d66041a7efb7676d70515c17a58e9dad16ec619c8a1b12262a7db45ec4f832ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h160fccfb0f59be1c8456070009c75d5b3f65e9607439a662f1fc7930a16a01f9853cdbad11f351a1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h570e8443d51036766e111145634c9f02259b03ef505b9ab03dc41945215b39a2229118646f75c9068;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0ff824a3bfe7e6a78129f013f10c45804f9dc2931c9df5e8127f48ff09e17fd636cdafcf966d4086;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0251e7e1a049ad2b5b6c6472feed3d7bfd71dfe7c9edb99ffc8b52685b694665e2d9c518c4303198;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb025434ecdce7dd8cfb29308ea5f534f77df52226047023bbd43ba09e2aae73f66f14b693e54acb5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h251acd61e4fda00e650dc2e2a73e6dfe22b220e89d32ed08ef1275e713a4b5cef4879cd30474896cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b3bd9314b65420b936fa32bacb91d6254f9958e8133e6d95a15b51eab4fc3c0c780787e8f9cf99e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb120e9f4fdb80fbf02d3fd80e122174e9577c750a057c2e004da513ceecf3e74e400402c00a3cea8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c3094d33926cc502a4c7ab14ee521a83b9c72c25c098d4d12a5db4b921d862800cd97149452f3ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc537e79206fb36370f17f72649468002c7ae14401b2f9a2768452d1c4ed075fce8853569ced0ab31d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9f159e38e797e0507f6a9971865fee82ee3834715b3b0b57ee6180ae6641d5596f51ad4bf68a2062;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfebf22ce652e9640c10ab33f94c70a69c3e54a7733d0fdda012bf98b416f21ac7e4370afc77b16734;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h745d65d0ea2715635f65203d69ae5bebad9d691af79f548a6c672c93dc9891c229d87f97baa3ccb3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8f24f6de2802b8609707ab2ef3620312a4be7390ca36d8ec260a7d684dfb641e2e2043cd27974a42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d620f4b405a2c869f120d8cea4c5955a1cb9736f99687222f02277cd02d6d94da64b73e34eb26546;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bd54f07145d8032e484298dcfe33bdab3dd9fc5dc8654ceb2808bf61260f9bb918a6482aff527fda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e9097984338a53652742a9d24a06901b57f1c28c888ba0d038e6b491385d544c74ae79d02bc22224;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h134c4c422cb2d3f432e029b86f443db462f8a44403ea265faaac50d1c5460ee7609693f2bd105de6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be6e57375413fd39a1a6129f8e50f94152f7c83a8a56269be51e8d15b964c54de12c0cf20f42f26e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc29bbbde2252f514419aaa5c2c575569a409cc925e9ac04fd73dbdaf422b6429a8a78d44d357ec06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf25c8dd94ac4f3794bc1253b2dd6da967d0502264f2bdef50d4af3dcfa5393b88932dc80a406abdc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf82b323a316ff35eeac5dcf4d9fbc953ed96d80cb968b2b900976c33289f0aa8cde350a33f16e99c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0045eb9f0830720c70c100d603500e99faaba6c6a8438d964e4578f64c18a2d1e820321711eec536;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a659bde9b0a648b53f53b64b13eae038d87fdfbd9a47775a3a54b208f80a20ed3e2e1e22cdbec8c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27610ba2df3c4490bef6681f5e460fbf98cfe4c8d26aa30ab284d7bfebaa0a722dba658b94fcb0879;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44243b1b2f3bc37e0d2a8066265fbda586e98b46f64817cd3337a95ee4213a10ed8deec49f2b76862;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d5c4dd72ac015af1d7fdd8c31324fb0f138660207d7da02d8d0510cdc2cc4aabf7375ea72bd8575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcf66f1b26d4bac4b61921f90cf1e37c7deea8431fafcdd00303b710de500a2af8f670b74073aa56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe9610d9d5d197eb763016644d00a20781277865a99d8979704843cfd9cda6a57747187e3ac809653;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h592cf3685d2028110000f280a79b839b70f48e21c9ed207e0935712874a42dab453098c0094d6689b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93ba6205369977e98ef623fa4f16f6d8aaf5b0e1fddd77f369acb5e9d50516d58aa5baabcdcc4494;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4636f7acba695877a4ad84f6b37897441294629185b27a74b45e013d138a4a15c7cd28a2003260c4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6fca3870aee98081481956ae0cbf571c4c56b2d4b5fa08cb503b5ab692b35160d233cec84cf9b77;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24498d44584e3097f74bb647cc8b40171f8a6727b8f886c0688729d91ddad50af29e218276246e510;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78440cbae5528eb282326703ad680811b49ba3ad04593923923c088296ab780ca177be1786983e911;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h235e1415579457401c6d5cf3904b994dd32d8f914654bbe17d15552b223dfa40ad42c526cb4be853b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7c4124c4cc72dd4905a87c60583c4750add3eba5e5a48959c81623dda03ff5108cd1ada4b497686b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f647691fcf9e179c0d1c1e814c6906db2dd82906ce3de072ecc55257a3625fcb56dbe9405acf735c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5a5ed1264040ca7d60f8a339404589ccd5e35360b8ebac2ce57a1a2ded105886ddf1c0fefc4a57f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab6c56104a295def2ec4d86551ebbe38368581c3eeb9978f2b36348c2a222ac893bf6e48ff674db53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3650a90db2cbc47b6e6b8f6f14d8cd24d31a8f3fcf837472f8d850cb2c8c171b5c2715e2e00ab35b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24224efd411825245075ae2edb8446492697db5d0027083c1f8145d2f91b0f02d38e2b81b10553eea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h432f47823459fdb10e54dd9664e2818304ec6f05f119c474084bf683aae1e3da9a7601689901014c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h419dfa40689d6741b3e6024a55f8c91d3832b4803cf39d5bb95a1451e6e0970f143aee673f5923b4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5395c51ad0beae19d6d641ce6933d58e45abdfe5273983061befdd067b5332dacdc6d2460f0bf90be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd682505ace3ed5358f57180c95de40b71624209cfa8dfe5546e31edbe73fc929e782baf984cb11ecc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c5a2152d3058f43e37122de284be369ff38fc0b3e6ac4db3d275eb7dbfd3bdfcab3d224ebf6c3e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf533bbf3081940c18869370cddc34e87ac220587d171a9a760dba8d1d5e6eb4a8e2ea736327765a5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5888588c303e437226f52dc3a69fc9c715921bf5203e270d785d2bf92d976898d240f7cbcf4e9e41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd89c935cd155df3e023cfd2501ea91e6266fcd12832bc78362934a7a82ea829ab78c1e1d944cfda52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1626a67c82c5d9d918f6aaa9d4ccac75c32fc63b50e198f8c4b5da6f4d89791e6c8c05fce2f5b3431;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57baeef5c3470e1ea2e4123f1182594ea20d42dfb63d28fc2c18c00334b1e875ec43e27b2176a1c5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42fc621a0317943525f4ab2e190620eff8ba9fbf2f01387538c82e326f46106a96f00f107bad40615;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha21d6151c3542dd15afa88126911901648e5344d922d75b055a85316e6f2a9b0873dd04bc8bd65a47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4de354dff590b10ea5d8a52d81163ce88d587fedefb0e05581dc02db79215daaa261b0097bbcedc4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h119bdb4544c74ab1a5631be111b804618dc7f583dc7df4db6953da5f3cd375679ac3fb52810c49f8a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16e4995dbf884ec971035e502dbb1234f66ca7d9203182743102f4eae9cc59d9e4d91241895390565;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d0112bcd4e33c9f4008d90920a47179553371f9e243b0812bb4974fc772e996c7ef9070e75ed4c84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe885e99b56b292679f25a0528428ffa4f25079d3c1af98757d6ca89cdb64db01fc840b8cf9f561d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h613c2ac429b6e00426867ba69098459111bf4d8f6cec9d24cb30e2f8e056b765606adabe12e80c86;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb615bdeb2525bcc673e4872a6f19cdfc8fb73179f439c14abf929ce0cb4950e8e5ad87f96db41314;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b66be74a040b010df0631be0cd86093b021047dc9f58b8ed6f33a6fd4119ecbed2be32803afb378b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc56255a741fa0f2b2585e59e28193b376e49bb86d4bc1465e59073c517c013bf89412224191c23b2d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfae8430d657df2efb353d8212cb5704594f60f7e70c0b253b1a8ed423c9d07966504b96b19099138b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha01e4b570f5146b9e0ea8509d01e978505db52f083eab0c3c9fa8d0230951d1b705dd2969ba633edb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf36c71056b358878cced68536988b1596ce6eb4db308011ae738a2663048f1e775752498dc8b3290;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19db6b32c8dcec6a21cdbbe631eb28c10c7bde2d411766844f773c35cfe549b1ac58b439b692c05dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fd4284fc5d50d25093bf72be2fb3459bc8376501887f834d2fe2b9b352d4a09a690fb012f3592e0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1ceab4cd61f774bd0cd58a0526d226f04e2561e58747d150c1d849ad15c1619d0e50fa68bde2683b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h549ee998e1f183b0712c8a1a2131281fbaae76e086644742d033d2661a14c9c1d53258dea1d9bd92d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h129df81b75b566b6e99bda0e9f70a6cc0653f815ff57132c08ccfc0e07671ab6641c88b8214c321fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a427051aee84495e799fe2394313ed99fa737352e32c1a9c2f3552d29f84cab9e481823b703aac1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29d13510f1988f56d4a0d99e7e638de87578b5e3dcc787b05baa4ecdd8dcfed55f1168dac81c1b477;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19eee79b792193894b6491170de5106bbe6ad2a915ba20badc0dc6b6ae15ce4e77a63b7bf0bd71bf9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92475e9642324039a447092324bc669a0d940d862149357a54a9221baa52cf1f9155a2141bd57c134;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdccb7981077b7d596c2f143ee62880e71acd8e7635d5e2baf49ebdf0479ad3fa5aa8ef0528ba551d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c00d5e0b6e365874f96d4292dafbe5f42b1b8bd56e07750790338baa5a5470d6ed20562d2aa3867a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57fc22d1022f9bb2be3dadd1c1d7ece55cce0b5d4d017c6773670fd953388f2177a3e0f847edc3c64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab45248c2db691e1374542a4739608111ab408cce63e67fdef77020c355e0a25ef44a8de5be95d23d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95f13296cf331a32b63190741e871d3b7c156fd5e79c21f2b1e3d233abb24a4f208ab181e44f0ff62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e341f99e5965a280cc8140424601be5112ddd24b13018185de0d110809ea484b93aeaf9404da88d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h316b9e095a0fc30b60923c17e774937ebd095b99081e6a7c017260bdaebd269d03d695f90daaf7074;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0b43f0f0a34bd056f37b6c638415fda228073da7f1b4436fb9e60030e59730535f6e2784fbd12b8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8997a553576013474a244979fd3a016cf6e9bf846ac158fd7815406b7819978598045ee4faefcb789;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4d0a0afd54736967e9cc8e1109489f068cec9356b1bd34197dae1b484b992f600c21be59c33c6688;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73520373ece3aa12dd4d64f1bc3e224f06f07ef3d1255ed9bd67aad18531bd10a640d5d10063b3127;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95adf4265ff8a535ed7369d03e102334aa0499aaab4c6a83eb0e492e180b14be44cad038e3f5555e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc954165440b5f1847935fa5e990628f0a49ee60784e056aa220d6e0fb11b72d8f137bf3a27a96889b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8feb3f983ee58805db782babc01f336276f405e71846be8a35c17cd88ef9832e4daebae97d17736f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7d4bf111930aaf794311467b5a38ee58c6d6baec5684751dff3b54ef580686fdb1f9758014ab5650;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e31ec3adbe0aff5b2e6d8c65ebc54c8e46cdb3978e0d0cfe5447197ee768ccd1f4986bb9f7dfb0f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h222a4924fd54f643e20b863aba195f4c491e5794a896cef25869509622f80a98006acf1cb7acb1927;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbacbe798cd1ebb3ff7eeb63a66e430f99f5442c5418291e263eafc3654552edb538a5744b5d903ea8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha83c5743c9837e85b5a26302d74d8be5e7ec140cd4a12f0b66de4b1abd1c2cf2e33f5f84df1917b40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fa8270f1bc10733d0f221ce80b4e04bafefb9f80beddeb570d15839b5a7ac437ad3dc249e942e4e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18fe2b505278415b170f949a5161f6062a10fc34710fcc5b5e69acb10a1007aea180452cbb4f9e979;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ebe78df5de9b648b68b153f7c63ae465fa692cafce6ef395c5aad5fb2c1a8876ae8493558bee5168;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha93fcca00298e76ff20615d5fb2d8f517db396e60ef66fa20188844dd028951a637be04bd3a97f911;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15b2245a8ea897e235b03f38075a1b7a1fe5999103805c7d7569ab5704aa64cf321ee509b267bf7a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a7f963590990587e0fc6df9c62fa5786ca68e2114db2ebd79225f274b516adf1f4f5d44eec9872eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3da6b2f04592d0c0787a793ba0a3fc1147ea70024de2c6d39247c64c670083af7f1cc773b4d51153c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4573edf0bdc7335f835f6f0879226909b6d0ebf3886b64fd9dac185ee77fb2430beea199a374af9fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be2832d493f5191d63d102cb3ca018f609f222d6cef8a18a78b4f0cd8bcc9e25021758554a97a335;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a210ecf8b99ebe25b186417eb66d277ede988c4b9c102751d9fc964e687e30b6bbd58ac019250515;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ae92c556af7f072b3f5c55a385be5bde2bd33453d20d755b70bc41f8a597b4c47f5b53c684e1e403;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd685a8302b49e31e9d7c3f4d2c929d43b82461611c790820eb3a2a4688acaedb6f127123471f2688d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb94f6acd9048077e92684d9ec82b9a7baee21ff7433fd2bd4a0bc187a347690728618b235410168f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6834cc50abb5cc711d064603e531d82550a2d61011a99443a1639e9a2cdf6ed67500d521839a883b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb67243fc389906deb787584e626ee0c0f78cad19e41a2fc209f3c68fcc166d5fa22101ac083563dcf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47455a62be314ed0ef29c56c1d93a690310cc56b908711454b7c333b85112bbcad875774340c49056;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba37090cdf5bff9e0f05b8ba45c23e7223cef9467d524ed09b099a2f9ac397a8a1279bc00c0298e4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h280a65b517593c5e868fb62626d5451dae84cf1e15902866b0f1458bb3db282cdb6e421cd2c160679;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36ffdf75f7189f60171a8c7605ce01f8fa3b615c21dc6ea3e3e05f23063381172a3235e8db6cc7646;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac1ed683e8e2cee89239b984fd8b5ba81815831d88c4bf2c1d23e6d07fe83ea085101bd9ab8499b40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e0d36678b07e327d213e2062b4e982348b82aa1ccbe0f5bb7ecbf229962faef56b22dc9a2408c4c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39b4ebc31d5eae619457c400ae4c52c5fa7db81567f00817e1afe7e7dc047e9d3d418609373b16b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79c81549c8c175cba5371b52f871ce7a168aa61bbb9a1eecc203802d8828a78b6fb7500de071d24f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55e7a84d1dd9980fe3e51c463359daa1101b1bb29d3ddc696a958e7f38d1571dfb7c4695beff1309f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heae857adbf266a5cb6d20ae1d909ed444ebf3cb70dfe089b3e2f819a44f839da4533211e13e69cd42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8347e0832ac4912568993d31f6b026d9835facce743ec26c937e8c369c27109ffeadcc0c3aae24556;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69ed8370e503a8cfc5a28589d197347b7a45607a68593344c741fdeeabf722744fe13453c4c3a364f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h943a18ea394cf9daa65c77ec5564dd5dc3334dc7b753b09604390410eaa294b39ac68b7bbbd85ff40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0a81e931007b7c92b2e5442385a832371df1c29de076cf06499411bc84bfa6d31ebb7cc2f3d9d79e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha79c258bef0db7a5b0e9ecf18c2a87b62cbd9f312e2200be096e41ee3e0966b90f08778b91b5a4ed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3ef884186ae241fda20c19f5c4c5f0012414d6a5b087a93a6d01f6b3bf7cd6bad7dff3675cacb4a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac7add071bdd797176f7f30199a1182be80468a870571ccfce95b2244fb0ae2306c6ccdeca1cb6214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he13bc78486cbf78d45b12124bea2847ad9114ba9bc7659a92c3000b41c0c1dafd6b5f0cb1085d866c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h505e25af9d7774d6a38ddce93af60db02d8069669efec3944a55471f5b156db5941fb430c9bcbd04c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf639d726311cfd60cafe34307789dd3f6a25a5a6d1c4ff7b77adbf210b29f5e98c42a888531f535c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd77c4984d62fae26b2fac6fc3cbb8a01d40816bb10c0c5c4e4f29a828e46d698ab53e778548911915;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aa3a956e4eed53c3eec215f3c6cb50a2c391ed34df0c08c1f639f63efb86cda5b0d26d801025bd2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfb6b5a1cfb742bd48e3d4734f63622ad0b9725554b95d7473a4d654dfb9df033ae32a09d54c5f848;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeae4171803936f6fb92558400d9b078da5cc9d8e97afdec55f8d2fb7d4eef2514803fd6ca1ea9e3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h148493be96e2507c2e734b1e9f84fcc1b27fedf6f1003c486ecabbf2e2a0509a5e8d86a7477d56c8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6559911385f485f1f5238c0a9b315b0598b7ae42ad425f5e9f8ea3930ebc472eb63420535d0782bf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha254f1fcfff4885a5151eef2a08b57f67822c944fe1cea087a7581efa9510acb369ace290e97bffc8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79b78cf3a3959d4d08d928ada419a2c97bf4a67c5fb460fd945076b28243f1fc72ca4a4411f910400;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7240b82e71330a8da1e7f6e1dad5ee94c3c3b7099c1230c8a1c3d72dd2331df359b0a5550e3eee5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha16f3d7a625ab5a6a66f4c89228c8fdfec3db1a45af496dd950a0f2d37b06e52911d1ed9822092c21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55dbec0d8898e76980e9f5a2b358a560027ca0e7b3dfcd4cfd7cc37cea61d165f793a407d124873be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d3cf17e27600f9c71c78a5b6b7100d203afbc74e5bd8cf29528bebf0920af570a90e125e4f04169b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e04831f40f33529633584313643e7dc920fc7267f0d023621a22997099f65629fd79689be9915ca4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e8a63e2a7ded1f9a8f9f548254eaed4b712514c182a5ac69f7d3c6b97d2d176f98719c1e2f5eee49;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heaa0e09a7796cb96255e16ba6436f6ef2c357046a24e068eebc7cc1ccef93006717757a172fc2ae81;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9741b59864bf674382515e01d07fb37135934039d9d964d634330771b2cbf5c99ffed57a527149a18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a8a6568e352f43589f1567143b17c7fbd41d094a5de7a22a1d52972f1bc5a7df56598a8842b1dc6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed2450c6adf9e27fff85d6d4604ff2ab1e8725cb1293b30f667671c1451df3f13fba255fd6dce4d45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5f43e0afaf50820fc5e16482baf3c7a964c663fbf92dce54f90a722b4cc21c55e79322aee194b1de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a91b293030f422228498438c725345ffb78733a301d173e3e16254aebcac1ea0e0b7173e83a5b73f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha71efd8b25cb56c83be27d565114ac3e5b32967a0580911d465ebe20109fb9051957203f588d1f89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76bea0a95d4f7a8562d141767e07105d8e79a632c3b139cdc6660328f0fdb127e24a95509a88c6070;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf79fb75b92d46635159f947c37c2c8c3bd00fc4c5e3de960a377bc6d44aff157c280923e79b6408eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15c9737030501300f4a2017b84a5fad25600584cd313e5737211b60e03db3f424680ebda99b4fd456;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfba209e6643714d91a960ef44075c316c88bc11a4b7f8086f924657243dac697d70c6034b61f56db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6edf6c5f15d5744ea1e358b4213947c0ce9c1888fa8a8ab4d35cbf222dc83ce9930773365606c1aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3eb8f6e781c5f3b48b4e9a747b2ace80a10c12a2652cc5604e31bb4e960f92f9fa81e539f20aa5eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc033670381f2a5ecdf058d60b0d97357a7f8e3626e70edb031d901b48a614effa5e2e6025e90c50d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99b12aff153e31b4ca978cc52ff4b7af4f6bfaa79cb9b4fc14871b407b7db93e7f1732bc8d4da3e80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9d9a105629882e56e6881b3363ed2108af4cfc864b1fdcd38f50dd22ecc823a8a247b2e9eabe36c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h305c0aea35c3e9c87ad5b0b228ec28d86e1280bcc3d6186d2a56c55e9b640b6a0e45e55e560e43f7c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba5c2dcd861f42ebf2aebe18b7af58a36987b7f1318a6f4e34c1c3471c6cc730f9afd0592e5ef8575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h588e2f434d5e8e8ab9c882544c1b9fbc1ae941f5c695882ef94b4785e001024f4a4668c14e055f4fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c23e29e2044acf41c01abe3d18266801f7eb29ffc325bcf40b9c9fd60bb71bd90e19c67baf748165;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0cba5fb341d40710f1c816afda5a8b1dbffb381f9e188e49ca0f90816cca119b38b62ad1a9b90340;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5a85313a4a1a6fe77a556a040af3007bc745ec30bcc0ce0c53923b53a356e8ae331043dd7ab069a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5490c001f2ad23e2d863fc71830b142af78bd11b20378ba925b0df3c4e47b2462762995c0ca6581de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20549cc97dedec86631d0cca3765371eb310fc9da229b70f7aee9d5f4a51081ee31ad4e098a74ba31;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3431f697238b28748f798c084573d623bf85365942dae44dacb92dac4f9d0b9f54532016b2dac0c60;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f463006f98fc7c8176bf94d1147aa56cf8d2e717f99aa43599d855cfe9227945e4e3aa14955cc495;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e1e533f198e61dee81313089005d4bd6299eed82220932d90cdf69b103c97586bfe137dea3343bf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7b5cc9b97d15f9b8b63929a2a2766efc7d3de85270c29ff8348f2a3cf2c2c2b92801131738b8bbd5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a9a3ff045e35efe6c31eda5df5def5d80f8676f40cbf39e179c928abede68efccd6c8509d08577b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28492dfffad0082af160c259c6e0a2d8c7c14ef94d6eaa5eb9e073b8348f066bfd5a3917c77c47f87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2cd2b9bbad8de6f2106773f54ad797ecc1cf7750ec7349bd164cccaca740389a7643be400efc3541;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb67921215a4b7db2728f379563d29913eaf680a3bc97b6bb108cba54fcd3843c0b6240b02dc6dfb04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98160b8262d9db7373ca0130049b9d33c9ed6c3f2f9a3eaecb524b2b1d0ea8460e3aae5953e40b3fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50c05c7827162462032aba422d1081d33f3ed10130213da6f6c7d71f82597375c0b11e588e12bd2af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22e946bf2dfa5812621b5e72a61e14c3f73eb03f3bf39ec8c19ddaa71e0e9ab96b4ce6153d7f65fcc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f9277bfa13b8efe6499c4acd891187b768ed6e9e10b57ba6a1104ad87954b4d17faf4b6d6d8f57b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cf7f981625fd1c82995cd67c11312fd2d5b6a82af0fe2a4aab6291a917ec5c2d23138e19de374f86;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38befc7705d24d3246f834f95753cf0e1e470b1171e225fa5ae04c1ebde6b5a0c3fdf439a5b77e32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb006dac019e2650e18918397639cbc0683898ff24d3d029a82ebe69ace4f0beab62de0a4587cbaec1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d9e6859496dc8b1ec57169538985f15fd803b4751f26aa10b67e542b922bdc56a1d159a617e58e57;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he840552143d0441c96d6d7b55e0bccc5b4b00fc510edd216c03e903e72e505d255662d75d61574778;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e45fa219543d40e40f88a280f61a93d3e8cd6c16f5b0fd22277c2edd1ebec41f07cd5872fc5b8c67;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f5dc1743cc2b2ebc723db184a045c60116e06f4c62de634595ff2dc0d6a96b01364142fb10508cbf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h190848e523cc5d211635e73f77ba223500add164882d2f47661e46b4a30d890fb5204a0678dedddcb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df4b1a2834d774f649cf671f50f0b99a7d27f5e71b70f22ce9d16af8262f2d6d176fec920285aec8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb539b9c41f607d5cc16e7e32e5c826cd945e7806efb65f424e79182b56039017c008f85ccc8f0e893;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62e6465b1fa4ba3ce6f7b4f1a6523465c44857be6f625590165ecb35dcbed2e6e0c2a4c9db21c52cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f609ea2da60003c6099ba98adbc41c9e41e801ad2770a815d10abfe94941177479f942f80f2aae5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9c977c80201330f667574ea618625806dc8491fc6d96d3e4bbdc7d3090198a069cecb70d4564d6b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb88f61766c6bfacd9b1d5edb606b08b462fd0553a363cb9a985835e36d60b8887b92f5a74a527e373;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ba6a61e959eda371dba6603a2a580136c3f7811e6488bbbf746aaf30ee788d2fd6b54ce97e74d5a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76ef5438e56e14540fc3b2178bafa898a7e07a9dc1e9711c02d9496ce18174975f9333d74d345ac35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddbbeba12bdc0ff40b51ef789059f1feb3b8e7a77718268076e95b3c0cc82554959ec5493336e6826;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h573459ee925ea5eaab12dba25126b334981337ee9d6d7e0c2b5c2e0961f3fad7bf5d37d01257fc43a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha99b98a135ad5e3dcc7153c82797dead1adb5c1787d6d26c7428c1af5408135cbc2bca4c7ea21efc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb371d64508da1d1ef14aa789c3cd1135730fda857cd0810c633638e6d49c1b0d084b69696aa28ce9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb99b76a05fcfc3450de2015371ba3ce08bfb41e7e81fabc5a2d532c601e5e6c398986ab727992443a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcac32b8be0aa176b1d0da08d7e05ba5285418412c7c89bee2e67e278c7730691267cd66b9e799414b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c57353d2db9eb55494a2f4419d4438f916f11b718659bb516d33f823a424a45fa5fb5065377537bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he645d6a824df0e86b824f94934d18178a6867cd4dacb8ea596c697815b546743cd5870e4533d03142;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h815eea2e5ccde0a735080271040144fd8aafabfb1c4ddc6175e995dae2578de6bbf2b319dcc3c06d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4391d1820c0407764e39e3ece39c2fa4b2124234ee187b03d2ee1c079e1bf8156f6abd4566e607580;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15639fbf5799243d62d2500c77f9bdad200fa9fefa07e57b2ff1fef7754e1857bf407b66fc56c22e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf59d44918d4056dc2bf3b9895c51682d1e6044d2c9abcfcd6a60b7a522dee65f15ecc8e7bc15bbd6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c3099bfdf0c1846abb3906f7601733ffea1d6a32de6103fc6a3818314e78c7c0e10f5ee743309e15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75b0ef1876cc7bc23bc9cc07855198c8ce3fb6538b263070fc9d48020f24b0250ec9ef2d1ee924ffa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a90af361735bd657cd1425c6fe0230f841943f030ebe4393ab2ee99e717a9987e924d53c7a525749;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88a5929feefb23114c63d667678d9110bdfcaae64639ea066517094765a9b93fa29980084f97892fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb749caa8d519b27ba6c0e7b855593e8f5233690d3b9230b5c6258e3a53f23d9ed329ee77af8554fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19b7b788105fd60a71175a9743a55fb9fc31ca871a0f6979a24582c110889cf046b1107654bd42e35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe7d3f4ed3a70b1972b2ba141c4344799a7be6f17892e77e798434ef2111a2ce88db91f7265be415;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc339df36d2e0e78a47d1769b198f3cead4dafbb824b1627eac25065923b16f0b1aa4d6f8d04a35d0e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e5293f019343a94e53b72f4ab054a646619262f04c7473f586c6469d4350fc74f639fe70394700a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ad703601ea5854e64e8a1ea0077743b0372ce6ffa3a93fa9ebd5410be434fdf4491b4770f6bd7bd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he927a8fce5483f443e14933005029433253d203c87c2fd2ac88aaf694453daec3982548d2822c559;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a27027e31dd45025091f15af2edeec4836de1c100252e00a5385bc35ee246fd5da6eb62426cf77b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83c7eef75dc6e1b415a9f0596f461cbe90ce0f6feef03658a582089bf5d80084bd5068170e5636beb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h375726ef3f9bc3804961badfbc15ec98ee8e89d72f74f09d35d256031bb92184003f0cabe7e707e9a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbdda273eeb5b3bdad23d215877cb700caaf104fb16ffa1d2a23d8762dd049e5a260f598fc298c779;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fabf152843dc231a3ba689de1d14d15a781652d40c9082e5587d77aeb71a1a6e8b19736d0bcaf1b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6a4b31b9f2a576c649f9821d3d5a4dd43db094efd1846b31238e5bc2703b127fcf0297dfebebd839;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebe000db57be6123f39ba24bdcc5cb3753721207724c105ac6c4b1071fa7f8068e14ab2cda14b1548;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9778c3200ee74c002e9440e650a779d97c74e65cb563bdd77178cf537ce29eef758c0ce056280f352;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83cde5d9b09af100895a87c36aaeeb73a0bea7382d2243fe92b0d803476141d9aad400a1b0fe53945;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75f45f31df06c3b7bf7516c1312dcce170130984ece09b2a8cc2ef4354312acefb77c73cc32517e4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11964dc02b8a9e2f21e864f9c4767daf9fdd82610ee81506ec8fc3823f2f62b2f2e960cc043450d87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cc50338718d90328f5b735c65c5b06556456e6b2ff0a4399e2e77e7cf494b1e117548aab87fa1861;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e8bdf1614fdd475012f8586a6b5f0d229208b08a1a5b5daf311dbc33a598a4dc7b1b1f80ed27dd92;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb770c0d2ddad89e588aab133c2b6987301ee1a14cf71a3140e3ac4ec3f7dce237444365dd3ea15a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cfd34fc81cd65e3e112cd50bc93d5a13e80624289a4d1968fde38d29365ec2ead87e581652c357d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecad5f89e74497b8061be4857ced0ff992bbf03a4e7456937cc8baad41980c459d63b6e4ddb94905c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fcedb4b19062a85d1e0fc23409850f879fce78d2da6c013ae3dea1aa9bc3d626bcb4e9596d9cd7f7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb70b91de2e3f7af5920add224a58528f8d07546ccc3770bdc589d508ef92cfd9162e47b7f9f808062;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9429235511d39127d424ddd576e1911c04ffae127366f91cacfe512e9ba22f6d00b88cf4730a30187;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c3318bf1ba8df108d2b96139ac5d9d1c3f96b6bb20e10bc79e7dc2d0f48453318a0d0d798cbf2caa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb47436775ae2a4374cc280b45d6caba8be0bf188969e0c7feb6c79676a775f4801c6826d3b434800;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b2396b24fe5a27f83d8bef34af0847c82efaba84f8fb110e45a22ab825d5df2cea34854cc60c41d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5eb6d9547586ad3aaac23847c3782a0f06f28da8d72162e054663dc127e0bdabe76eb84ba2886598f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6875f86ecaa66eab974ea3611346dbc2d9f5921206c85cc496f01cb0271f78ed853ae2d6fd5152f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84644ed3ec91a2d552e9f4c1a556f878f1353e391074a4da014f32d6c1fc6a354287da9b9d8bc792d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea3e92d8dd7d33ef1f7fdc2317a267fd0a9c32441ec378e5d122cc2e01c3228111b77e7ef86fdfefd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa8ce3499aedf76f0ca4701db110715d9eb6ce034bea098c8c6c71be4dcb4d1c13f160883472d5e63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h555982d5271c6ca2374eb193c8870dcd1744b7aea0452dd7e43a29877abece451815597e95b417af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha41cd2f30c70a89c699558fb0bf285b9d5cc7b6a15530e841866be8c6dac8aee31a0c783a718c9a3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h874ddfe7fe7325bc524c0b28aa4c90c8a1710adba0c263aa4856ffd1da8431ce855d5a8c2a824e368;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9f3cb26380108127b56aeca0d280669fcd572975a7ba0e9ece7b5b08fd141830722925e1ecde024f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he44c71243f265d74fce84407ca6e042b04cc3faa7ce1e9b617d6ed3bf90166c86a6732cf359fd84fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h647fb16794281c92f06e5881aed3ec6340b4b1d7a789dae8a4af9f74caa8cbbc0fafdec95d63d785d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bc2ccddf90ea73b16d577f8045ee5cfb4fccf9723b86f30faf9ec0fff578cf0aaca04f9a290c42e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bb1334e1e317c33102474acb14f2a613da12b98454223fc7f578092f535ad8d7a44570730356ffd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e585b544838160c5874ba1f3ce899417a04ac74ddad99119141980c5e477c73ec5c441cb59b49560;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1af1dfa13eb21ec35369a608eebc9e8dffe9402794676ce7a3b0f281f05e9587f9760fcdbdbcea74;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha35cf9d4adc71eeda35e63a35c0374a4ea8cbcf857b56a4f9695bfa9879a7c5c6ae4258d142d4749a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb973af7fad69fdc73a1d6a5f7b4dea13536dc917d57ee6e13101136032fc853e120947a57cc42044;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h383b170326dbae0975445937746ac4e719d8907dae689fccccc0e558e062a66a4ea081e5c975faf05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bc99c015a8c94eb49c96f8744f12fed8884938c02b4e26f2b779626fca8e37b119126501f8b074a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35dba1fd9a575dc4a1e983313b45fdd0f9f1ec94444b4bb6f8afbd2872ddd87419237b30eb87bd9fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f43277c961f21a934a8d5f1c3533f0a5c0c20f034793e1c2266ae6132bd85aaab769e7758014cf1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1522714b221d935da413e2611a5a2c908f514c6793de3d1c6dc43848e4440425f9c8235dd0c9ca7dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcdf0987a9af4dfac0e8a5ba7a41cd392a34866bd73ea0c2d70b44dfc2f023b68c1ce98281c439388;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4efc8b03b313338deed435b0e2caf107871ef588d0bfa8e13db64c52124540c6b2ab656ae486f8e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94e5586d9c63c2a3be057e2e6c2bd2ca7ffa9bfc62b319ba27058a8110f87e2710f72b1f7529fb7a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82de3e8ec669f90e51fc19510e671dbaf15cb1eb4a02896af6c683cc26ee804b936dd40d60194d6b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63844e14eeb6a37c6db37abbaa477858ccd74ed586c8a73aeb361af2e1ba348828706f703e93fd169;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98d067d31400e7fb2874e07ecca2fd52c956330baa1815224076f55128be3401437766c06fbb5daca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cc6d0a523e79d22943d3870646c4e2a8febb6e177786333d44c497411ff04b586f0174c25d9e3361;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4795b2d9e86ab2f2aaf7cea9a64949cc45b6db000db069e2aed79891fe028e0b84ae6e2f862c4a8dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8e9bc8428972e53f47efbc57f0bdd2403a682e7d18f2ada6becff7f44e61921ea87813cf38d4bd6f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cf351d918178aa06d8f82a9e97c4820adfe98dfcb0e6c571d866c18ae1e297ddb9290e5411bf48a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97b1aaa84ef25a28c5a92ddf2e7da6e138428e919c056bb96c7e703d8ed3543dd50b3ab2a5736bbb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca49d3d4b8cbdfb1c567a3ddf8ab9eddc9792b1e761c4fa7a2a3376f2c7532f8d78c387142c5b8f0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha55131b0b36289bb8642a89e8b891553ac8bbb985fe6ed9c85758c9085e3a17fa47a37a25c3aae4db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h129285744fda21c54c5f17db888cc010e1c0d4a140aa81c69718d9fcf0108e74278de21b596e4e40e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1633bae2ac512ed1f3ef689bf93ce45880c6368c02d55929e6771a9c76759b2e0b29785843c70d8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a329055bc3625173b446bf06307249a4cb44c018f9f58d768d83f998cb3f42754a6499e2d3bdffde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e05321add980de60eab8721b8cc27fa0cec580c4f4e63b5a1889dee439e50a9f00e9d223fc193082;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h286d3daa9115dceec4718e811688031d5d026b349fb047ba5c9f668e81f7724825a0d0f3ab7adde0e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ef2bfa3974186990f95569f7972553ab11a8b09f6836504a26a8484602e5285abd0c3f31d44d0423;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb00a963cdae3ee153b2ef9ff4a71e03b5a9633c42c3f2c064113a9710918c62a7ddca264fc56b3e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd58685179184e334681bbb936324feb48387dc9e7faae793173c4ddf1a6eb0f60ed9737b5daa9cb1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc420ef90f91130b23358692f1baf2a2d24021ea9d4fbea8e9adf9ada441fdbe22fc9be7ebbaaf2a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2050a33db8cfa70f50079dc5609e9a3ca80fa061ed54874a83f035023ea13081d472ed3ee13523875;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb9ad5f41320a2eaf2c89c4c414de8b134c3d85e9f36bd5ef60c5da1abd9bb4314b65a778185d7281;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefe7cdc1fff041d5924067f05728bf3d3db40dcc319ccd86b32c703bc4a40e46fdc94d6dc5e6ea5de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92719855f02aaadc0dd4d83a1ba0a424fb71109f3a25cbe9185026ec85a9d2a77350b775f757fafda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46f59830b018b678e965e08e269f244183eb6cb0b9dd5e09cd7543cd591e91cc51e879bb42b20d920;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18943c3ab4b6f7566b3accd23000a206681b59f81b960ab6ed6eeb81ee674de875f11dfb82465e805;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51d72335c42ff5f8ceb23670cc566cc9b3bc80348864b041338764beaee4cca40e9bd42a4bd69e1db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc58e068f37814323c75107a671324bbedc149704d1740fd2cfb8cc94eff448373da7d2db94c1ecd8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a7c6b0a693f636fdbb7aa315fba9bd860456ba0be2189fb23ae29a7363c328c1f6d02c612966fc2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1d592c0a5d8dff8fd4a89a3e79064a3ceea7547ef26fb748c4e8399dd7d4c3d90da7ad034a8cd49c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0bd94ba6adcbba1c8690db07e0bd89b36155576e1d9926fc3a247eea248511869756acd1337f7b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23391ffa98582de1496fd08bbe6331ba6b5383736c77f96a5fdbfa786110884af9ceca1524ec48ad4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97277c5baf9a659b43dc95d049404debc7ff68b296570859e6aa115f863f38f71fa98e1d58fc769cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73ba1d7db8df5cc49400b1772e26ed12113a904bef85e74d0c962d4166c66610f611ab1af155a05ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3492945f6ab8683b088f7481c5a0e722e97fbe6eac22f86f175e0c5257fca4a24dafe62cab44868d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h601427abcf19be1beb65cc8b0d69b48f3d00b3e298968ef49cb01dee09a4bb1d5c51951a21ccb1c03;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c1ef1239e0d2d7a64884c2cbc95582bb7a151187c338f33f0c658dd793014926bf5cda277a68435e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a3bceb45fc4d390a435d93628ad68da77d1bc4b85a30eacac89475ce2b33bc75c586c9d55f9da545;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc5ee58b860ed8a4ca5fc89b1c929e08a43657c020584f40a9abaebc023c16581d4d392ab88e3d1c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94f04ca7909017a5e9836a157df0c9636085cebb99d1ecf858206ee8c57903ed4803a67b0e4e1756;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc28d040b1371198364ce825beafa8c081777a490b2008c9039c60fbf818552ebe01df2edde166f1d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7927cbc9604652ae13393d89ca9366d85a3e02d030cdb272f06483b53630df943be2291f178681214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he46c2dda2dc1062a78f5d3e069566080d451ea92d4bbd3ada52984a9bbdbb15639d01f71f8eedf9ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28c7edda12936c511bf868b50e80d1e68bcb8ec6558d4ae3f515707f0a3227023ad954bc1f9f8f6c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dccad17bf41c34fe62efb07558bce8382cdef04365e97502c111fa21be849ca8c3a064d7015ab37c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd94f925e109a715d0b7fb0b713a26ad4229135571228b0d712f7ca1ad45f28315dded369fcc30729;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f77d764fd0b1dd91c156d315526f399ce6029c38c656bc443e4f30086b794fedb6f78ebc888e9c43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1b35f848309e9436501eb76b491973499f0477bc4f5017d9c729372037932795dade49cec0a53f16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cdc01fc486498c3a51f4e98eb6097cb777625d096b75725f3166acc6f17d0cb1eeda5f98a6774bb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16019acc9ee259936f64db5001440c8598dc8dbf21d05322645a62eb29fdb7b798a38944ba9c75347;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66cea1e9c6606302bd44998c27df7ffa09e5e17cc17074ce61a866b2dfcda2dd3efc8c9e4656f06bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5335f08eb8f35eb2567ae37b6c90efa22b24ba4f27b1c2949729254b0b2b04e99453e40cdd4ee30f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb1846a0c9657298442bc7a72c88a228910348a2254146fcece1376c8c8ae2ad95549edbd9f22db8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c0443b293b3952ac901483b7d39fbef4a0dcaf69fdefd0235b52b0f0ca4ab82562bfe351ead14410;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17f2d8be977614d003f2b72ebcf353be05d7cfe62d30f6d694e82cec2090136ea044eeaee0df63009;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c9dd4a0d8765c6928d2c9736a8ecd33998a4d01c4959fab11c7bf461d59e6b1947f4cd743d854dfd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71806ad9c5ceee67915d13adb12000b2ee78c82ee8edd6a54520d977cc00eb5be0cf6ef3b26e60207;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h752a4c60367fa51a7e4e73bd2d8eb900f6cd27a089caac31548a198ee257ee436a54823d224863b0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc05265a7d4b67c5e4656508bb6683369d8622744827dc8f8814bd2d71f68d65a442a3f68ffd378d9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h697af835602127a71b2397593cecc99794af011cc4608d1d53936d42ebcaa605350654990dadc5fd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54dbdea8673fa53aeee89708076e7cde73969e7dec6e2c45b2336b3386d02632be59a1132c82665b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f34f07174b9853787ca16429cdadc9b1f0245906563c080db1443f8591df317de0b98795d4ff8ae8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83dfa75e1f1852f833eaa541a78ef282db73a46c6e9555ad5972212c0d2bf6223b96db0c29d062038;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f54ee95c119ebcb9e4e8ff95e5332f7b0758a2408e280b75d146e3739b677cdf8d8ad0c86292bd44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff98edfffd86d3597738fb79806fa3c1661fa03bc9dbedc8db7c190aff053b52ab83964547bd83e49;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a1ef265698f30d59409a36451232e004a30b73e0a15f129bf83af84ec8155dc1d6b2cd98be9a6b56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h535402b8e56d3b94ea1a98f0834dbffefd5d3ea6ba85138a6483329841c5d884f6f578d01c0405340;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac370dfb28bfce94bec204986dcd1d7266500927b5f48beae5898e57f396e3954ee561cd2f31d0069;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f3f47d333321b68f6609deddd48457532793b4a324fdc175722304eac9544399eb9b5d793bec2da0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22dcdfcb4ad380f1f5cf1a2a25d5a89f0f29b46040ea56807a3960c194ac2d6f40b5b140e9190ba87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h766ca0165dfc9e2610d267ff2468be5db82a99621caf98e1c70487f1e4ae8b8a65a16d51494971626;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcac9d37281d5b584be892a475e9ae7afe312827733d0f81feb1b67dbc5d1676b7ccbb7c6a01a8971a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fbe2ed14e3e70fecdbbc7a887eea74bb367e0394cfc789da2bf450f28504eb38664f50509d0bb8a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c79998aac9cb856fd5f66221a098bd312f2e4b2fae69587f2cfcb621b44b7be1fb6a5c2add1b74e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ffb65a5eb03bb4c27a0afa61f5ba4ebb384cc84196b441d1bca36dcf51e49b14ed2d4b48e2661edb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bd00215cc1881f7de39952093a052c86944387e863d2968d7bbc853a74c37a5357222eb02d5c5a89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h521ea45dd0ce969644bdff593e13d96994447234e680bda2f9a2575029da8f7b9a5d91dfc65f41967;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15cf57f1118bbad9dfc68a7d772ea6e897e8a6f0e75a8ebeeb1f7eaf099809c5eb1a97566dbceca0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17f15cae2a97b7fae9531785ec2cfd0346092c9e9856dfafbbd26325f646074b107102f333776081d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h924f37edae80065275a78285c1afda81d51e9d05d0640dd095fb7e6c9e81cee15495fa9cdcb60637e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14b76088647ab2605b3756c6d2b8534e2b239d6227080c04d2daf07cc6f2924d5b93e2bf55227bcb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h514a7e0c6bb73d729ad795df98df3455886fd507f18cbda4200cc79f2e83a3d9483895c4b58ae1d04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90804a3951750bb60a44d0c0aba0307283aa0fd5b2d6a5d0c08547a6363217c838544bb7adaa1b68b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22284e928dfb01a7273483b5b41dbb909c4bebde93c8cd55f1ab92190bcd83057f3c5ae78dcf8107b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc99514aa1515358c577f16d906e3ccfec3a604e9bce9d0071de6ec38b764dca0e14bf459698c1a76d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4a7111f34e5cbb5d9e004a3183be28305a24d2cc7f8add7edc66be67352683e695d25729f5766192;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h660323595b12f8d0fb41802bfdb563da1effcafed6b18909bd1f87a81c0e27efa9bdd17bc71f53775;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3d21d33321f4700e3cce00d3808e5eee172b2a50fde47785d6bbe2b464f8b8e5cd0cdd0521eafa87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf8cd0dac6807e7f435450c88df62c88c0090ff022e5d5a7e1a348cd578b7780d43269c83e20283db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd838e3322e740b15cc2a819556c0405a02f7098315ad79f1cee1b878cd3d9ba21d0a256f2fc3bbd7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78ca8e0c1b6091f3fba45d5c106721a876a0eff219ee81c068e6037048bc74574d2df6e42b7021498;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56308ba6bcb3d0cb7f1d7776755f2faac9e1960d19ccc7375f97fde40c7c4e5985ea8de233ceb04d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8767a82d90612ded8e942248b01c8a8ef55179ab857740fda80e445c00ac9358004185ec95ff8ebc0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf49364212135795db1029a7aed39dd47783f4b31524e99dce7f3cadfff9320113f265422a70a0401f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1f06d165d7b34bde37f9bf0fa82b01d6bbacb008b7a7f356346d95dd16321f69f611249350bd1204;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h251af5ad5ae522ec7aa136cbc0965940e4cbf079f1740f5b85d6d88a07fa4995336898738e64530cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93272f041211eef9dd9f342ede5dfcb68b5c888966bc797a23ed314cb9d7861642fdd7bf0d43c35dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hface9a85354ed68b4a00e9ae4e3373be3f7e7c4386518436b911cfe72a807105422726dd74f17101b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha70c559c88918151b5d4d61baa5d65d478b8256f52e581e626acec1c94b97c49014d5722a353e18f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c3b02ea2198bff35a2ee3a3532c460186f98a36a2e0b55ef7061c34b69459394c8539521aaeae708;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefaa513b2a09c193f87ca41c70ef5381b584593e52c759125c8a42d7043710f2044ba2542e36f8c48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6976e892f255fc7571bc962c5201f8aaa15a168b0e3c64d1b3b754d9334647f1240bd2122819886f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4a41590b9f8cc2e9c1d11d8e60cf6b548278451392217e7322c1fce7c21423ca0510bd28cbec854e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9850a9bcbe4357f71f217f60428548d9e937cd48b80395ffd178364c06501533663e13bea88472409;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h193287c92efb46a03d197c1d69b6bd9c32e1c5ae0c1438a6e6d6634bafa2310cea1eba56e5d2cc2d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce667456ce67d0811c6e0c0babd87580abd9e3bb096f01ddde1207011539015a0d33161fca4919d97;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f0d2b99780b0151a478bd4a09a92af77d35596cfba6ee9ff268dc3c352f53d2b5fa0d70e372baad4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha427bcd91ec1fb47f9172d3f68f4ef09d941e2c98210ea7063fcf895e098ee0ed96d0ea5e94ff6c62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92c82aae40fd5e43921f91e8a6ab17114c25ce777714d915d91a361c74525155dcdafef125bd230b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h782813e6c5a347f2c82b7bc6b59963b86c238ce4367a347ac0cdce775117f9422d09ca99208f4b7b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2d76ca492218d2e96a7cf16fd6a5c00e6122255a1445bf59b17fde47b8f1e7f13d291a9a1c4b3d50;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h156ad241aeb02b5ce7b1aad30b77b2bb7b71356db0e2395cd2dcaa0458c422c413efc1dd1abcfd57f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf24b78cc5f430f79ab4eb920df333fa124c33de16baa92273defc391f0284b315384a4a86e610a3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca122f637555acdfef26b246828df6bd4f5fe0d434a2050224dff9dcb7c1e61629e1610a6bc19a145;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6653aab0650ccd8bb9663bd217ff2a3f6cffdb0f2b202f058c44af75d71ddfd625d09859c46287b7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c19f2a87e2500abe9aec79c127fa9474a8b4e7f8c982f44db21a4181ce089e3e750311e87305f2bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf567e8292382eb01b613ab41a043af80964c087fed970487afacfc1563cb751b40e9c4800017be3cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h435b6d2023dd258e7ea1831e3bed7cf083df637022343583c40228ff713fd48128e6068237d89b31e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h283e003277877725e9a429d365babe955b526f93c21cfde92d6cd7b663f4391ed9e78e8f2e00aac99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb3e1b7decc6752f0e10db3799c2b09c91f8e809eff137e18616809797c66adcf6ea199dc6d06b35b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac37f1fd57250c18cee40fd4cda673e5e912f0e75e3390d46563be5d31a46a23808b970cb933b670c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f4ecc4d02cedff6d611984b8d7addc7e28508ef58acb3ab512d33b34cc076c887637e99e45f7d503;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a46fe73160abe30fb956af45eec9ca773947f6eb5eacf838daeda93beb93d2313d0cee23a973359e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67b12430a4d344ef8d49bed094ffe0f93675478297822725669fea028b62ca78549cb58a9e64750c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h927e73ff83d564c0ec5cc403a09317b33dd27df3ccbef438ab64e7ce1b17ce583e4c297de83d8dcd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0daf7a45ab486243419ff8348548545f90cf39929200150c48fb38f40267287a96bc79b2ce803152;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12d54bd0e0af7a1ec6902374c6b95f544447a745e0664e305a85a9b1895a4fd7425f72849986c9921;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32b318d34a8a8c9c9bc83ed30ced70f5ffc690ac108e19682f1184c6644c6da1d5392e5e12a6481b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc41b3299188268b1e5901345db5de56e9705f81fb6c62905b5de333051f25306019d010eda0ccbca7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc008f123e5f6d094b207648c5501a8983003fa8d599b9ad09780e069f7ac4fdbf5d7479b3c0ca8a50;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44f0eda98399a7cc37f030e47d1f606eee81810969877aaa6c5c9479bd3d4643d91ed68d76b3df8ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63be0fae3470db0bb2ce07d850dadcf0ca7e78ebe1c5f64312d46fdc4d09aeaad253b9b13b8cc2dcb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95f17994481b542d35781b2d3507fdba3d935c87c701f9f2aa5fcf10b502d61b3331df4cb62d69b66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80e4a0ff1d765424033fa1305d2c9f8707afc6198a332852b778daeb5e3addf7bdf1b86eb42ae0ed4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b275b60625bf659febf92e58ae13951eddf123f2cdc9431a620632668e218498fa803e7bb08de4bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d61082a1159c1a1860b46f270c239476414928078a9807cae96311bde317aee7ff0c74f127feabeb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he74b9b989caefdca39955e153a4d60e260a281b179a51ce8b516f6eedac5db03a2712b0c5c56f29bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dd19290ffdfd82977a68b60223700f2fcaa9c8da8e35572a3ce01d75f8b686c8abd872570dc6889f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2010ca826aad1993eb49577289abc45ac7d1ef2d1a1943b0b7fd285e4747a073aea7cf479503a76e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95f9278685b15266da0b75d84e03eb238a35d81b2bad7f1e688524c419688e0123d727d5073e7f7a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6566dc806306a86d41a2cca37710e9b9aa2c449c4ddf037b3ce816735efac9826ade2836f1683bee0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54dc4d6e649b901228b2e2aa6da4f94c5e2c57e294190e7c254a5e494a99676d7a3b2c2ec1b642961;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddd441bcfb17650f12fba1fab271c97f78c30c4f6de83a66d3fca4882bfefdd1137b09817f3ca3914;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha14fcf3566e4592c3f9c6979aaad994da8d4260cc2b2773ae0909a2f9e2565e62f948261c99aa4884;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5920f83982d28e41de4b68dfdb90bfbffd9742b9ed66794724cccf38613d38d130b5ef0082b40a940;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36feaec5662785dbf31976ee512310038e4ebddb5bd9d9a2166cb18f40288e262dcc9546c617f1443;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72b38b35c3992fe1473d36ff2ffee8fa09578c939eebedd05d57d521cb57d5f953167a90961de1b35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h794be86e21c2fe2f46c2e4b1da5adc47c131da8bedcf5f1ba43b2019439a9011d5418daa746ca5f58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffb897429dfa5b47080fef140b5ebd3e7c9102a25f16caf9911eec99d5651651f2ab8301af49cc61a;
        #1
        $finish();
    end
endmodule
