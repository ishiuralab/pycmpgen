module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [22:0] src24;
    reg [21:0] src25;
    reg [20:0] src26;
    reg [19:0] src27;
    reg [18:0] src28;
    reg [17:0] src29;
    reg [16:0] src30;
    reg [15:0] src31;
    reg [14:0] src32;
    reg [13:0] src33;
    reg [12:0] src34;
    reg [11:0] src35;
    reg [10:0] src36;
    reg [9:0] src37;
    reg [8:0] src38;
    reg [7:0] src39;
    reg [6:0] src40;
    reg [5:0] src41;
    reg [4:0] src42;
    reg [3:0] src43;
    reg [2:0] src44;
    reg [1:0] src45;
    reg [0:0] src46;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [47:0] srcsum;
    wire [47:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3])<<43) + ((src44[0] + src44[1] + src44[2])<<44) + ((src45[0] + src45[1])<<45) + ((src46[0])<<46);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccebfc6e2050aa128fc338977540d5afc1be39eadae8438af868b2da0a7736e4d3ca9ff4b38cd5df6083d7cd09d9f6f225531a7099671e1867d5753cb5d95e8581e78a61ba3aaa76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb7cf27524281e22b1d976b930fdbcfb57ed772c280cdcae9aaf0f8732f4250f2c1c24ea9d31122743fac49f09db3068b7110aad7e82bc6ea7a6741d41cedcdc3b13662ef573176;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde1696810eae6a27c94b558a973cb2e27763410e723cbf0775c656a2edea65679f60ad704a8ee6d03f04a5eb6a2a919ad221297b84e3255573148939957c0d6b768709c658592bbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3565555fe642368ebf68dca430d8c248832e52571dd9b638592c70e5db8f02e2ce4e9e03318d2a7c8638ef701d2ea94220f785d5ac55004ded9d1198ac17196d939c9b984bbf4292;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d16ebde9676abc0d144a6ef026a0cac44fab764937b2009226e8279471c61ffc7a2d21aae4a381bbc8b977fad458c68f7b6cb4ffec955d9dea12dde57472ef9dad932cce01c2cd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf902da991d94c87929006d019ab72c0a5ded3bc4e4fe39bdc936ded6488416dd7555021cb4ced1d4ed2327aac2e7637089f16009b592b7d0f01dbf8d7f2a386f5a1b52cdc3143057;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc882eebaa3c954520c5bdd9e6f7552041a1a66a4766470665be8d9a8bea23ce94e5ce50835c5ea96b87dc98294c697468490adf891fcadf91298d65336e30e6e0b4e210e4427206c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2567fbb9f71c9fd97e8869a8c7a18712dc510af9a0862cf328549bd65932964716faa78cdbc551b65604158db279bd3f999230c05e9002ab6ef7753c36f6139f0b43280fa244c513;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b6bd11f10fcedaf9c0edcdfef828f6942dcc3b5c35018cc0d7869f7c53d00ed0f3f5b990e4a9ac4db47b0341cc44b869b741af884eac14de7ef9877523eada1d395d43e15c16ec2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1964a2ee7e81ade3571d1dc7661d01713f5194f3ec4ddc93682d2342196de4982a25476cd71c19543f1f5b07c3fb1b6517be605a3eccae9f589ca4067376cd905d5eda8dbbac782b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefa2c78f701ad2ec77b56f02fab977dbf231241341cff17482405b059ca056851333242aab53f8b10d8bc11fcd4164c346c3f2f0b5c8969f8908c1fae54add7801e5825c4fa3b507;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39c110c465fe10ce6784738a07a13f23fa242ff5c38a5d25d17c78ce9aa6c710eb34360a36f572631893266f8dfbde160b346b103e2dcb19dda0dd0ca8d62e44d8db8165dad8bff8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74efde655580ef3c3b5703b31a06a35641edc4a02975e6faf64a3d34cd72e1e00c72e957ff949de14a58693215be8eee70aa492503c1bf84ea1091c5ca9a8bb21c3c9714934d3d6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4257cac7fcf13fe217752ce43ddc8488c6bcd3f633bf62fc8a6dd1433d75b8820237c872b7390640b9e915d5b220dfed1496e4efe1d9a5a093f6d50decdf7978d182b2872c165e35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64c9401b8ce541ca988b5a604ba205b3dac01cfbb3d5903c4376f0092e9af0c2eca024c07429cd5e98528dd5a08566603932cdf37073cabb53cebb9791f95ede717e6b9f9413ac27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cc4979b31abf0bfdf2127abf453969854e2ae0a7f5f2c5e703542a70a96582368efc2163d4afb547e8ec73264b9f5c1f11f2fc36e1715c2ae9e9b3922b5a2bcafa8ce60931d4667;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebaf0bd6abba38bc299e5b0e682109b33b93295aa80a210376af28f5b681c0c0ec40c94fdc4360d0693099770bdc19428b61474c18e40542a94f4394726a4e848bc83adacf14e0a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h262dc59c0c69aec689b0af23ba7bda4af61604d0b06a4b89371a42ef2c9a814195960271bdc8445cfa80b6072e469642602eff6dcaf037a18594d74c8f13097670684b8ef13cc381;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8464b662734e39974fe1df5a26011dadcfdbb6a23d91b6009322b2b8998dddb9702c7bb4ad9bb79e4913fce5bbd68896661cfb003a8c4f1290134311fbc779c084e9ee7becd7068;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e8b93e45cb8ca48dbd70bc8709388777b664e7d0ccf6d7c84baa16824490477c112d4115d81066d58794f612044545779bbd06f5eb04be8e2a824b2f66b014e617d5d3b4c38efee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78e1b448a982da7639dca6b9899071f0f187d0ca4a4d956c0b4cea99bfc24a5267d58a417b54aeb0e3f5bcaf02740289d9000dafbc824851fee444ae04ca10b091cccb1ce9a290f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdb56fed924404c4a9821454ca11328e69ca19160c75b5f419e3162465ce47b009061497b2747c37ff4a1e672baa1e26bd03b17b4e9ec9e2d75eddccc8301405218597e935ce36a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd6783c8145fabf990136e89d1b10a673749b8d1d39567d1d02bc3a9ab9305bb3c169d4e801a311b1c7c2c8fd08eca3e46762f7a7393f6c288fdf6ae17ff7fc4e7b58336a958d30c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda7e29e295a356103bb3d1e00f6188d451348d5a19cc6c9f596ed1235f46c52354b5b6f5ec87832d57dec5a4ca38f3dfc81291205d682e5daa90bf161aa97417a9eae31d1ae528f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8abdc2d170c80faea801821295845da9f50504c833a73777b6fe6d7d947293cf70b9161a15c1509e90ee16a8109f12f0066e211fb547687ef866916df98b9fc43af3e7345a13decd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8577d5d86ce1aaaa3c45de4b09a63fee08ae5b5dcbca5655043a1002fe2bfa78e754ec24660580e19cc943dba66e06094838a27d184d1cfd82504028b4d120082e3d2affdbfadedc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ca532858dbb0bd481788192250f85827d402af481fd4da5927e7889f90943df6291557560b6dc997c35b94ba97e177481483551ec851e24e5fb3d65c03793fda9fcf7d642e6f923;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h534befffb64ee4b29ac3502644b1afc2d07a35b78cf3de3f69551a3a77415631a28e7df58d63c1d4bba7e7b64dc2234bd4df9d01fd62e5571376788107f005f20d0304ba78be74b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90bfbb976c6ac6ef1769e392364c23e3e82b7df35d054bd037de1ba91bb8cf48f62e3f8e060086158e630bb85c23472b0a5d6ae120034649ed61e82abb15fc9e71764ebdd962ad66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f901e4293f63b054758aa1fef039d97db64e2ec738240a51bf4bbd30e692aa8e9d66fb0a98c33ed92e2a45eafe0ac9b5e9b7f52e52b2f979c3716739a68e27b4737cffd44247780;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h895939ecdac3fa98e8a2bb3b18e60dffd9513925b1a94270093e6490dd45e4a814b3e55d78ddd342d3842bf19e4ec0b5be7f10250ee4c241517b55e34a6eea7c6aea752936e7871f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dc7393b82cc3f2730f7f6ad40fcadd479578a4bfb3041d10c8b329f35611f130beb9e8301b2feb2f34778e89e31b2d5767755fb64293c814f218209bba2adc69db7bef1ae7a0a1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h990a68d21a5cb65a1bb5639d0ea4ca26275b8d9c2ed8d656c085ff7617f995328cfde35e5f52837597e264163042ccd8d2ce25feeffc9a5d58ca897d4346df6f5f4cb0682e781a12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a4f2cbae87646bbfdb0394c507548cbed17fb5a2d1f21187734963f313b083a2b47240857d4138512a79776b1a37f28d3fab28bd4acc391ed6043e1f739781e1ad72fe1f2829c54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86fd47c39d9be9ccedcf6892d7836a5f85dea13844a5581c150d200d0a6934a8af161c6b3636f1fb4364c0b5c42912ce4c992812255ab9d6fc32f419631dd137c8ec7e4c176971f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfba729c08678e6bef279ab569e8d5ac469a11beacbf4f081983a9239516112ce67d49578e5c1b2f1116c923c93a7b22eff5ac306f19d91161fd606b6e6fe4fea7d7e11d2bd435fe9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6494ee38f856134981297bc0771935e439c8fc760edeffd2ca3b0297424c468d8cb072547c995441aafd082bd4d8ba2f1c8030dd07b7228b71561dcf83db51eea2e6a777bf20db8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f8a5c1e8f704d4c8ebc038a56f9f3a11fea096336a51a3e9ef62db47e6ef44183eaa2e15798fa67158fb758e655f017e43b1acabd89b97aaca71dcf57ecbae7c3423b74cab7e20b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had6c20acb13366aaf4508cb54b2cd22c8acd9db2d6ef43df53db4d7cc6a92bb7997b354774d8d2e10d06ac3c62e7763b968a22d8413964a71ecd260e5158ba3490d5605b976b562d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32d4a79a7140f8bce13205db1b6e52fa71f9a0f617fac3aba71d4761a7ade58fc4dfe6f06e1d529d47b0df23eeb5439836fb8e56686a3f66d5e64d3893c2db5dbf0d9feccc52c0d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90dcf16092845177e9698be37712452b356d9dd5fd8c2af58378f1acaaad42b2856b872aea6012980e074fcbee65f7e153c6dab21031d4f89eff30a68325b4c0c9b000425f8df298;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a664eeee437c00635120fc5361ec923eff0a7bf8f5cf6cb4fdf1479d1d4f7dbb0ad3bc73c3c1b30c1de2e0f182dee99c6f5bd2cd36665cc2aeeda4163765bc3b3a3053c1defc166;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ed4abae4bb5c97ce67f822e19e4c3541190d4379c8d0e0e2ac76033c4c4a86e5ed3cabb5db47593d7da71ae7565d4866817dd479d7a4bb131262d1068102b9476cd184763f154e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0b24d2a9dff7483636a88ae69989887bf5e694c251f9e5f0e89781ea1d64998c85535a5c46d272e84b0ed1b0e014aeab340abc808b4e81d8b3db9e8e4c1a6dcee458b06c8317c9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50a073ea24094468f4e17145dbb18c7f26ff1c01f4e3582902765803d516bd1490af759217db9939c4e6c1d4c32203b7c02f37152dcb58dc8a5696866cdb57aaa34a0ee43dc826d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec3ebebb75d46b530e1dc988349737044bd7758d205aa7ef7947fd2046ff1d098a751e8fa08e408ec381ef39e941297b5e3c0a1633f886e58fd5eef02ea88ec8640ff3a6ff28817a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb619540c98c5cd2aa5c8dc7760358794ac4f4fd47d6778ed1968635531e8bcac89005ec1667307622b33b40e5edc6d2d5313826fb933fc78861f2215ae328ea43c05c8bcda6644a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76e410202007ff7c4509c92b5112c11e5283da9d877903a31aa85a0e2eef5d04afc4df538f510a43d46812f429df449dcd3c644749057e8edbaae0a0e2288348e8ab9a5009632e3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa6a6caf6b1fed1b0e18d3771bf9c424fc26689a1294aca30fef81e1396aaadbf6635f59deefc1f5c102c889b86b433fc28a4f8fcd8ddb2a4e7ed5c3906be50f515b0db914073d19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8f1299b01980db348b64d779655530b0284dd79c85b31669341ea5922af3e582f0dabafd54b9962a3fa453dda602cdcc086ddd25e4f6f75c265fe1c4468b1fb2f018b460d8ceb73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd052feed0f82a8d836a156354b75d436bd2cfb46a298d1be1f759cc489bd5fe6b30f57e809ca5f0cff85fc4a855054862ddd65283356c122f5935908578ee5615129361523316a5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bc94e4cbc2d5d682cb8c58d92cd025fbd2cf29dfe5de96c33c08a2be30d930603afcc4b050c3a66c8bf5fab507a818d75a1543427bdd0146d2c812d02372fe33908c1faaf6fa36b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdfa11e7eb9e25dace03df687082a86ea23de2ce20715c109d3e37149a87eeae9627d5976bb112cce7ef7647754859f0bb6d31aac572a9d3ee19eaa430ccf58ad33483581c204323;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a8d0d5e8b8076815e835fa50fda62ade8b9c4bf354465cfb774b300e1ff7c176ca50d22bda84252e40971a73edfe4549f22fa21a7033e081fe0c53012ad5f72bd75027c2cd45ffd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h391e2dc5cfd3633ddd1f7305430f0abf929a9d7dd147bd80c82db9a29ae08e68e7c4b64c4656839509f60cd98203290b887cc9109591b523ddd33dad4bf7f68af9250b337de4011e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31fc028f767dbc01f60632657f566cbc09ff3cf140cb39ab741e5f8562379d8b4b00fc2a5acde8a17aa0e860c1544169340055b72642b2082887af7de2d3dd266b3f214ed9f50246;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bc4b7b24c1535032310cf4e1c70fcbe72ceff74cf1003209755bc4ce7ada23c94d846813c9452f0f52eb64ebeadae8e9b362f21dad6e43d5aca088ecdb03f85f09c18c432530616;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7803c22b95748a5122b7a0f7efea73cfa8e983e916645ebe6a83bc768a28e993872b09537fc60448fb4936178c0b069fbc098fe0111edaa2dac59acc2cae14985e1964032800c475;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h214be3ab5794da9621c4d102c5a3f4165389bfc7b08d7c40c75e240e94d3d591006021d0610b525e38eee76b6fbfc41f9fc67922135f0fa6e534c22ed0151f1b6b5261c5ebbe8d49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c26e6f6eab439d2077b414802e05f437715b00ef38bb20cebbbaea4cdddb2d47261c38bdb2702bd32608f3900796bf2e23810a8508ff2978a4152d9c490c45778e5c56178d2996b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdfbc6fca1a7d9633b55f9cd3a6916e24f9f5e26ae87f7aba10f6d7b436327416a4bc6943442c0b33654c8bd6b9c303a1c1034074494a36b6ed286eed2a795b3f85e610e85d95e16;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93939ab55b3c8f4e51e444bf99d1df6f5d6e9a344d9d8c6190a18554f98eac2c49960012378593808b823fbdd4a4520a4db0c8478f16f39fc6380063db2f99d884439ed86ada11e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1842a4fcca432ddd158f755d3708cc77f370f10ea5b1759457098faca056c2b88c318fbf9855c03282cd8d53cce82a82fb8017ade8b3a5175f3d73f4274b605847540beec474c92e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a5b1c92e548fbf07116a06e02bc66e34c1787f6ae8b4b5459cbf9fced3f1c3e19a03ad6a4033187ebfb9e8cb698fc87643aa0e346b02e8325b5f4f862874e86a9c4e7990e22b781;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4645c6333709595fc8dca4517096dee6dedc70996544b1bb68014fa6b5674345f1b675adc29f132494acc54409576104c669c8132ee455032ef2dbb1919129260473c4700966214d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c056662cb2e03539deda67ebfaafa96c1d1e595ce561359a59f152df97f30b43ad9955925f6f7bbfc3b7a582921704204005153a2221f51658d998cbdc918c7a666eb36c18171bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4dd742b8bb4233d5659fbeecbddb59d2c7d1bcf18650c512bdd5cd808f29fdc02a189b50850f168560a1b5f1a4df5fea839f50e9b3219e60aa2dced4a67cbb25fb01dc1be8dce3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcd6508ab63f7cbd14510442cad46c518c92ac08dbfd10e24fcdf273322189a82fc252d397d9713c1efc770c05e537b2a9d2603e5793b5eae2beb1d1ed2776ef679c40e855308bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h562da4dc6e7be652a70befe46c784c5f4e33b9be134306e5446757c57d6bef9d983f078adfd611d423a49bbafddf058b4e4729e687b91031aeb185131f266ca648b0afa40e6ee6d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80560d2372ba8470bd053aa6685b074e44b7ee75b185165d90eba1e3843f155e13a80879015b483208259ec1216b72b0cd71ac5e39b9a1823a8a17b8270da95e61e6b3ba308189a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc371fbaa987a2a7386e9efd38999fcdc513e9ec1b97a1f70b38d5b6562109b22cdc0e9d5f7c40b1b2b73303a7bddaff99744e09bfa58e6fa9772a88a4c049664ccb22c3cc10b475;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4047017d5e9292c23818559eb4c7fdc7298cb09b6eab94d46be890ba5ce6f5740c82789bcd2116a5f6e600bb36dd115f488b1cd0366026c62fce562345d18e7c01decd51252b5a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5be4c07bad5ff74d8880de1dd0119f02cc9cd98a9591900c224154b457ed8d2eb7c290d946e42b04e1fe73668c06e1890207b53fe140acb9ec19b1a8e1d71c537466a32dcf8afa1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82b72513436770151fc9fef83d34054753a5afd3cfb1922b5a869768f86a32bb1e0c7423fe719a10c96c43ffda70028df445b033048ae3c7b13dcae7c00cb77090e5e767d15a23a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h995c194a07963aeb46ba030dd897510938eb3f3442908d684ce780fea399b3c02477bf03613b1fba8723e0d70d9d6b7da0f86b579af806b676df6de5377d18ea920128f564765b14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3587222daebd657ceaebca24df54dcf550828946f98cec023f14ffde6587366254e87a0a9d8f24b9cdc4514f740bb5f231b1b2b2c27da17192d29d913d0bd021d329589b9d92a82;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b1d36c90dbf7dd3e2969a9adf76ce16e8cb25514ca2965b908b3246a0cf37f99ebf5e0592a9433602fe9f3a2fcffd4e626ab45fe225ab71a4dfe3a009a238c928dca4e390fc3b63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a3bf050bc2980a7adc34a52c9d60008db843f01872d027c7fadd018f0386de4df7720f417bcba6678f0cc462ad079989eaf3d28c364e1dfc25d84c023f335499ba7bea542289fd8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33825375794871f711db268dc017587841b07d15d693b94b621737e9e42490cf64e998ea23462c88018d4bdac0090d1e7da9b8290acc689258c3d639525487506106a52b19b86dca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf71ec649b49f3e6cf0ccb3b1d46e9c086445314323ba11f172777ebbf83282179d8a76288e685c81e12ddea6895c4a494dc7f20bd4bb4c11aad5611c9e5d89ff20d038cdb003c5c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc74338be9cfa8a133bfdf04c137f061f226e4ac7c955f95eb6bed8771e1cceee6916f8f25598ef52f02dca5f18144f3e88057e15f5b36a2fdada03e2b0bde9f444cf93f912e8010;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae8b94ad0795d70569781fec10cd547e280f50fcb6b7276c993e2838b9772ae2659b755c49e9afc3b62d1c0f33ae6a6fc807756a4c04a20dc6fd566021398425002aa6910df55f67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h365863af829034f5f91d76c409ae6d3f3bd5c13bd14d7979a4c9956e0b66c95119cf2fe47b6ae9cd4857c4bf320f7d97f55fa44fb3c077b17bc573622daf86e7002b50a54e59f042;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h110276afa3d80a30b7c97b246e39ea3f05297b6365ab4047e473286fc320c5f5ede01bd8089d5960897945375a06849fb4bd37cafd5662ef48e11d7c635b4a2e7176c248469a2e39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26654348ab584c47e0daf204a2513a6c30b8d921bf13fe98f4f68ee0e03861c44fce3455c44aa6c7f06997bd68fe38352b6a97d36df1339dcd350b3d98e4b7f6e8371d3fe7495332;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92d8ac17c152ddbe721117580d869b77a404858b8b6bc375063a36dcf75b1f17361c01e519679ed1b820848029979f823dffd1489495d78ae487ac82d5cc40030024c40618f07c73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85be009c5f82d804ad7d476194b1e3542b9e999be9631c086d9c17d48b1fdc8244053baba71a741396fad932bfac3e3ccb928e3e72c81f8040e6d6bd7c36d3a01f879878e78775df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd97d81d3ef4af7ddd137ba49413e442187e4eb09f4c410fa5d6140bb295334141772970a7752daa17874866111025ff0dadc3ef4735e55f2484ea86da641da2935142354129a5788;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72323e789d001bac3b6a61319ae6132b3e3ba2d3bce224dee75790ad71d193208478cbab45d43268dbfeb974cb54d823a6ceb30f89140ca6e86d57e0b7284383873e474de0877326;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd903511ed11dfdd2116327da7c9cada4a76046d9129b1dc91ddfe49266458882387331149accbd8d149d0d5cea05d3f56c3de64e73bc6e297563ccbfec2370f65e21283cf4b73029;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9030709294632a6ea448aaeee1551e7296da6b4cdfdea9b29294cf044ab692da903198a84d64ca37d0fbce8d0bbb6b6dd3614d34f3748118faa479ed79b3b01ce77135fa281bd06f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7ff7fa93d76625c7241fc1d71ac7a0373424ae6248ddfc63ad9b6c52b67e78df3a2d8ed5c52c547689e2e45db7613a4e20f3f5467065bac844f71295a914ce1c1d97773b20da210;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafaddcf393c9a6ec310cb11af2960deb322f2e050bb1c505bd17ab15331211a27d477a0123d8f704c27a638e9af3bc8fdc7663f95d71061db604e9bc861ec5f327f16c03d037a1cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b011f5517fc3031899b10a88e9d411d139044a80c4d9d82ef098205b5d1cba92f8015e4a6d95c4b76f7b0fc99b3333ae1fa4f5dd6f7545cb454cb417e04786dc67a67d277b2f345;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ea6b351cd3816da38aa6eb0616c085d137baf0ef8604337826c2b42114c9986687842e22ffc737581bf3ccf9940737536f09d6e8ac2a074052c72c20591d8f7c6aeeb1052a0b2ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h330c6373e0b34bae918457f30ee8af99f32d65737740abbcd11443c51a475bb4aebe324e0295c8e89b2f7a510cacf220dbc051d15314c8a5c74957dec854037d2e25d0a28e9969a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6472fd9ae262e52bed2e8380d7909f818eb4799887989c1178a62320cf35259c6d799b37253a180464a5d2fc02bc9a303e9731fee7c6210f6b9b8784b662f233574e4f1a266776f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8f1baddaab568c7c88c00eb0c3e54be5923e91385e4e8d68fd295d5f7c80e416d244501f0b3b76923933c380cd480a8fefb74868f2669666d9ac9f250962d920b1f6e3f6f8cf6b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2da4995f598280f6b0c996ba523342c69dcaca6a0458446b3ae6dd8da3f130d73c2d41d0985e698fccc1a15908179ca7d696acd09b62f1e5b7b711c5418d13580c7110d646f4f534;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b1b5b557705a62a348425880ebf55c7191051835c4ba431226b797603860565d212b9be9df872ac8ae7f7a1ab9c0dc76b322df4bab4ca4ff62b273478a7bee825fba83a8e3b6855;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd74ee6fc9dda524f047c6e9af6a1b213fb525ac54d72fc5d556c6d51bd11dba3bbf99a6b14af636a1307e8d02eadd70fd8c2617bc25aa6e97e7558a3fafbb461da6f1236bbc29f16;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72757983ecda5cde66627f8366745b532b421c94ec499cc4b98a4cc9e12c94d253336369031f30cec7240834c8be2f1733f9d07fd7d30b1cfdf4eb6a30f4e428582d1fe6ad514274;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb182e31b0dcdec0eb8eeec7c5fbca6da9396df9d627ef27c49a1274ae44eae4cf85d94f1a7d5dc806dd56738fbfe2a56c023c09b5d002f572d929c64800a18431e18b6b536c478c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c5c4eb6f9835e8c39c58a2caafa209271cca7c6b47d07a7273eee975ba3a595a0999566cedbe4828741e2698dd245db36149257c376353a21f0ddb39f1003f20a16d44b5a3f2136;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd29a7f24c808e8f4d7fc0651ac633dd42046d96c9875c9325ad7ae4dc9c8bd1da0a3e0bb297bd7e52386949505c5f4791c765953498d747ccea38806f58ec38a68ec48987db7caae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3039b0a3e121b6f5a47c4cc208483e29f9b4a6a197d16d64f45961f8dcae37197fca745bad86baa2cdbf2a884f66e76f7b4c524929c321412ab092f8a11284ed1ddff0d21c325d04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d724fe88fb7fc0215bc64fbdab492bbd4ec476cb3aeb924b506c748724df11344e531ae94109790691eb515f6d0a4aef0be6a6ce9f2962963e1eabd28a4448f8be181cdedcad40;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a7fcb1a5f3538bd563cfad2f2a17a88c7c143b3b9d9e964558c50472fee0b774e554962395277be3cfa2eeb9c4167a679f0424230e78579010f466f82c8d219a12d596a4aafb278;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dc1a8ed2a6755f1458e19a3b12175459d41cfeec76aae09b6d0497239cc42bfc10aa535ff29b2e8df54a31bd0417194993dac6b0784818bc227017b458d5e12c3dd78a6f1d1bbfa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74178c7c17221f1bce72d1cec910906b306282a14168984ef4929e2b13349213a33fec4595f77cb15382f5e977f2059d9718b59aa624ef84f41c269e928fedffded893b9659fb399;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h751611bab365a1438fa361775b417c438af2353fb2be8f1a5ee6a6d82517a1fd10751ec2ef6cad0e1566ccf403d65146e3d6db18ead0a6ada3791d9796e935c21a1985b14e20de19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ceed2c0e82f08c1ac64ac2a1dccb58e9d5276a011e2b3c56f4cb96b87af6d2bc7134265b087061ef3ee6546147ed43d5ab8f1f86e7d512b0d078c6ba5513197dcf848d8813955f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9650c586ff9683c25dd71fbe2d022da50c438c7ba6da375b4c0f7ece937e1d5b0e6f2c0b4d1de6779747bb9e6b40f7001c443aa78d40ee007b799aa4f260efb9fd942be5d7ee832;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c06573dbcdfe461e68b450a34b5f972a5be867b6a4a58b41e2c98d802895e8adf09cdd3c603f64455ecbea8d503ac5d8efc1edd6430fc4f23f067a3578c2711a40e504f5fa261c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h785bcead2fb48e83fb4afea8370ba85429ad57b8bea568560d4969bac729339f43eec26080a88ba449f0455fdf8b48c470ae92cc1346b955b180cbbcdbbf58364cfc54dbbe9c3328;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aa98af78d19872af87878fde2ba06b0778cc6a257bd3d01adec70ed9579b129387e94ef7e8db052dd6aeb776af839e42c8c683c426b463d700758d26957bb779a5bd18dc2c2b39f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he67613376c4395c989bd8306f42f4b606998da91020e751c452c4905c1879896ba42f8222deeedf99b71d57a2b0ba99f30f3320443242046bad9f9c463b49924730b8f3c489da476;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca94c49ddd5bf4c469640693322329687bcbaa436b218c7f298ae7ed2cbb3eef29801953ad47253bc27384a8d6db34da0ea38010f86aba71699eab2138a1061a90cb2c03642b98c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2208d7b1b5964d561f65d6239f8d4219ec5a93048e8622eaf18d5739586a6d0b15dbbc4d1278226a0c0b7f10076ffcb2f17cce101e1fb43756f76ce7abb31d89120e722d17d5e5aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha883f71473b2ab8c09a07f4b2ef7c18e7da4ffbe84e62c11ff2a0862d4c1e5bef9af29c0de28ae0f14ca9b89ebf886e3b29b664050c538cbf6bd0658e3c5b0e05a5f46e98ae826d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4e495beb10943c975fa31e04f439814241609a5d893e822dc37407c2e64f8c7202f291db84d8ae17631909c4e37c16d565e06716627b68dc76b91b66494438c591bb410d7d232aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8509a21d247997df3216b599f31d020ecf003b7dc3aa779c1408c92d3814f12a81262b60cb42718d7271c34d643e1c0688066fe1691ef75e7d7d9aadf9b85a71f8d261da89f33c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf0541ca078fc32d6d6b71d4721c70a4764c8f70eea66a6f3fe837522f04dc0fcce36ed755461cbd97c07ab80b612b561aba17582d87e8c1415371e13806e8738463219d60059613;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7838ce10291c6f45b1ba18e71a945add2bd8e1e0fbb0fd59eb0d08fb9f547bd371bdb7e6cb5a3d7ff78c13794d665f31138e9d20088f0af8c14299ade51e39510144f59c0b02b5f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f73c12a617e6a5c4535a11e3c9830163ab75fb7a80130487e1e8a55044252325a7bef6bcb59f9312742bccba04802aaae6403a176da6e156b0276080f7d888b63dae67a58178c37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed1653b6a340c9158f4eb5082c4f6c6b8022a3780c4cfc0b7858aa12960dc7446c21d521109af8aa52f54bbfb20b504b654f27501943d1c9796f2efa94696a1720a4d3f9142d16ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h552e7dc93726335593608b615ae2eef92adcf5c0b6cea3d64769f7028e4802a31e61d4667c89bf51f5557c17be36ce3f7bcceb84fe5593179a7a68b247b357d661fa50447ff14f61;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cf0d39b981479af2a7044ba928798561fe0bb39813b66b95157d047a622c83d1809fc9fcdc4f4cb9c9fcb223392927daa2745551199298df48bb3b4ee04d4383c5c73f67c728500;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bf7e87c01aeaa1e04ab26f3e5a69c89ae92a5317e952d4b8a557229876ffe00cae0a4787f21de5bec432c017f9276a62730777b33dcbefad680a686b6b503b509ceeebc8946aa45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha349a3c5934b71c8fc237573c0c2f8ad7c97f76236b3ac5c983ea4b1c45208e00e080acf470307e16173b24fe4d81bc3847262d46b3cd0425b6ce19dcb57700b4f937d36fac2b2d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12092b33d0f3cc9e5d66e4bb46443c77d5beca56ecd7c9c9f79ed3e9d1e8609e0d445d33ee44f65e2505993801109defda997c9b0c79367ac039efb3f2f8be76fb2436e26012bf47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h361c7220b89e8a456a85a4781b131047375e9932f9a8b42d19016defb523d1bfeb5d69b11c9c310768542cfb7698659478e47fc006fda5f2092db5945460af7c881e39ea53c753b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7d9e3166228fc75f1ee00561bae745f0dfa6ed2d66bc5bb337e669e76c24d8a9f6354bec692641227435e44229a471fc0d2c498ad8986e6883769872bc38057ff1db42bd8e3297e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bda138b0bd7f54b71d8d5e4e3f307aecc12471c9d4e565be9753266274c238accfb6d8f90fbc141582ae1b989306bdb3991e9521bb59a8068a5f76475b4c68d440588f39b1f12f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b8433acc37016b3478e734703f13c4b5b872863a8f639e8e35cce06ce70472bf3d6000fa028521ba90dbdcad470dc56c47e82d3f873856d1596d4de0cbbb3379a52c541fdcef260;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8556265dd939acf196e54d1b369c52a58b20552f149fef22c12a75530139abfd30f5b98541161352d42d895fb80eba26d5c6029da9b480a81f3db85f7e6bccf59524e19414ea6b0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16ad72bc6a1f4b5ef8c6b64f4c66eb1fe02b462522690763f6fc00eaef57f93ef8cc720fecd122ddea21428b9745a0249b54bd5b388f20eba07fccc03cbc164030c7497aed203674;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd713645649146ffb27f1eafd922c5ce7b93720bd474766d7d77f526cf9910bb36dc55b83670c38430a874ae9ee73b22e31b6f7a2978275a5e466e411c64fd103d7f52f97a0ee46eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he443094666eebff91ae6c4af9b8de85942c714d6d08b5a3e2ff1ad8c9a7c504ecb4d0742aa921756fc20cc239e62b9cb6ca5978520522473e722d7d19963c3d5bf6d398fe89ece7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d371a94e42ad092bffa4e31b50558a99c45635d24c33f0074c23add620a99c65af2bbfb8bf4c5616b33cf3bb67d897dc0b9ac0a5ede4a59d7bc339e1280b5e659c92a67565d5e75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a1206b5f4d41f448152aa86ad599008ec3ba690a74e171e55010023d5c22a51797531a70a0bad2816ad295e826c83bc8d5d17517424c6415079f16c78931b59be482df85bf98867;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5799d9da08cfbac3e70901366abbc4d5a089a2b158b0600b2fd2829f6be74018f83351bb199ea1a394f3b21f414ec6612bd62f0967052e7801b16bb0f46484983ef280fe4ddc2c19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30957accf262f47b017974474e804cd15676211c19b526d314d751842258756c64495aad0129da2e5bd9111cc9d0550a778f1e7da35c9e506bd60018e0af371d50a95455222aa6b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89d9dfe39515d1791c2a80fa9d47a07d12c4732bd53259e57d61f2386102e9ef6ecd62886f9c941d5db58ea152ea86507e61deb4e3df756a7bc3b348c3654987e6d91abe2141b50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3cc94511dc6c2d1ef0c5e3b7293dc281209b170d6ec1d404eaa73de014bfe779a33c730c3d34bdb171b0823673c19cdfabb24ba4c1c7128b140ca15a45b201563d802dc5994a9dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffc8b316285f1c714c78fd52683b6bee3bf0d48704e33f11b53558cdfbb501b4d5ea94997606832b982adc9405188eb5ae1721a9aa0a9f9e89372b422b622dd101e8e28c368a387e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53dba668cd02d60ea905866a981e2b29f2fbf8d7ca6d84e4d976542f9094f2ca1a59a22ffdf8f5b135d917ff5ef493615da26702215b552323883fd887b99b4c9c92c12c88ac5b1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf1158219d18b176782f5d29a31c45668ff1705dde251bbf173af4528b16fa91dc5b21118f56fb2c98fb44fc975a4b0c991df9c51d7d3f72186bb43c6330afd530f05aa8181e4254;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74996993ee8ada36b9b34e3fa6e39f7a24e2c98da048f25f8f17e921744fbc74058a75d8bfae1e076671b29ad131c87d36cb38ca418098662b10a621bc2477991db35d390e07ae69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbbe009662dff7c1f1c4a8dfb8d760f97b544120d15e928c70fbc24e38382f9e2688703f6c3d9953d831120e78a98493f9dc02fc41d4101f6356726ce546dbb22911b0af830f2e4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58683370e66232afa65eb76826fc725c9201b52da5e83ab9d52c1a50b4841bea62ce7bf90d8c86c11bae0001c5b96a80311307b7e1d1f1edf5b1aefcc5d23a72e3fb2080964458ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10917f5f44ae01bfc62964a2e6d76db7b7c525b639107712cad4d398dda5556e7c2f789e5b1a8922577b77469b21a6d8d3d0ad9a9207e24bbdf39cd51621938b6196879a05e0235d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c9b0bae730b56a6a4c06538f833086b78b13d97072fcabdb8920d764f9ce3d22a955344add7ccdd957938851d0b079267e5ad2cb1d4e1fa6b0cccc80ec296f19cd7cc38ad5e2653;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98f413b8a8eeba9066e8410489fbe7978b010dbeafb4b4f4c0a445df6f1ecbc1ae68759d9776ad6d443098ed0d6e781f6cc3aa0275810c43c4ece513e0055909bed9637e982731e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf8402cb79043e584a32a59af89ec32c3a98e0863ee259e5d4515e9b819f215e4afd082b4bc7010c06e52a24c2ec61dc6524eeb9947c721ef867720347481397dd65809f64d6b9da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e0fe1e976da4dcc4b04f58f6c14e106cd4424a95bfed7da1893c9a603d622b1f5c2acf5b1a33e8cbec4bdea6365189ed778885dedc6e31ea0032549c24a1dfdc43ba7b00e00001e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60881d476093f1b2c998f25d978b041844cbb47d089a8347b3738b7195111de24c2043ac90b405366adb00eb800a374a27aca02f8ee43e84ba9d5005efdf429658320f5149e8883a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h950d0ce0c413738b38af1ec53f58d1af23f947c86d5cd2ab68520d4d19b4a5b1d767f107db3ab54eebcd99c0ebd2082e5361149d6f1c727e9806537386c059f63e8132df5896c7bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a3545b11917358825c29730359144dc29cc83336f8a2b79cc26d5149736bde548f1dcc42461b49a3d8f0ea007a8bf0c8fce9b7a36bd9fac222eb794fa19cf1ebd360d47cc210091;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h723e18085d14e9f6437bc8ab3705f50d666ae57c05783be197e6189526b087d77f224a5bb11715a155a67cbfddc5e0617c1cc14a8192e53411b95476b59ac69cf97655546c2cda87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he34f86cf284d7bae5ada18aa67b274c8a043070c709b54e6c2b85f66992757dd0f01d5085772e217e794dbc1b06b2521b4883904520b679efc4460507060ffa0f8fecde2e5a73212;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf198ea6216b5892e0a67e1e766ccd4471ad0c77b9d1ceb0474d437534d87a4d5bd5e38c9063c64ed3e591c4c09efe69c222c8bad877539b384070c7f4ef807ecd9d09ec0d09a2e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb4f9b76dc7d7531c11d41059e97a794b0f67b0d0fe1aa221ae536c2f873402aa89eafaaaa81522940ea0c4e1e29c7fbb64ea18ccbf5a2d892a62b67ff32bda62957514fa3cd80bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf28a04fa2b903c7c30be986fd38134c69af026a8e63c1cfc555592570501060dc463b6e11ea1a0cca3bdb124d78a5603ef6b2363b99d71e507188c0df499fd4471be7e673086580;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdcc513f373d5dab6dad69dd1900a8d89bb294d5605ffec748675fea33359cafb2149d40798f5f584bb20912f29a23b5fa28386c17f9d714e90680f1abcc2b8c736e0ed2447d851d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc87698487f3da4bc1c178a19055835481ec70afc34cf23e05f5c3cbfbd4eefe3c1d94e50c1f28588c0e8e89d2eb7fa00091bcee65cb549fe0bda92a4f90b8f9db73e48177b2b5b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3c988238a94f60cf163538699f981f19c06abc36bad75d838894592f3f18f5c5410e6323d66833d82f41a67056d637315ca321d872883abb898dbdc84444b6714eb484541761ddd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ba10f5f5912b8a43e31d8f679bf46f255cbcf4cc514deda40190966131180ed255cc0906d994481da721d25ac42604741d5dadaa77989475858f1090ffa8ee7601ee84aa7ca4ae5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d351c654f02fc242ecb7d60da2a469d11874bc209dcaf79e3318ab7a2491f0508d9f4dbdfd64ee417a394f35bcfb86b69be604dcf2334e2f7c7b6cbf0f7969dab1f9bf28b6bb8dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb84406db379fabc30b1d2a83b54fbbc09e0f38301b06318aae71dce546622d97b6937330ffd92446ef886cd49b5e5943d63290572807c31f30d260c30d0d9d05ac6725badd8d2429;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5254b587dfb98d42aeb3f3de12d736c854b352e9c8596824cab30ed41bd72cbcde55d826ce03386139993c052d4c59812055ce74ff26655517d5a2ede25b1fb6446ca0b5077f1a9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73d8c39f46153ce4fd414908ba5cccebabf72821c133eb0eb22dec5f4a3828c7360940fdf1e3e0cfc30234d2cbcea91eb57513b7d24ba9a0b723250f81a0fbf9e7a422f55edf22b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4896c83966be3a63e9b6ed616324782751f9a02eb97fa1e11cbbf9712bddad93b952bbd6647ae701d77adbab7be95dffb6b5ccdaae889358fbf92640ef7c0f45d97e66c3b9862c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5afe08357d792f169ceaf6cbf9e9e9778e8c0964e09cd6ac4e305a22597822a33d598055abb0dfa57712312845805de47696b59b127f76f9a464c9cda4ae60cd13abb0ca1e52fdb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f70eeb9415bdbe3818e5e4113c39f295837490fb5d99bde33f6005fb88c9a9f29b76f731e4e33193a7ef14230804c378ee7cee329f711d668769cd76d980306fa88a3768bf9df37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52716086800f9094c08557017c8f83abdaac0d8e774bfa907060229427aeb3a6ed7cfb0da96b095e87b655e039c9cdb658329331c1cf029b35bceaaa67c89307d3faa2bc264315eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8245d24433546ac1deb2d70c1a44594a191187e6cef7651bed234905bb2cc040b037dfcc1df856a51a0b4d9cb384346b4fb1cd083ad108f187b268121aabdb2b9f1930fb771d70ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76e260adbf354230a663608693681caa8403c00b98ef1f0e1032c6bcf660f468ab23ba41594acb46fdf48592ae1d189c6846531edd2822c549e855a70b92e349559089fbb36fff33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17dc5ec805cf9257e0b3ed704bd48761dd809a919caef35059ff5a426e10056c3663afab964c91b9e117f6743fe18f603aea83e1ac53bc59c237d65aa2c0555992dcc170740f7311;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha888f277eb950166baf2ebf7286d2c4f2160372d9cba92a48251f46dee548120d5538110cd042a84c151ab7b70de396ef93c60ba5ee82535b7bf89088736579f8ddb87054b3100ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h134e6b6c28cc5ffde7ac7164312807b8ec0382f2cdae00336ca0ad2bcbaac5b891d2037bb6097d997c0fac6f325e2163cd33f932d25b5cae38bd44c71f00ee1b6af3d42720f01782;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haec46652c5e9a544d9534bf1fbcf1765057abbf09a2bac9d7267ba49e6fe747f9f543d8d88d7250ff1aee556534cb06f57c2df9668ae86021ee9452def27b745783a7b41034e4764;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89b05386c8d4af3fb5bc174336168f4f62846a96447203d199650463e13be0ba059d6d510ee56335a4558acb7a8224a2eeb466c07af5b8990d1028b16c0bf5069406b3dbf52ce7e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c8f725b3a5e640c7c813d1eae5e45e2035014850e5d54dd95253b8bf7c8cdaf0e37a6a3f472adf4d46345f5f8b336b0d3ccdc8e17a3619a7bdd96b42f36b6bd810a467d2ee781b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31bf69b40aadbecd0282f8ce67e84d6c30ae99d81c43e4a6be366e0d70092901e9f5a217ffa71771669a81a5cfebc93463f9346fcba9b33c004afaf333832943e39f8711a622828c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h120e6dafecdbda0c001539b32c16ca9b3b6661a3552a7ddf0c0a190c2e2eed96b7d41b7327055b88c1bf05a593300d1f506d829b29cc24dd15cf1c04b8fab01e4b09b176abdc1665;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb60f482588cc1df7ab37c808ae6eb5df00b4e73910a7cf0a2e8a9bd85da767ee68b4523af42928d7d44c7ba327bfe2ed27a297a81b0050ccfee3798fba7d97911c34aa2f73efb0c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde71e5faf2f783d9402a2e19f5d420ff00bd78774dd7e4dd10ec3eec13955a5ffddac35b32d88e71084117e33c835b90799de535bc9a4d5f31a45ac8ed5a777cc6ccd532b82e0c25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h130f9521ff59a2158b6ef8b4746beda040c31e2b95028ad717d6ccfff4791415b3442c39eb0f6a68cc7aa8b3f56a896d4435be53c785d693632942d0c86acc071ffb5768bea3e400;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5549f536b0f164d1ddf5f53e2470c65dda492f9cebcf2835166630d6b45e993d4e31fb0b351f2fff76a98430b41937eb1fc466d028d12d669962c1e290e27b85116a870e8a683215;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2567ecec98eb6febd4dde0312aa017144ce9b5132f03573939e30fc26f94631825cb7f30c87b1ce94164766898ab36904baa9ad3e9ff43a8cf6ee22d5e51d6a5b0624db818673e04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb64f42b1ae4a502369db328316596d24dff1fe53dafc36777a460c65ba7ea8039cff2f0e6197e31c0e1b5a2aa5b6994d812eaf00059d09a5fdae6a70628eaee84fd2c30bd7c84768;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a3c19514b2318c67d8498038a39ad4f8be7484dcd013df985ed3a9ec315bf221cf2720b29085af2487aca126a235ca2fb065661a0b033746ae338ddd3da4032115678679b5ba0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aff4287cda1ce82cd618a42bd46cd0792e05b19294ac79a6d71a9ae9464c2f52ee36bc8d0b0072c682dbc8959a786699140273df2b38727d35ef335a8378631f495f230d6c0af30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf88336dd925429c400b383778df4c8bcca73bfea7a3972dfe706f8d93ab0b23dcbbec17dac0a0683b496dd65781160bb85f54fa895158cb16e9d1432a77ac05ee0e4cdf5894f984d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d4ba355bc74a99a46e277a95c21d5253495f8a51f763d42cbf5024e05577f6b5ae212ed4f7e2da038b5f0ff4620335ee6e2735ab709b649fcc5a7321806d0d4894e61caba6b22cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he309d0bb65593d2d404cccf89f032508d132853df47e77eb5e1ec5f2f613b74e8a9d0bc65378ae5ff0e5fca6ce6ae7a66e598aaacef6440610c5bb457e2a9f15724d2968d3ec28a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29f376e80309a2b7b9dd6d609478581943748e38b409a6028941fd6be491032b0decad98d8780c4ac740d0ac14a7d3a6c324dff5d9b4caa8878287b77665fd4c27ee10a84907c91d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fb7475e751f1ce902012f1fd6e9e3fbb2f60ba73eb607c5df2cee8cef54b08a53ac76540b2a79b7252f26548a008755ef2b66333d10d9e3fba12253015bb6333e568fc64b095e90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aded73055e103766cbf350270969972c81973c4de7b10671a29f543ced406c2b528dc6cc04efc07031dba6e0a0056abb600ff6994de6f9cd768563f9eafe8153f9dc0544e9fdbf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4c02350ec7d0f361c4a9741f0733bf6ba9ea60dc330c33ee6efdaecbd1c01370acda5bfc9efc78d999c56872a5e5bd29f66cabae07337f989da90f95782205a454537441dfadc38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4207512d8055f4b2b1b650d785e0008b86556c6e2bdacb0685e40889cb698fb2c842b91556683ffbae780ed4d70a20ef2df4016a21072af0b442ca0f9ba411b9f4bd9e0a44fffb25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1b6243784b8a3b03400154c1e553115ed1ee36b231089d525aad84b8a51408fb2bb1a557c1cf9611b16b90ad43bdffd8c3191c125a74dc27f5988b675cab86b58b5712440236e59;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h208daecccf32b9c899087b0194015819e6d16e3ece9e896a83e283b06cb019e41d7b02fc7e80b1fc38d4795b3a94e651bffe024d86b123128c06d98436622b7d5d56b9c708247153;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h682073d189c0bca35a91a0a7f4c5357266fc737c1cf84818594af834ccd3b96ed76c5298cac71edae39600f1ed4b688ca57976de15607dfe1f93b320ae2f03962bae166de8cc78a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d48807586de02585d0e0237d979b7bf042c96ff4232aff89f3cac64a3525e0d628353f8599af268b919dc13cdff229a6864a0f731020c3a3e81dc74d8d9418ab07bfb772e893102;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95d363f1a7c58c328f26ad0a32cf462d862d1ec937ff72fb2e508045cc075a14e92af410791058486dc85beed2d440e8b9bc3dd11d60e0886c464f941e7f848660403bb7ce85bfad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1cb0513c1d3c336f7da06512a8fef2eda24bd6769026c7d1d8ba5a323d560591c9d97708fb079f0f674a97f77112e39bbbfdabe250cf4e44f112bb4a3fd3c1c6cb1d58fcd926d5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c203485602202c9615ef5e6b246b9353c05627a7012e8e66c33d594fabb041500f3fce29cbd872ee0de30595d670e417ad9751cd60eca9615de7947fdd3fc6b15c57a0a3918bdf9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2412ea36caf10b965fc1d19dd58c0b22ebf845e2065cda7eafa6693d434e3bebf2d73551e6dd0cf16df89b59dfcf28f79b604ef431c40293ac6f9c61fd923e147e10c2b12549ea8a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f0851eedfd9e00129ed4593d72bc2ae89739fc6c66f1b5961a076fd9ab16faefa3d85519e95d41e607097754349655b5d2b266516c8d749fc089735403182a77c3b3062a8c8ef3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb868200438571763c850268fc12dcbae5a9e452d96f597e7f625ecabe4634d599d3adc129e8544b36108749082f2517e572bc7309e87e0829d3ba75e7b95e7cbca0f5dc6a433bcc5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8910708920425c9e4e393763fcee55ae27783081e861589242e45359c711482fa8769a58b5e1b87041e96604f50447f5949a14be819125b873c75718e470b38c56a392b83e07ce61;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50411f94148a540113963e50d916b1c31efd0aa450064811dc5d96bb0ed3988689dbacaed1f75a539e0b069d21bd7bfbd44e71ac5df6f86924b3523ea1150dd2b86ceffb2f359bd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a32f45e223b24bb17885b3b76efaadefc84bb91a7152f79c3e943cd8fd45e6a136c6e2dbad062c3b56d75c7e095701f841bb2867f09c38bb66b843860d1ea256a053f9481865b49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bd53131972444e3a98f0ba3c293cdf05a3fcb66f5619b8474418817e8b6c589fb8e13b1bff74fa562d800cb13bf28dbd7d55150bcc13e464bf2d51a4a25f5d5f7f2254d5269f8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha41c389152162e9089ed3f9f5224772610db18783fc013d484f740485a2da95528082d27dec1bf68dbb12d203f0829bf40f514aa77481e35f9180808c4e3f8ea75f1c12779e08897;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3764a27ba715b4a7f150d597adf6eca4b9abb4b21f1944c443a4cc468cf2ba885e6ebee75c99d7bff520156ddbba53effc6c1c806e72334ece84cf0c1b62b6089c2e018e24c9b694;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h483b138be6b7f9cbbcdfc4e3f7f2b0cf95022e6e0e55e1c13dab9bfe0c898f952a4a46b8cc3b9225729946b9b44fc501a7a46d73bdbb7d4b32d3de1212df7b1c9229c715e7ae3b12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaf509b62f16cad4837008a36afd493ea072b76211504866d21e2995e677962ea7e5280229eec36e70230f7c6e6533492ef1a50c4574e13383905269a43059f2bbe0c943cee376d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h309c01bcd381b6829a68a9dfe69e0d9583852f6a0d234fdea4879ae8e3781f1bd2018519e438b80086477bc611bbccf3805d01ba1e2f819a365c5272e1b21916d9df9ed85579ccde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h261d6e5697d6ad3761ecdb18f76656b94621b8e0f123ab06eefabd99c7911453b816b6940ceca3737900bdc1796fb14cb63ad9f9cac3b392615557c2a25c7b0720ad525b61bc3c29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3e63276130d8d5a767b0e82b465c94081e804832f2d26db504fc94dadb8f32b573399eecd69052e50a9f63279cc3d2bd191ee770590964ad7a759f3863921acee43baa2f6125ba1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c47a1e10146d545ff5cccaaa7628e6b0121f4e4d162af5997fdcd23d9a41033f685706a7ef8d43269832332d0e40313c636c3bf4750a1746b727874f823e76e9cb2f74cc11e2d58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h280bb7c96ced97e4fa49ecbb4e2260a267f4036507c41e6787b365567257f1840af978cdc136cdac61632feb2153c72509d6808b20686a3b05d7787437b4aa1cbd30df93ccbc2ed2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aee7e0f1392593f031d086d244677c9c6b4a919cc7a80a3977646eb743386397c272f369b92c0f21c5f3dd350932297d1e3203feabb2ea525d859b9c2912dd033a1640cd0e711c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6189f3c9f6ff8d5aa628f284585f497486719415f806fd8170920d1423e46b7d1008cecabc8a681beddd9f504eda2a7b919a769088f371e76154f376d887eb631cdc27385ba42104;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had23c9cdfb5fa9c0a7b37a767b7ebe41c3ae77f6965301536c88f908831dc13489538d6cfd2a85c716d01ad4d063fae748982689b59789fe846d6f5da809b7d5ed9e46c55f0952b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd23f026f5984cea2a037ca7d83a1623ba0afc2e9c17013111c390518b536ea577e4cd00d51078e7cb3d4023d37219d508c942967c3f8a3780a071e2576854dd3a7ce40d2eeb6dff8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fe50b5af9ce0b4c8adff7b9c029461459f5eee71cb67324b161ce4bcaeb5f8ecff62eb72d6c191d222bafd8fe6f3a23bd9665422531fd9c8be6e8a52456c1f282766df0f54f207e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc53e7cdc3191ad57fa472cf7aaa83cc123f3518a2b0fc0d9e268a569b3d6086055615feb6344f0e8cd9c746c7b9d8c2e73261bb1172c44a1be56440ac75e518d598f61ed4c02e984;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha722a1dcb3c164dec859e0fadc5a75539a64cc821ee87fb2a3fd04aa47e9aafb2e8f6af8cfba60c430154f751eca2d197b7ccb9eef607d438274c2e44bb61ac71f941597d7cdd0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1367c96f8b05da289b3b1dbd088912bb0e3f1ff711f841f68cbbf36cc1eb1e481ef911ed080d1adbdf9cdd63da30862a6e20e54d58097e99500f2e0fc97b9b0d9a3dbd41c62cc2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22ab3afe11410801e81e1e0f96d81a13f81ce9ee8b518211fb78a167d2f0565f2103b58bebe9412a5193c65e26005059aa6a96c606546bf13c27c6ac68878137287fb9c1ef441944;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc196f3f570207d5c6840435a33bebf91ef2db24a3eef99efdf35aab21310582f65788798b802ba6f8965084f7d357c8a8e43b7eb59460458efb34e43883d665936a5c6dd3bcbe4e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf83eb04c447b743fbee757597054cde4f01f667224c7c6bfbf5a1398b84be4689c71473018c81a615a25c49bd09f8ff52ee8aa80db62d8fbe757b662ae9622ccb15fc30d1b03d043;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5ac3382db7e794f056bae3cc059e26f8801f0293430c0073383fe853dba1e429282855dbfd3ddf81c7e29802ace02c85249c2ce655329a8edbe7391b06656e45e2eaf6d8cd93603;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f5c510ead5133effbb68b13ee938f76d1d208eb3bed2d9b49ab2349eba12d87d16d5c16a4e6f24f146444311ffbc7d2b999364d24de3733e2065a4426c652963a91e5e89b39167f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a6396aa12f9931241df8e4e479852572ee01cd38be79b31cfb5adc87e8c940f2eb842e2d5c34cdc887e8191cbd63e60fce5c9a29c07cf5d172e0cc9bf1a59c299a8f4bf96454403;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h470f10de7858a130ddcfd45d6b75740b0c8067e9c325348f755d7cc6e1b1d6c0daa3a84e78091ccbd34314947c818a9b5cad1a4254f45a98a69e4193bfbfa8fb24b1eec57443b79e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb314a89ccb0611cdbf49a237f19f1bfd8f15351b0850ac4ea130005222f4bd1265d3426d4576a04e4fb040390c3aefcb36c2f8a9d7fc5afad4d4071d916d4733a1df13238b7bad5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf34a84ee093b52e08debdfec9e2cc8ecf0157ce31041513f5233eda8d2b1a6936c61c5a4a47476953d1b4ac54e0764c7b80c5e6fc086a5a1c4cdbd118c661784ad7f46235590ca9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d5f169c26b860e8e75b538f312082f4577e19fede5620bcd86f3ad47d7b78a04feda083c888e8e0bf154504c8a61ae085a1c7e87a90c01f5c88679d3d71679a065484a4957a2b9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d73a48268111ef837d85a4830fe4e64346caad32c10f899e1601aee74fe94d86ad6152e49d812bcd299ac7e724ae98de46155cc01dc4113392d1245d34482635e09de03f4fafa27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f75a6a003a53a115aafc613ceaa398cc5cb4b6083ba778af39988b48ca5ed8f291200c7cce71c3ed0f1c86129cd1a2f6f76be36329037cd4aa82ff743dbb2dbc6659373625ae4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha80f41191e57c32603aae8e9f0740f5263ee622d88f9a17f9f06b8907194b2e63ad2c908125968f91f1a2c642ce01ea4d8453ea992a372915bae03dc44380aefbc44dce678c70ae5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1493d0a64488be878c4c6aa472b9f84bb45e94009f5f5c7e2034c17131a0157afc4f91570e51d098d1bb880fef66c62d813e7fc032e975ed6e41e3b8b31d84f6c210dc7cf552ee77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4eff3e3017e6185ab01d02285bf558673319cfd99a6d38e487b74f9fd15de9a71603af0c5325365bf2b820438d436f9082dcc7ac4d35fb65119ef7da5487ac5e4a9edce9238b772;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab5b89c7fd2d1f4bb958f7b86772f2e3bcd7638bebdea618a96a59d64318b35d2cca6bfd115017c2e12b90b20e2153593a220fc0d9bd9ffd7e46719f1aa6d134c24b79617973ece7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a52933db5b959d9e3f5a069a3d544e7c742cfad87ce6ee675e4e27814b4f5dc45aed144ff11005e8f0471dc431876cbf3fed8614e31c3609adc873aaba53f2d7839159444c4ec59;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3692889b10b6c0ca7262c1638b75ec43b4803720d54d26c52162d30f37753da1a0452a030fa21da10e7e87f4f7ad65dc30126b165d791feb29fde64679b908e335c2dd47bf1ddd0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1046dc73e9578a2476f155c3f7bb7b66405c8313bee34c7f2e1921169d950fe851209d20e178c5140137dce647605404d4d8a49de89b8a09ce8fa77db4d07c75e59258019edc41d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h448c5aa30aac4a1bf79752ed42413ac609109c1249fae526a5a9d945939f00baec901eab3ff9b5417805462ffd3aeee29ea546f5855a471cbe09404e84d1c831b7ddad26804e2b46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e05920e99f2a6bea8f53e068317f5fcc8773347e811f6275a477848b4606534a71691d17aa3629e65ca2ffcc335bf0b1b0b063c06a630da0b08168d0e9551f4003873464ca744d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fda134530947be2efed11aedf41f3d4d20e8d80cbd1e6fe52311060b9eadbbba3335514301ead7052cc78e3f9788a7667751aefd0c050af99d884c879958e9e04158830ba603b4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25b92d5cf1205d97ddc4a4e4b300f9fe89dc04b96f784da9d0dae43b70cbf2b86249ccfb2dd966c2f7a4f1bd4b6a40719425dd052883ad3da9e0b3db7cb41503269737e6c7401fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f8085f1475d0303b7516f17cac7127a0ee2e7dae9ab7c1636c0f02a4a5bc6aec314acd438bc428a51a44f4d0bcbd2c49a582034c319f971781f55964166f9cc72e14614cc49fce0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd75cbb19250ea74797019b2fddcdf08a371a2676714a9544b4e121fef546803d32351f2e719188a83762fb32c2b9f3e8fc46392f91022e93e4b8f92bec6295ca2f6a1215671b9f59;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6826a626a7494328194c729b5ba0800d7887a1bf05730acf9dca694ecc7b10a608ef3154ff40b83d651df0f2573bd66e36930973b727144a707a7357e2ed15303346648eb18692d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4c01fd1ed688f26c993d6e492de1642cc41c3d25a7f03e2c3570a2ae34db87f18319d60f784cd37764a0b7bd4c79287f99daa6a09ee3b7f50cce868ca9d21c6aa99e197e1ea54a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed9c1e1e383331b0c30c0091b160672353422f7e93feddcc14622080faaa01d721b30305ee358e6b5db5d6fc178bc47a95e523a8ff4c9e9d1bc14eb3984fad822f500cb6f2f2f122;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82e4f3728b967a4b41eed9c1519cb5bdfe38a169215a53e8663856fc3fb6dbed52d3a7010e4bff5155e2e912d3e8ba1702d03c7a4c087acc925ade921125b767ac1822cdc49d14ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1327e64c0f9c27b55a02aecf1e53d0554bd38a05d6c2d5dbc11bd04b0dace49f6b014bae0220e6bf622b60b1b06347b26e351ee962c06341fe65d33a5f1b0170b7913878efce3e1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11e63dfe3243e36725933ce7486c79d7144820703438f0349d09944721515d46023d66b682a107f24f7185d7000edd7380224f773776a38307e70649cc0bb5d0a2766b286c040a47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb1f719eab234d0947f94302b48d509ccba26b41d76c661a9e269de349115e0fb130f39a719e4c843b4c059972f333bbdc04b9202184074cb9d1f17a305d53ae51d7672a0af0adb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbe13c62b853cf239f18f0bde3c1c6ca128af4054323335c661c30381d3ef9bf074f262966a3f59e9f62e3b6d3f8c0e643724ed274e469c82fe9f2e3fa5d209016c143e55590a36f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8611073421d24e3ba6f048f030aa69220811cd009529a49f0546df77863e4718f6c3fb2163ef64d77fef4cbbd52a71c71c7a9ac6b56aca325d0d8a7556ecdbaec28a7224d784bc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0db8b0e615c63d3d3f4159d1df1ab916dec73f675ca9bf965b9a7a042b1f502a6baa0263d2cb309de2d6c221d66db479b941c692a1ca473ac448ab9dfbd5e5c3486fcb321eec707;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h523f96612762ff94ed5ef468a4d8c3bb9f284606b73559da94ea24a8c0fa64d64a4707a9e3a7e7bce177ae099834f82f1392bd24147871c1e0e8bf51eec8756f06aa2986ffcba8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h874943d7e9e6dfb167dc90cd4f24117227617a270a8e88b44153ce57cd31647c748da216c3dfc106918187103782f33b84409e55b18368e5ebfa7429fd6cf4caf4a9135a9031c141;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h732178d59de6b698b62b69b2eac89a927c491bd52c22df5ccee81ae181469e4a4b053661e7f35a59e11d5e914a8ccf5c1cb8acd3365903f27a71f2ccc4b7cd096f1575fa22bd3b80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91f34c28f4e795ebc8fafacde9ac778e1dbeb3fca42180f86431bcd872fe0af54f87b4dd10538bd77aa01ca25dbaf48ff29b401e1b3a98776446e838f41a2024aa59fcbc19593531;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8952a5560dcfd2c28a2e2c0056f86fa4920db27db2db47d67a091d64b04b279036022a592a27f67357f192bd73ca7bc3ce12cc66b31004a95b2bd0fe03bf9c283cc61f535faa71f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4629fdb7b16bad6f734dfaf1f531a17e24891f2f987b8e69b84b9f58201a01148032088dacedd24f07a4f63464111f2e3fef148b1d7010a654c6958e6665611930ec22dd45cf4bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h732b0ee2afabef23f2ba1ac67915c08b1527948e7c2c4ea54e0663a1d50b15abfc3c2811bdbad0415b93042cd5d800f7b516e8c57492c949b33da3064dc80ada59b1ef405ff8007a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0124d3475da7359f1ce919210ee6b7a119d9b1594c7e4ac8eeb2dfb9ccfde400fc23fcfbdeb6c2aa0d2ac882ae46a4dbdd15cf6eb340742ab94df7e3e8f99b309b57f4208dc416a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12cd4bb371373b02bfa1230c2dfb72721f36f10b13fa97fcdf9255abbca7ce9616dbd04a719a3e81118ec12245b504c9ee79659d52aac7091a9f57e1c1b56d8c5c1538240b29c101;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he43cd1c6bb3079da3b970e71a676dc09ced17944c0b21f1c152cd07290f9f5ac94f648cc9834ebb0200fcd87a4097d265772c25b8d35f8ea6f8390da19cf518d6f1efd646c1d276;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb27afe99c76aea84b23b1bc104465d1ff9a47b7a1e80908e0f8044cfce442655be70c19fcafa98f919ae89f587dbbd2a5d22352180d26f6cd4edd9ac74d57de714e8cdc913b4f564;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc25572b5da73c48990b8c042c71fac9a10857eca678fc5a9c09b8208f9bf4985c38dfafb76dc2a1164e5aed953381bf54615d0bd02209c63508b18226cd71bd7064d46e8100a103;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7cb3837a5d0cc0545805205cf229cb8859837053083007693a01c8e456b4118d859f325e97eebf0d76115505530bfd36645163d21853b49036b9792934ee0949af7af916392b312;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a3409553ca38d6b8d700aca0394761bd7033d5aaa7a0c0bb9ff95eb832abaaef5622ab52f222398cf1cc39ed38c970133fc7f74ebe734b7fe4917a51fa87053471c44d4028573d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce956237859973b5553e3362ed824a16f10e3009dacf041f3b8aef904797fea900a109528f3e757cdfb32ca68a353d96e0c4d0e35d91301e9409ba0fe463e35f519c2ead9cbf8c9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4c11f54d3bc1873f0ec3e7cbc66428f363628ffbf2174f5dbcb28f92d5955d562168bf7118ccbbe8bbe0011507341335cb325c31860b883f3e7dc05e6d906aee8d7a8bd2c7aaf77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aebfaba95edfd475e8faf6ddf60c171cef53faf5eab7d30a3c2d9ca958a9827b9fbbc92401c41fdbe6aade98836ccbd43fd3faa17d397df351db5bb89bc1f014a6d3cbd80511ff5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he79d7cc35652e48e22bb28aafd594bef36fe3ffd396b3b13f8ee25a7e761a636dc345106133fdfa4a1c906a9aeb99452cf69193b9fcd935cdffce1b56dba09048a51fefb01e13ff8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bbdabe4b6f20e1ed2de7d19ea62e7f250ac2ade186dab10e07d6ec873622658db5abd2a6616d98b3dede9d48ce92ec41e6e144193fa8c8ccd6d6335e00657674cafc398e21a5754;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h452e4ed5e1231dc0271f87038f07bd1c32bc29a1f05b2985bb579980757c025696015bf0902ad19f153f072dbb09d8fcf22cb06ba8aab45484739cc7a03d90feb62f9619ba41086e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d71f5cd1948f01a0280850d9dc15f4ccbbc64806641a949d2be503cb3fb88f120ad6451c8a1025e91758374933dc6d35b1f778a4b09289f4c62bec519b4d89cae45596e459310a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8e1834580430ea7f973d615e12d395013a60654b154a76df8f4f05fec3ef0f486ff006ebde2cbc85b884b1bd97855aef46378faf2741de3df52aa02df3c0bc2b024c6c9c92e4816;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heaf23be5209d88a232e7527c167c222d38ae8b3d6c3c07f68f2dfcce29a637d7cb3d33b22eca385a67ead0e4020c169e8fcb3c391633126c04a0949cb33e9fe7f57423385c82da0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8181a5eb4d1e8ee9f60837508f1237c57577149753019bb85f77b57bfaa398f2377481a0aa289ff7ca74345fddb73c1a6c06e727708c28d988d13cd4160aceabc29ab006c9459b69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61e65d975f685406b3fdc3981a8f2981a2aa4d649d160ac52170cfd9b3b43b5f44b04217ad4e86251aba8a5d0cfd2f884e32767c7a211f653b333361e2425956d50b6eb178a7bc08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74498619c3fb21fe2aade8294925ba5d44986ac4f34ca56990bd707080fe74c7deb6ed73b4b69db9c735c6df75ca5b61bf06d18dbf48d993aa12fbfc399684301ef482d44c3f3f4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a66b2d62048ddff2e18b25884047f4d30de8192f58eb217cdaa4b9e884002dffae66085cad1671fd9f7fd6f2f5905b3f2496ee85f3804767ded42bf6fd6612a2f14dba300029a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be38096077bcde734dd37658326612d96a7fcbfc98e51ac99e2ee1830c4c259a6e8d33c47a3d56a76335f598a554b5098535a967af4e8d1b719161e8627a5e4ac5767b889c9c6d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc421b2e91c7f95a6b70b3af09aa3f747649ab7103ae7995325cb2fc656b90ccc86eeaf2a6250dfb193ddb991a19f2ca050a67691ea0c4924f2cf51730368b2be23d6beba8c74fed1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he76e0a6246621058c7a99db1a8449e0fcd17fb485a1c9ad24919ed25825de3ad96f344ba9be7a77fdd2e4234fbca0c15256c27239adcf051b06661a4225b2e887d328da2e6b829d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd790007f025158d7a2df1e99cb8d03ff7da6b6495d27a4c73a8bfc455ee955adc0a1983c03bb55342ef3544505022bf57b92e6a79795c432b256d559263f40b8d173f5860b97af90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9025c4f76e96c0437237e2f04a35be915dfe5979d0ee58734b15531b89afda1c7f44bd500b16cf32f08ec79fe0a22da4a5ea160ea2bc66906e54b7c8b1a86b106741ffd6f27b66df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc209a7b7e14a0601716613f69b4051681d2614f12386b819a52e04b0805ffde26d64164442050095491bab2981f24cc57cf0a752e6582d8f96723588a143c3233f04b4cbb560d6f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50076f528910456e00f6a670d6eeb8fbbb9f7603de1f5338911fa897ddf69a26bd1622c1413e5a9f2892e29f9ad4178f1cdc63865e304c978178de5e9355f4401a9c176a63db9b66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42a33b0a48a88b26b5cbeff548f149b51745032ff33cbc52c29c36b5bfa4ea526009aee178dbded9c0f57edfe7502719d498598a9a902927a9fc19134d8c1304515b1cdb3580c56d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea3bb52786a7ab59da3799b2ae062a95a8e82061b8969f793c0f1b48d0dafd6004bb15679b2024c24a33f8e851b2891a826fffcb86966e5a62ece18322fa6b3543904b976729c39d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2712b2642fed9af334be07ea8339a7aeefdbafb0ae24fca1d387a597e6cc05c85b0c67418e0ab9ab70c88220cccbad48435aa49a81df2fc0b258362b1b94baa29f4cdf309937d4e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h940f71089e19f5d3965213a946e5d1efd8eeb88b2a25a75c91cf9f1d65d18591815f3a1c65d70d0da6ae0f364b1f586ff86d2d569ae51b6c54d2baf9c3d9d4ec80d2dfe8589f0543;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h985161acd31f9167159848fc7ff2197eed0475f7932b9c13f2343c447efbd5a40ec239067da52428fd70efb83a120098e558e167603f6f82a7eb0b119d4612ce8d4ac2b28a88e44e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e7a302c73e90dac686525f4c718cd7586e3214641d44265b03ef7a89d862b2b338f5f761638c5ade6e50e9d50cce8c108d38ced30d86ba1f294bcd6a5e5818e34a696ff136ad5e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafe4e1686b9824b873d7a0593281bb2d1d71986d6fdeceaf6def9c2e0a12787b33f6bf5c01d6f6347862e5ba9338eb09ea08e2b1cad60acbbab22af2e91ef6d2d5a480cd282f43cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3675edd86001eb5c78c752959bc632149c817dab8684750aa96dcbe4941210c1f26352c3a61c2b7ce475c05af153192e9af14187659b6a03e8241aef472c3e2ec216f2a531b067d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h652dda85e9859382de0812eb23d5702111460de7b06d40aae29ea7a5cd9ccfb104af26e9ecd1407c14a44561e5b3fb64be55ca98bc663d5bd02fe27ec40525621c0aa7527a8a894d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h282c8a4250a2b73eb59d182d28de5d4b1dac2811c85db6f29bdae0ecf0251684fb663af19d7dc907edd7d688c281cdb4f2452d1d1a556cd34a2a67cb8138134839bb3fdb89bab4a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32f5f62b509e461ea4daf1faaa0f5b4c84cdc9909367febd4883d6ebfbfd9d7cec981bbf592a1ff36d978aaea2e62423c27cdea688d4a988abf793f038e39fc1e68eedc6e462688;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29c76ece35684262677f66dafdfc9835db0853c1f2cf2c18ba9dbbae14b66fbd9eb3a434822cc06b8a605ce19c6c1147d7358a379fdaa3fd835dd0733db21cbcbb854e036ed9f073;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8da10fb2723b73a154813ec5617c3307f2fc6bf308b2eef9ea6fc3d8fbb652c5c554d5a5d0cb42ad5522680ce3c01da91d6c61d8e742c5e6cdbbba47fbc7e33ef631f5523e47dc23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6318364d8cd0d9fb7e4e6910179fad4dbde1ea5e283979160e74b69ab6c73f8730fbf6a46576455dd821dda9c58671442c3d01fe444fca6bf6ed00854059c7b490522964c499287;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b143095e1ebcaef076ad2f743b128b6272debcf7fe6efd55ca729154b864b25bb0e671ba893efa6ebc4714c9fcbb729b2c9706c364720604ad45113ec365a37ce7ed57fa186545d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79192f0dad10950c5a65e9b0c506af232b746725d6482449d6dc9e83ba34ded1e56d2c8470c308f1cb19fecf9a7788f2a320b6d63a6cce9a2799b20e03f5f07c1308b8862a385473;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c2f72441b5bacc8a2d7aad671ca7dfd18730d5bccaac43c6b35386b9012ecda8f246f8ab96fb8ac3337e8f1e81cc9f51e81732fde525f93ba1899b38c68cf732e165a517c329110;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h530dd608b38ca37eb7f39c822e217c632af539643353114f160263ef225e03c529c7935c72f8cfd8f45bcb5cee4c70a8b665a7e43a3fd4dd5fdf55ba4a6c74183a5a8a14ae675067;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d4ff95ae110309ee26de44c8ba59f063675a7b06344ef647efeae90cd9018fa73fa888cd6f5749bbd77c68cd651f67460c526942d6e36291ed2274af3a1578fa75f0587fb069d3c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc628faf5a2e8725b5e6ee01533f36595028b4750b57e6967d5a3cff99e86baaa3629486e9492f7a3f1bcf752afc67e8cc02f39114980175d073048ec5b96afb09258dacec967e71d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd50feb2d47cb1a503ba929b3c875953d1920a67b3cd2e97d81ef74fb9ad2c2f406c66d496ae3f0b826b325a0cdc30398ff6b8a3887115e6d5a84b63da350cec0c47179e834bbaac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha230fffbb8b3f32ddf0afd09b4d5e9ec328748fda734b2d9db7f95f859243a1d4f0179d5871f665403189334802885238b298e16c98661d01ed3e569f081dff399fcc8573f5cf627;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h376605871bc61994582381a073649533d3258cfe447d4d5fd9f969a8ad036eee10bb05a7c843b65893c2e7b2cbd02533d84598b8aaad4d36d886bd01bacebbb98371d34ea6f457b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5513a05be4133596656b31ea6756d8d4c66cf12dcb53909b36553c96aebb3d51031496a4ac93471752a6a4d504e12b05282b2560012ea3761d823dc91865b157b946961a3dd18066;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcea81c7faa9ae15f69023d72c0caebdc0f32d58e096702ae3f05b51fec887d7aa82c9442087d68c51380391b7ef5034682bb1f257c3d3a64df4144cda3dcc5287ca95030240dfe26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1bb019e992822360960dc450e1494faae1c9da3055c5171d8327a307fe5d91cd7f4a0892bcfa8e727a99c74faecb798b8efb1efa85d157ff0befab81eed1d26d21ea7f74a804044;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4abab0726a62491199d244e8fc45eda1106c65ef703b4c591db2565d991a26964a23a0a8dcb15342f591c83358bec492d1844e1500a14fd84af2eab3783b9210eb9230f1948d6fa8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had5d89bb23529fe7c3fd40194cd190c26469c2a31bbc167f64604f741b3800eda986cac3a81bec22e245a940098380269d50bbb8c2f54bee75280157d86674ffef676c3ba8897d9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d22c28c644c7de3ccf4baf60859efab51dfbfa03ec6a49b2ef0a278405cf77803e8910d860ce23e2f7a1860d25395a0c2b36a1456aaa7f9b88f5b2bfb26df0700a914192153d2da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a0c91e292397a5d42836100ec110d9d7cfa56baedca5d1efc4d2d18173d3e5f23b81b57f079aa835467511d3b69f931c1874b23a6778ee491344426e9d60b3b82a5d890f3d1c203;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe6d9a73ec398be11da7e7b7aac6d8c4bfc3bd3a4f298f8f16d4f3962a9ee56f793e85f32067f271200e276e816e0525b083f3872d2f6a83eacaaeb1fb4d1f61cbeb572cd4536e79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e5b2440017547140cbcf0d90fb7b9508db139347dc9d35ec8fd32e18d1be99f96484df59a0ab2414fad79ee621d3d27d14e733538cd20787856238073843ddf8f2185876db97183;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1acdac992692a27c142e0dc96b9e5c2ba17ce0f72a615fe926a911c369e8fa7347cd990653dd9b30b047a7247b70a72c682acbba94ea0c3b94ce5f59810d252b3e4fe7b2c521db9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcaef356c2a4e904a61adf90d9a1510b7efdfe94a7e9a4ebf9f528c2857b416a2638c312c3e035e735d37427469269f514738408367305fe2a88cc57bdfda5609007a1a12c9eb7a56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2b656ef3ccbca43ec414707457ad475750cdddab7f398e646e35ca5fcc7345ddc05ea4e6212c92c946da1153021a84b63a4a40289db8c82a11d1a41c5032969e9523c2c53367762;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba8c5383ca05e681d45fdc608fae52166f15f9da76d540fdf94cfa7a437d786a2edbac8f83eeb2f4929942d7e73e685377cbedb549f319b53cf07bae01b843209b28c0adff77581;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7042e68db5ae533d19676d1071579e73b3bdc6e5758dba9918d78037d730da527ba8fb12db82560939b7d8448cbf220788cc09f6b81b9922a2d641a397a4e614c00304f670a1c369;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70807c944f9f6b25504a86ea0768435ced5e909925d37df14a3e7f908d62943fea00cf9828302f1048bdb6489c72dd3be8cde07dc8a3501e71488b797ceeafe08d981a772c654a2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h917470d11d52b812e58b924a0080099237d6587f977bc47e7fe0fb5468c2fa5a66a3cbdd92a60f377c9e0089ed2c4cad467b3f8e2ec54539d3d785baabc6a42144022c589d7668fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h931ce46a7a1453ad478dfe209341354ee3fe64cbce2043fc790e224b8d59886a63c75665d3d4fddd9e718e2e1387c767df0314e108b7c9b98cc62021c874b052559a6ee594cfd6a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5484c04c0b550de473785134a0db553ffabf2b445245f64bcf5fafc44759118a03c172e1dbf465578fb9b9513b0777ad5a0c3d2b2c62bcf5404f3826ff4f1c1b1d24dbfe0b436a64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b75349f54e176bf756ae51a001439db07992e764de27e84b471d40cffe9df4f796c4e45bf25ee679376940abeca822d03af3d341cdaed333ae6aef7604f5f2932fe5d39ecde713a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7af7df260fe7a4c2ceed95bf56d886b3da847136d7a86aefd8403d691b81a65a2d8d523b5e4cdd46dec30559c993ad554f0f8179d3fa39b1d3b8060662a23832372e38a67551ac4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h212eb8d1403bee0d1c74af53fc414f8259bb03ab36f10b4369c8e291bcee68074e5187abcc699e10955fad5196e7c4bc19936828670366a139222e18d6c2ce1bd48cfc92a4d222fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e3cca586de6149fc34370378e98baea403837eaecf9f43dbdbdd7459de985e114de126d560349a6a21c1c312c18facb63a155a9a10fd8996b53d9d46db7f853499d25e6ab4e408;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h190c0f4bf4435872c878af01da0422f13c2366a8061f4edb34a67af1b71dc1cb876640d9de1182638bfb69e7f5795f92fc82d2019b08b3856c7dae0edf6b9dac74dcce749e21da98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h770ad55a9db68bcefb303127ccfeded3392789e45e435caec6abc992dd91175078391b25cc50b7da649194565f705aeb47de9bceb8f5698f3093d45b7e8464f2bdc3f303c16fec11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe710f5f419c0261f36832546c63dab18f3a975ed7acfe05def9b774160d9212c144734d49a46ca40d2d37ab71a2b947009d0e5429098ffee3ea87ce7915633c03dfba7407d860b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd623354456d284c4d385ce6d1bb6876779007b2e363699fece24bdbefa8b308cefc0d72f175ab398f24743abea472c1d396b49d1dacafea9ea2fa386211915371d4b88b206854660;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f0b6bcf2930a1f4c5e8262dce0375c8114c4dca1a2def04d78fd4ec9ff1a9081560fa58d907b4d54f82f6e1000f5d4aa67b019e02761098457ae7ff176a1d4d9804c7d761cf2b08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0c3fb9c07334d52a25e42caa392aecb75505ef5a51ab279ca4db8d71fa392333d560fe6fa1a5b9324a8f4638308653a32c643e9633f12a21bd1d518ab79d307ef81c315485b7a79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bca80de1ef3e232687eff933c6ca521d87f28f144253ddb2ec48ec1405025de618e5a100836618fee9baccf8598bddf4eef296aed27787dc50c6e40398aae6a021ad59d25f1a98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37cf1755b9a86d6ac99b0dce098dfd447b8f1329dc8e9becdd897586eb6531f94780d2bbdff5cf9cbaaa1d627333cc02eb3483f9879bffd0918650696f1dc81fc1ccaf775dbdb17c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda3615070cb05f2f61a338a2174a7a58be9ae155b8f029c6a7c3b324091b1adeddfd0edced035b5a416762fe878278b111eaa5bd90cd13032d22e294c72aa018195db5ba2ec14693;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97ee6adf38d4f60c68b5ca6fb15faae267abc502c9da5db5b4b4f8f1cf8ad9428fe18d08b2662bc5cb112fcf387b9adc6c83004f32378a3151fcaf498caef57bb394968394a637e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd45935239843c7b3f61ecfda8b89ef03b6f20e2c57245e42839af37bc4c976e7f9e6f70f6379521db08a601604752629a5049504b6e1b8515d9ccf3c0217c303140d84ccfcd11a6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb651cddbf1c3a43c68921bbcb24ff7c9cd65b8cbf585a8b03d3227d41961acdb0f41cd047e68b6f9296b870145cc95ca553a5db4897c585489087073afbd1ad3f6f27de3c6b7c30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a7e7d91d3d89dcdccf06dd60f61848b32811b42d336481409ce674aec43a76cee18728db95909023e72f02c5e82c8a617b4e5dca987e60ab8d330dcf64c6e19ee9adcaff4e32be7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79a1000889f550fb19a1a83cf839dbde4bf69a4668997176cebd7d8f7ad18cf123b43761ac19351bb6c82a2b690e67f6b79c3f7e0296380b5718d86cd89737d73601285294600fea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0bdfd56985f3b0194e5989c3704982bbc8f30a88980eedb178aef6dacfa566eed2f36b1b078022a91e60f39d0fa74f41643f05c65b01c91cbfa65802d147fef29e3f013b2382cdc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h601fd72f204d2bf269ec8ee5411a4b9c1bde108055a99f3d4d450b9f31eed6e88bb5fefac02dda7f672a1aa3379bb70aa50b2622ce4153edf7db5f87383bbc25cde5715c8c1de186;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h274388d1c7e56e4534e12bfa45ddc28380822e611ee12870ea9fa3407bbf23e19e747fa43feb1059a59db9407bd87c4eefa0113ba7be2558dcd7d51fa1afbb36c00fc9364c4e4866;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f98ce3d27d71bc38af4d301e916ba5a97f2888b13e0daad65b5964e4b70a5c238035d75ba738b98d17f8cb5c1268f99b9073e637aa456d3e9de137d31dc1d0d2e2589d239a321ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9de0f60b783d73e0b05ac0f607405733d2deb04f3646724f6aa7f3756d17d7bf5401a8c778e83f538f1d2d6885a92271be3599fd51180066f3a0ac8f47f2db5d110c96897402988e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9eccc787eeb5f1b95a6ac55741a7905a99b8f5490dee4c87f0e3a61e8a2710e28b667a8d3e69a39ebb51458e47660d4c3efc0e0933806b2d90ab2e969d8e1cc018f0620ed1cbffba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habd92c38a9492bfe6b6e56c32e0a18c5e081a40aa2c0fef6829240c9d40531a51ba1c6d913d9870a75aca55412667847f2437175c086cf41a15bb232886ae0bb761c58c45ee31a0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha42fa81c769b4c8503deba364a60a310f4212b04ab5e78fe31bccd5e4ec688ae72439fec43b0272370ce2445e6141e88d5a67c08fa39c4adcc636c7c54049d726d03c55539dee365;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedf9c7a4fda32e8a456449e77d2ae74f37c2bd734f6ef601d05884129c79460df86b9f14fadbae763022d8b31d213eb42d84600f839a88fc2fcc981261db34a5b1074026619f923f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbee786d1fa08fccad6a2274cc91d7d98a95d320f936f2ba4d9f3ae65b100fb4cd45722a3b18cf5da209c0bd12cf71c9e31d4733ec403a0bacd6dfe2a1190de2d0f6e194c2808529;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb99fe18441dccb6d3e39ca7f524dd06e83cc8e003cc8aca69f8100c677f7a0f071363cee50dfbf918010a4a1926a0aac135e7471760072592c5554b89e7eaf6d3592a1d5af186a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2a791f5f50f5f8ffc210379cd4f5effc3feb0a169a787580fe8518b3318c39c33cfc72a3e7bc894329238d97e8790668a9fb8b9f1a403e679ffe1c7363b03b2ec5daca3e0f8186f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8932452154d3621671a457ce1c872e7409d92e15d1ee0b2e64475cf92cd5bcd20b65f195dcaad23837209cd124ef1bf3cf944b7c6c5a87e1034c0a9b8453f9328a94a113252bebe4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haba5924fd9392660284105065d4b7cad98518552bfa4ea2575a71b32c52a0e37a3cad1d9637ca25ea2b9fd41f053475ae9ea0713fe9d29ab6cfee94d76b404572826de6508dcb153;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a6bf316547904fe27293f28548094747fd93a7ca0018087f19117484aa62d4b1b1bafc5caeafe28b16e5fd9c3bf25cd84d0d246cc1dc7e4116a701af7b0e124c66e7e6fd657bd19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2938dd6761eaf4cd647d111358419865a197fb63a6cd4fcba43b5b72d7720cc59582b4848bfb2c8b73658c8066f197123c80ed803c52d6ec08a54bd22128628ed03e6c9ab6e58b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb85d0fc877dcdb92cfb0e757ea51a0c11733f4322868c62f42601e910e051dd354f9912ac7f8502b2a125af092cb7dc3a742499296c74d5088d5bb6b7f60aa48c501c561e732b38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd54e152bd773ee862b1d69b8855051c747cb05730753693df4f6cb690d2ea89ca2231b4b344d27e4491717197eaa76d1fa688eee0265de7543951b55b43f2e2ddb9992c9b03acd7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b969368a9525b240369f271bd8b77be18985517915cf7124b2c96085139ad05e92c7369952027049cd17c91e9ac6351ba70a00cd2730944e67d31369c0e34707febc45b0f6385ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e5a8bcab298c1aec49029aa1c1678a53f968670279332100be69e4dffa4eefb210e88c49ab8e74fe9b19f04d9abad3d564cd24e3783b2684772b9b1e5842e75da723a5a713b412a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92da444e110e7a78028464f1112eee5c161936656cb68bf24391c0b3ff3d3d948dab503939c30e93a4c6edac46c33b6040ab3209e2831a7fba3f35c19bde064146ad9f2e2d8f9296;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea36ee4108bc9d743936f8482ca9ce2d91632bfac884aeac22fe7e6b85ce850386b57ab976299c590bd51a8585ba7900a7b0fb4cc0f5bdc75f23a9fb62f6175f31d547917804c716;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf3555f7346bf09264267b2ef384c7fa0b49fda0d1aea604a78d5ae22a008968c90640f175cbe7617fa3b0d9ecf03bf292abee207ab7400ca31cf73f44a8e170fb8701321ef3dfc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h171ff186367ea4d43f22b89ac2b01e6579618283670f7facb1282173551fcda1ea5bf2d8d4550532b40923dfb66950fd5a587f3d9e2d39e761068bf74a0c369e94bc39267a14f703;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h335b0146b71cd29ae90aa8b4cba20c881b34e211e07d93a70ac8df7a60c4275895669e808778fc7f5b3117e698df675b4c25e5a4bc732932a9e0d178ed1b137c0e7fe1d303d9ea3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he76f56fcf504b90c5d5a3d0012f6915f0a9cf0788b75c64c0cc93dbeb0c5c90d14a8c7ec7dc4ec26095dabb98c245ed3ccc4572e08c7179217c21dc33df9fb7c1acab86324f45c2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa5b042c588fae1a19b75fbb1349c26e3b3b5914193923d1f840c7605933b750680887e77082755748b6b048edc03cb64b1c51e1d976ba53a899c9b25b9f89a1298c28c9af9e57e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h336cd0b2a9036bf221d492d11977e780ec8feac2f95db873db784ef53d6a384b5fe1b262e62650390ccf5fc14f72c152c3fb55be0eb242378af6843f893d195a566ef6f4f4d9e121;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67b92cb604baae2f9f8ab8cf6b849b1c181558c4956fda0933ffe6caa6934ada95527361f16967845a759e91de74489ce7c5d5deed947e4561aaccd1993c5a6db875d18fd0839d75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d6868a54377c6ce57fa476009489e81a569eb8313d2f260fca5506009c3cbbb4d35c42a7b729ba194b34658548884e352aba38443a84bcf7c2901a94beb6d836377df8dd68876c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35b69406669712f0ef6a7bbddfa7ebd29711f23bb32121110ce7ca2c5ed73a2abbdd6d52b6750d354eb850209c803964d23e70fd9bb838f2433376ede74625062df4971e377396c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d58563f258639c5b08b2d1becc18e526ff4b617dcbdc32044427073f2f212b0add812bbbcb8fd79b8cbf228c7cf5ac7184b0be0c8dcb20df6a96ba7d84f5cd186332ff5261275f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a208bd1eb00f077a20842958b8c6908c679eb1ce1f280fe34b236d9b3564faab0ef3effb45828438e904145978899cb4eb88fadf8b80b284242bbe1e438f2c73bf5d9f96678d8f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bf88b03240ed1136116828760496f34a1963c163799ebcd79421f13ec225b169be417748d8fa6644a5c294100500e141393ba7ac88d6123222d6017578e4323ff2e168c1a941baa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b11f2e6e6ad2af81a79d189c8babeb33594f2980d0be3724401ddb694ffc78a46d1b82e4c9d6db89590e838e3c15d1840b0c1d5fe2236ce3480a9cacf190e68359ace37d20f1d89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha777f69943479c495d7f6c6d57b343f05381844fb428fc0e018cd0dfecdd04b5f4a735d327a38320f840b3cfd9e635a91e068e603e3df5597dc9f610a261421a19f1159dc1db7389;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba8d682e7571bc1efbd15748c2f2b79c17a637455a13cb1eaa87bc97a50c6c7f6540878928c8b17babe4e206052633e79827cc56f8b0d11fcaad1e7882b7224ba79642514153f799;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6774393a07ae95adac63fa430d0139e9bdb75687c7bb57bef0b007fbdb487000400d2fbe8949473120e5b8e5b4d4a65d3ec377b0cb133cd42d417fb3c82e60f2bf4f4eae73a9c01c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3bb463dc55465459f191cb584801168980ec1e3c50b50dc0d902b9b3bd5eeb59955ccc2a94b63d3ee2340b43a2ad8fbf884ae8782b6d42789676eb68f15f0a023fd263e93290259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d6c61df5aed8ecc788270a4bcc67315553774d0bf28b58b66e7690f5f401515d9d59bd051187029a05a697387a71e8b72db16ca2aa8a5dbf4e50ffaa7a8ec77886aba8e6e9e5798;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1a116dac61a1ba09e557f90d446cd0700a39a24f975d0c28ab62a2fc618fa6e4f6ebfb8412cd27c79ff3b40be1a6cf930fd27638a8312e70dd2d2d3aba67b48be8d05493cc86fe6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha299bf3374602cdaf36c650120097384ca848881f50802b2855e18a1c9ee38751e1e2d48e7dad8927329b901839c0def2727d2c6f51ce5d64d2b065515e73f3729a533eeebd77b4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a3b3f85799f70804c5026b8adf1f498b26080681b9b2f9039c3768dbde1ced1bfda809c661a29dac8b7c26515d60ce4797482f78c3092d2c069439fd6fabf08b7d860e427d5e4fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26aecbf987232dfaacc7f31913fcaea6272207279f92bd5bdc8b5c3c5aa1e622f56e29f296fdcf1dc883d14e5a375d2de0a0eca6ea287c5031107c3790189f2191b007b01612cba2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa4310475598a9c32696feb5813c5c5750ddc5dbb0e704687dca822d25b28f597b365a6498fffc15c63adcaf761412ed34f0705c9004553211cca7ff2267180f7a33c46529bcd627;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h672b1b5420218897381226ce8524551a32ffd126e4dabcb0ba668d4d1e702052f177c5a41175a776d1f91860c5a0660b71606e9c487591c3703359f0399dc43e7ee4f51440ff117f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd36030f1a5f5780466c0dfe85e4de61150b356049580d790375957ca2fe12039b7f15a610d05aef22bc5c0485d89563666fb2deeb478daf1c049d031a0a286f6e11601111e3711a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22308bb453de6a8daf267d126434a09f482672818f077cf9043524cec19f8cd1817e8047084d018feecff4b5cf3f73f0c243e8769dab36f2fe98e4d8f3a04da477bb05667e718f7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47e9e4b4aa97da9d728245c16553d8e084c8806d0f069e5d26565fd35f53fd0d1c0a206a807e10cc702190bbcb2783218046c706c7d94fa5fa2e2b1d567dcce82469908140b8f7d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f847d86d4497ea8ea6d17a1bd50c0de3d286b562f37b129e0a7f8a9757f71bc88fc6547dac11d55530fd1f5ad176a2c832ef8510e3bce663268356e71d813f66de5d7fc75666b15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h356594f019e8c71529450c395ca73e1f530ad3192e7cae1310bede002d6ca70f4e633f1e79f1dc7e84c90f3741b4709db0b25f197cc26f905aa017866c054c13761c4a0caf9e9466;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heef74a1099d8bc55d3fda5f72b4825a0ea785ff602103baf30d2cf61a4004c9e7ea6676a323f0bbf3fed91059b0ffe2c2c814cc826a71b3e4dc4ef87dbd0f03ee353f5986b2b5403;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9d5979810357663bf67486884674c9f3897bc94d3efae4dc774686e0568147014e39771eacb8edbc1ef5bf5adeb479771b29ddb12642f24efdc35d7430d070317b6584f5bb1d99f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e383fb45b94ed1287a2bb1129829a157d58acd308c5bbceb9ae2ed8df171089774f88e143939e5346decdfe0bcc1fd22d0491996ef1ce9318a066a57ffcdd2823cfc8bc2841abc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a9a41fbf355352612fdf51f6230c17b022a25b82b72ac16c71fc99a27de6853047f2868f5573b33da5f707ef5f766d236ec54ffa405d17d17e2ef1d57faad64406f385c70e9d35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78b900dca77d289a65189a8bae2277dc189136825cb5585b4204ca15ff84205bf221027eec0dd550ac9d2b9218996ff3a3b8eb437c32ffb287cd55c249fb75922cc80196c3c828e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h456c44a3446e47ab6c01829dfb903709f90ae12e562bbadc69755491a9739693fdfd632df742147bbdf4b608b0a5863211d3838b98831de11848fa7cc41b609e43c64c61847a8f7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a7dec02df3aab56cea46ce912a0702f9e7d0ad54a24c2694c6d9773bfad933d22e1bc2613261b60fc0bd28e5ecd937ee501194cbc39f22a9cc0bce143256d1943a328a9e490ab00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h540b4f8b0fdff857d9b7b48f61bcda24bfee88474b42bd6a16332d24edd93d1a3e9b23abc5d17e0ae53e4f7ff3fd167d27cfb8edd971b992361eff02cafbb05d887df94ab013c6ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h927ed325e11ace2e45e45640466bd9ee0a87d196acdb35a449015abde5beb98142b1ca036a337e3d3c69a914a49ada053008dbd8d8097cc4d44ccfa0a181941e98a7537faa811fca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d75b92d6f5675b716af6a794a758583aa61fedeffaf290e8e2077a8ebbed8d888533e7d581761b4bb29d2bee279c7a44576d550ab82577137a56b98fe58918379cdaf4ea1d22abd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95a1d01436730a4f843c1bebaadc7712f1211958604dc4c3df49943de19c789b3911950c7ebb66457823e47b4da2864f420d004348ea70d7029842c093d97aeb60a7db33666c0ea2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54277fff06321fc3a1135c8059c63539d7534d814c7696ca1fad007a03c6ad71e364170143192221813de67bd8ccabf18f46371ba534dcef11eba3412aa8cded66ca7a8f3d79cbcf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bcd5d56b66df2e7cf9b3f4c39f49b389c075b98eb4fa9c78519a6a66313e7e180b615058cf0922181d08113602dd2aad47ca90dea95fcf457740ab877038783e7c3aff843ba7230;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f72e3c36e03e23c4d89402ac86df88cac5f20f258a632057913b87d1b169fd511ac1a852c45f155c7678376700b2e45174de2ff539a6f88f48275c20bc70c0eeb9f7553847a6f84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he79e1277a6c513ee0e028643581e93b0e1e8398dea5f24ed7c0eff77d6e806e0114a0ee181610c303f748f1724e79a0ccec952284aca7b7a512ccae8363babab3c7209a1e6f114c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3659d86ea9036bc125e5060c64f286bf8b63aef03e4e32f52bf4bddb9aebed9672f1d6e265aa3041475805e6e10597738d088f72d7bbf89b47d4679b6e78c6344fa57ea8bfe3b337;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h308df34149e1fb176ab1f745317820d0a942e6154395d9661505567bb3a1889cac9228f840d31cba5aa7800823a65767c325d77682daeaa6292ce93f91667f8090f2e9c683e6d118;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34a35ff35d483951a5c42bee0ddf08f2c5ca1d4981454651a0adfc5b1d664c9382e815918af0dcec8c048e84ba3e55a133a0f2bf3495770be26cb3f70d1007278d55d7935b09338e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h704f5655bb24cd2cd4193464a3aa486c85d80d0ca7c4543bf7c31030dfed6ebef04593a7da63d3b400a761484be465944b621f112b60650112d844d9543057815ab5e391c6eed46c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h259d1e9271f0a2c80728303274758ed3ccc00b749fce96c175957ddf8663c43b4ddb19026e922f0a61ff77cedeb35d9fcd660c59031224467c81080a623ac07ddb7aa621bbc070a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dad1d93b6a023fd2e1c23223ff58f32f432c69607f348110e92d89ea0a7f88063b60525ab12236354f1c7bd91b0d19def6009a283276c0a2df5d15d4372a271cd1c2b3613ad3d68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7005fbe1df48f2ebb98a8d0eaaa08b4882e0c92f6b142870568529bb6996edeb757ef40bfc37008edac851da3c178e304da3e599bf2d4f981e891b3c29ed88692806767faf8d358;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90237b1e2ea1973195838526ce5e28d766879459555296896284f1e7207dbd85f1deab40d39cd29d3709a5e956b99aae9ed23cdca09d6e74efdf01d57e32ebfc877bb2d279b06c98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee2784191d879a9f54b0229a3d552dfa5c880a5142c0776715f1bfef1df61f44b5e3aa8b296c652d35a66ae0318a8b4f31cd65b1ef2d7c0929cee5153920c24f151e854eff21daf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h502c7a2604f384b1807e156d41507e2d16a5462cbb410b1d5bca9d55c5d440a061449c06e740e687db314937a85551479274c2d19ccd1c2de0c9f71ce98bdf85e857fd1af632472e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a5f28f9bd7d647441cf9d86cb89b3724d902714838a1ac60fe396b892c0239814ff3614196c030e9ae84f6a6183bfe65286367f2e5e05eba8edcf404036f13d249bbcfc1029698a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha158d12d10d93d15c7be5c944e49dcfd8a0a6e0dff0923e40e8e79dad2ed3d765ef97e96530498e05c3edb60a0bb5dc4011cb9b04ec3e4fab1706fd169945ded673a8261e6fa1bcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54215ae90cc9892120f595b939c17716c40c31930c3c43ea5c0570b2d1f98a2d9720e4697dcc21623113ff4a6df2217f62e85310d6f2a337a87eaf118bfef1c16a7509580ad2742e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72f314417c4acf30aaca427a2c009ed0be7ebfdbd35ecc5c2413e0e0ce83835d070c923108065a3ce571cd8aed1bb2eaa42e3592bd2f3969328bced02fc3249c16a823fcb311c94b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d1072cc3e0ac859c63be373dfb4f2e77a420588e263ac3fcfee2f409f9416d4d8bc50a01c9b002e811d0d54df873ef92dc8f307069ac9517903c457db9f76c12769a57a952e6d73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d0207a11b0326e915a95f977954b443b45adc6687666d0fff59f26fd6dd8de4f8320a6d3683e789461b26462a63e37d80b27eb1520e10cdd34b1a1e0cc7f397bd074e5ff072f6c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e733058cb522f658143b08e0b46ed12f6c76d5406478582177618f33f49e3599d36362e22f9211572f7fe1accfbd08a11c8ea31e2a57bbce0554ab321cf38e16416e49666d0922f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb524087b236e08c2f713a26bbf53f7ef0a7f79f7058e54785545a8dce5ae804be148e1e64a29dbd3eecbe25a68572f8ca8c6109535aa6a4e5ddcec9741f6c4152ed17c466a44cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a791d0d399d659e37cf5b1fa7327f1fc5e5063743560d09521f94bb5403cf330f207a41f0cbf4f639a3e5a7262ab57a1b7074cc6bfb9304b98c3fe5d13a032611b04871a353ab50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h924308daa9426a0bb4a25584aad4a71b2b61a42879838476897bf364b6695f59d1d050882c2591a66185e261d18a014b52f794f27413ff9a09925531326b8a1043cb154d7401c41;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d97c8f0ccbda13a8f8e5c17f284146722dc576b65fe859eeef51e7fb719a12890e89b1510fa493ffccbcc5b860a8105368aa9affa9227f9a68e218da7e9ff9f86a6d63b69933a9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bedc5a0479a3d7f50203d6999f5086b52b768013d2a59298f59deb52b3a7f1027bebc9e30a6f918faba9d13056559c15701641f5495ad261c4ff8c5a1dc9f6210feab19dae1b02e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd90220cdc485eb5ba1a8a21d95e0af66e140aa113ae790e1223d3e05a5d698d73665283879db855ed8567e43bc7b6af9cc149fe82dd4355783208e459ae2bef3660e1d6992a4f554;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dae5b4dae4c60024ad84bb112a5c0b0a9a1369a435d223ca86d875eb9f9645e08572a1b018044021aa7a7648744583dd1261d0a5f31482f2f113f4485b49b2062c305c2a8c9d9af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36406cc46e448e8156b4bcfb87e346554fc915c78dda6f4dce2b206ccd7e5705d0b80a26daeb0802e273792252bac34cacfbaf4396f26f2113f8bd546084d294435ac961aa8c4785;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd07f2489277a0c68a1bcd6ec0a4692773548839b4d64c363fab8eb32f0feed90d69142bb5c33ef84870d72b7f69a8f985ceb24f3167c027f70f9bbaa30267475f6e5a15e9320b39f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef9c8823b8a71465a3bc84827e9893c2425305620ab999ac1fa5d637d7125157834d7fcc21a5e462779f31d5a29e73b72415378fa5d6b8b7960b21b73e5224e2becb5db6451d72e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d508ed869985176f835f35570b14ce9ff99028c755bc2581da07826ada068ced35e70bd0bed5da5ec5b0f2b98824dfcccdfa720d6a19619669cd600202c5e99d429d4f032828f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h258881e5426f85e3356a9e3b9156eb1083e581f607886442ae61f691931bd16621cf801531b3c3b1d51db11374382012880ee0b16b282ba2d0c903316761100a52dcae794aa886c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43b6212eea695d179c9374495e4d916232ecc099c7918800a7e40dfde512ceddfd59a77519fe67bafa2ac49f9d44d5b490bda4967126ec04faa4cb00c22b82db5d7afb11c0e0002d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cbe1c648fca65399b096ca4d149c904e5c271ecd2c6362965cb211e81def9d6a9d4a00fc8d01a5b29f80e0e5b6e04a005c598373b093561e241f444c0c3e1038aeb07c41354ec93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2183b520d64c83a11f5cb6b77058463c6c034bb3211851ae2474060f87c5311482db21ee1cd1ea1785edb715985600375953ad5d800ef0d76f19000bf96d326b32f24160c64ddbeb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had37971c0af78cf2f9acbb5922291880752dfc1795b1b33c3e2138c9aeb416a62c14344281387a034ca65757917f17615f180b0f522724f033588df59bafc2a3bc5437a8cb753ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b601593f312a76d2f1c5ce5a3120476886fde272c4c62d97517efbfb7f3a3373e6aa23d8b8a6a27169c2ec358a631dab5e57f519a9392c38399dbd1b72e75c4817e7f5fd74b866;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36a3f3afbd43a7376ae72dbc8bff31f71b8a9853f78bcd3586df0a257881058d0b3eea384bd22470b654814e47cd2a3fca7169b449c492e3b3bbadcd782789d8fd106554b8c6af4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b01f994e38d0643930a17a74dc9bd229cb28d33b1433b60f51d8911d6875508a3c9f87e0c94866d97449e26dd9c03e8a5cc740e54af47b90620ccef319c4f065a5305bc47096561;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e47749974eb4fc6f10bbfce15707749f657219b29f79d8b6a1a2f9e32c19129a335af7e3c19c8e6c2808ebb49021e0894aaf0b98433599402deccfd8612674cf390ddfb56caa4af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2867a147e5fee46bbe52fe14654824b5c6fe9a7716fa9db7080df05bbff709548cb6790b30da23ece5320e0f4d7bc94042874db736a534f8a76a96494f30a8a9beb87cc8a1f5148c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc9ceb135eb20eef0bb73a826bdb967155570711619bacedda18d0d7430d8c0ea7a02b105972b1156aba41597e97ad5fed82b48fcd4db700f8edf743d7b788f78f9efce1a7351ec6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf79deb362bd5674ab5cef0de2b0956e45a0316ff7d6ef0400253f78f7d36ed1d852c03dd0765cf2e73ecbeb324906e5eaf9c293f14ce9c7c5c585f9a88797806d699ef2c32e29b29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b71f1f9b3c87e20694f1c2ae40dce234ab1a22ca4a82714ec6389919eccec24f6ed8a1dc6ae8c7e62ecccdbe85720b85de42ce88862187cb172dd1bdc75205280f8520a040f9638;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ce24143c31a37dba13be56446719f43f127c4b090a74d7607ee4b28a9e96557f3c17ebd3ffad149926d305a855eaff9b146afea95e9818a706ed7c4dfe1985da7475f31ccf1d3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e8fe5001acfb594a7ba1f18bf187a45f0977144b2da1024f62e8cc4a40af59f72ead3b9606e3a1b8e7f4d27a0862b72ad8db00ba6095526c4240700637010dc46fe7a756d8cf49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94384bb37bb2d24b2204009d4ce79187a75c72e8abf2cee2bde48c66cd05a2c0abf7dc14d9955717b31eda5b653d7edafa5502aeaef158dfa36fc57539639334bef228aaf222e734;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7241a7b2b300fbf5bfcea68114e0eed8e14ce8dea425843886ec0a48766ef311226e077f1aaa57aec59106b284deee0e239830308cbefe5b208a6ea1e00638a5b4f39e45a64ba7b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a690e11300ba8f51ea8ecc59f0e963a36de6743636e56948c831d925d0eb220eb2e08b9f4d6fb01645a21d305b475e71cb941186e0d1a5b23f07e9f6bd4bedf4877e97d56d1920;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18c3d30dc33894036f179b0449383babbf2de3743d10d22762382ff3d65da679d06b3cb353673ba781dc7278f036a84ead06235eee72fd2a69b2b1a6d88affc24787498c7b06f2a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h487f0ca617398489c171e0eedcd42f8d0777bab00a0aceed111b325c910ecb12d05ba807f22b0ea593e269a17da134cea3f1d34949b287552632b6866530b3d5a0a32e767aaada50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fc6902b6a9178c575f68083d802410e89be4a8710e2d4160a48fe2fbfb53c9a0e6bea1e4b508df52a5639da49b3d75d4ab02a27393a31d8ade4ae43a2b9c72849dccc51abf55d80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heab77ce85452e185dfe07d8577368781152554307c54c8fa436f1f0cc0e6923ae8e6ec23061011fa2204af06f78d8aec714ee4d065784d564fe392e2cf063837db5673b81266e736;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9ba3ec612c7f5e7955bb459ebc972ea046fa69a42d39401462e841a1301f65ced4a4cac1fd9565706265af2c4490a733253e59bc27f008c96ae4b9ff13953307ef87d6c1e772644;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d1e8800d4e93751e533fe032b770f34c7da12baeda2c4084e9faa75f96bd6bc13766d2704e191637a8d144f9d5485ae86bed587c6c07001a7bc41545dd8b5391e4d0201f7a45651;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3286f0e454c0136200004676f00a456761f82350e2344014c390f52230a5a415a3211b45ab04fb7c8d909262be0812362a17ded87cea88f98c30317feb9202896bbff1bdc8714644;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4c0e24a1e751fbe500652ee7313a8944ecfeeee8ca8cf45ba797f3b4e2673be8dabc2243f4debebe47e97c6d2ed7a3325d8a7a5543f3b90c714429dd5c8c35bb81535dee9d665e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h198a58028a7b59ba23d8e20dbc3ba8515666714d76d99197b16d8423c0e46aa4142eaf8bd7884709bba1475d410b6893f807dbbb0ba111d2472ca83827d9063f6c541a43fd5dcdc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5052582285dcc484d4649a52ee0eecf421b3812e060c3136875aa9596f02948616bc475a5991120dc2fa1a96e0c2e94524aefea708fc5dd2fbe0de00ec61f54f589961c29c498443;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf67dac7d87b41341b9e36c444f5d7c1f0214a1110c1bef8be8d811cf03c114683c1bb67ae7fd51e661bf606005ad79ebf6b3f086c0cfed72676ce229bf795ad5f502d0129d19aee1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4692b7b405b18aec13302a9c4c8b3ed2413ecf24d8d5d0ed6493f28e77481e84d4748bbb340ad23fe5bb378601f58f79979237918eaf7371c25aa7cf83bf9ef0067e007acfd6ef15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cf98be1d7d2b3acf0eaafbcfc02627ddf1b80f6e8f266a2abaf89c83a6ee9d04d42897a4484a0dbb71ce32bad091d11a135f2aeedb628d9d33e90b171ba1d67845cae4cf7f3b700;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8142a887376c01fb4b0f2510e0fe0c391ff98cc947d2e5a2937bb73747efe40ff14ec263272651786bf66fdf47b90342caec69ce9f4397d0e6bddfb294dbebd3149b64a9af3582;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86eb471e07ecb019197d347954a63eb9fd2041c2b02684816ce34d5f77086be753fe20ed8f8b3b85e2bde32417a95505133cc6f296aebb2fa49d8f089c27b0af6d4a38ab58a82d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b3c55dfc048d93bc83f3f219f008eedbca0a030daba2a1c698bf3c56a18d8a10a66839de375b3e5cdbe7a2435ec26183faa3b674b6f769cbae2c34938b75db67761da07a43ab810;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e130f1f8608105556803b5395a9ee8ba0b33267b7239c7786ddf7e6941ff1001f6e71c07010c084ebf2ff64cd450337e5bdb55af3ac7296282185efcf0d2e2c6828c54c780a82a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcfd595f95b9103cde2fbcd5577ebef10b86f2dfda065f106b607fdd1930131959fc95f80b46e2f5b63fe1c3c1549953582f57cd5c340e7bc5149a23f7c5973fcf7b4e08d03d2805;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd62f4cc4913c156c10154dc844501eda46b6a3875b861b0b006888c3c9097dbef2104ed9add11398a403acb5a29e6ecbd2fd3491b8a318f2042b99b9889d70d3a9514cc9376c43f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb5ec4aa7805e9d071e26beeaa8da0b6e8d6693f9b093cf1b57ae2c59e3a136b85cf8f1a513063954aa3e666e769c19db388edcd06a5b5bdddff1905b4c2dac9bcd6f35994c1d6a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52415e95a47a82c0ef5168b2370cf8bf033a2297c4dc428ad263b34f07af4976ba589ee43ddb5222cb35b7fc63054bbfa1759a1e726de31c5c2582908880ab1ebc39b18689d92ede;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22ec34df06e7d9596332beccd606672ca7f71438cd1d2e5e564fed05c5ac7c5291d2c2e3677c98fd6466855ffc65b7a3d755bcb83b4a26796d770d9023008bf24dbc93b38f8d1bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb14bf32c5a55592d9b37cde0d8ac3dedfddc075d39f9759c6c4c720c351e978fee47e51e292bc4661896c8b7813c3264b8fbfb1feb94f76d3d9c6fdd858210516e26a4305e367ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7eaa95b0d06edd9a95bccfad8ea8c0a074d69bf0678a60658b365a2b80d82bee2ac0b24550680315ea8a84fffeee33b33ec81fc1b3ce655ccd5abf28053730f5a9aaa4b1e421ee1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5595338dd523b490c05a494324c2908879e2e1153942d084efa96b1b0134ce6d9896a966ca7c73a3177e77cc02562a87a34fa12c1aefd86e27d00e63cad997b8379aac119d5cf10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1140d4efb18cf5f15c8c17347d5e485ea8c67ef8fff601282577bcb3ad834e03c6a9b4b1e1cce7b4edb7de5c7b4cc7b22661fff2dd31e27e649fb98e2e4678263fabda54d860a94e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc1618931ea7a5dcf3faaad338f289207e604f4c698e28634321bace6f87294c52b00dc02af0a1232be07f90610ab73a39fcee641fdef5d5defd2359c62cf335cfcc5a365ce85a99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc90a532dcb521df2e45440c954ae3f296a90be2de9a43d103e1d72d8a7353410202b9ba0f9411e715cf59873a6599c41aa84abbc21236ef9215b17bda5b1b992ca5f98a5393a81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h317b71ccfc186f4ccf8aec2cd2ca642534a221e4a710a8ee77430959bb35a716d454f05c041af684533715c7d4728fc8b5db7e563dc1a13416a76defe11e76ce79208982bfaf9bf2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60a2e9042d2b345157c6dd19584ad9986dd6e7e1f3f0e478e761ee9bc285e7fd649675b23af2e861e295a08f2ff5c96da22e04f85efb70e1ddc909d9a4ba5dd373b88b20761941e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffa1e8a99e9d6ddec12d263ed5404d43bb1bce80781f9d27045728ca77a6e05b9530c57cd3ac412f6acddb00e596081ad0363d0774730c7db2fc80dd3989c485d3ea0bf36e3225b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h627796da79f5f3a1730c5627b088ec563deb931c23269e73ad6d64202abe0f81b41e06dfa8ce5af498800278f3d26116d6a55ce8885b14a112f1f78ac0cc2554f0f94778a2a8bdfc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ed70328b31d44cc8d56da636014800b67c3cd5d9f9fdd339b0bc79424b173900a51c7764d4a2a6c7f2eb708be645d6dff0bb84465c94853317826665ceff1f13b387ddc575d47b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb10cfe19314a0a3536562099eca937448a59042e2c3e54c5856e604ba306a01925dfcce6f10ef61cc7ad2aa76727962c8ee2935d41b81482b0def4d32191c187405a35e644b8f09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc7395b51cfafc82ae3de54a9dce7ddb403f9d1d8abf38c17c73b9d5a2a8c4b3b9407ee355ac20a8ea20fed737ba865d5aa674cdd9c5fd165714a5e0660b23c64d97a5e435ff4764;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbcea1d30426bd75bc0e06b823e50ebec1018d79b5c58c704213d9dd3d2891c9ae3402d159db8fa7ef99b8ef60a3707bcf9f7ca5b2661653db64ad13ab706172365648b9b8ffa5ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee5d79fc044cc1b08b42ee0deadc98239d2804d541a0c14f6fef1c51a98d8b6abc8dc698bc75c088923fdd2431e4e39a7b452228cdc93ec4f6db5a0376e7731e2303ea544f402c0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb71dc23b3c03496e3e5c3fd11fa356e9cff2cbf45d492c34d810cf4c075a08afc2bd7417844742d66060b51b3dec7881684014e266cc07ffbc5608e72332de2b05b9e781c9bcafa1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f488a2c796989a016bcb350e0a197730fdf2f0690a472b5ac4ef62fb81f8ecf8c5a6692d60ec8a91695e5b3c5c7bea3c8f94b8038a77af0bc02ca6a9954e46d0c54f9cedaad77b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h859c2c66044e3310c8e14a143cbb3577076c89e258ec7c8ee18b3adf83f431417ad97eccd6b4975b60c7607885e88a294c1f465998cbe7555ceeedd76ca92950f92f86c33719bc09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41c0a985ab14e607947290fbaed93588dc5f8e36891751490d4beb5a838c866af79d58fa2573b4dabee1abaafaa66e53e12df913039e9d772b9f54280baffc2ef94484261349bbf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f2deddc30cd75e2e369ccaf6862e6213718a052fa7425a70ea6cce92ee0f4d023678eb64c6df2b5fae38e60ca748e52b7e6d0feeb1fc836809aed9567e2c36e7005467f28c02e86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed02693dc86d2faf716d1be5b5f4f6802da03cb55e76fe58afd0549b55f5e65a2ee09bc9303f98aaa52ad0cc93af51313722cd1b4659085924ca434b61cebb8281241cb3501207fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60bc6351c4ab1c60573bf7b8e1b28496cf1ea0ea9bcbfaefa87664c63ae4ceb1d7a8ad4e3a0e2251e3ada176507851975319cae63a9733d78801a4715e9392ff366e046edde3d836;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf01918a661deb993d5500f427b4a9c539e5620a662486f0f2383b81ea2f000dea58c267b4606ab77fb71b366390bb42acfa3d7fb3077c854078269da899d2bcce6cb2b6e99905317;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf98aaae699ed31094ed45595d6dcd765050ffb043b70297d0136dc417be0b28a1d7e37bf1521f7171e6249a385f405a1851a3e001e2ab7115c4adb6e17081e3883291cb223df20c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6d3aaaa3ce80c17b5867cd18d9640e7a9863813016e8cc0a249327d91a3b1a2f960a31bfc26e182f666e6af78efbc24a5be080e7b5f272d834ea9fc170706b5a480aeef408b867b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cdbc8c98159d2033f0737e45626f422dbb9ae2658c3b3256bbe4c7b8871cb9179811d03543bc848750a3da9254b5ddd18f568bebeb4c584fe1351d03df8e54b05ca9feb371753b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c3d8d84c40a71ee2792676140dbaf6192a7c9cf6a59dd185f7b5ce3ba3bb9031bd591653dda71dbd16b7a190e7e161d8f852d0b51fce4b2a91329d6ee4e98ea86f41ecbd78be17e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdfdb39dac8500972b70113492c03805fe6bac68cc624e6f1ea4cb4e418d0b67c6186da3f87207cefa19711d6e124395719455cfa2cb5352480507f4a3c33f90de3cf5c09814149d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6647d7c9041ad6da9cb63421a734c570e585e4892e6510d12efd1d6a4481b024e639c28a2a420183cdc461fad700d9f9247a83d0c8d0c9f7049ac82a33d7e86733e06e698075ac3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19b8b228ee71c851d7868db201434a08b28cba61331262be173e1c5624c35fc0d00c4c6b1a30777e34ed878eee8d8cc0ba064e581c54c53c8d9e02207aa0140e3d0977cdd8f9e68d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc02086f859842c8c418a6815e2efe92c4fecaddc152b57267a4068f8d2f098424e1be82b80fa6da3c9a019e4251b1682f558cd5b697c543dafa14b2ad99a7397f812074cbb954cae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h450a4b014d48c1aec29f89df3103a8f0bcf666615aacf992c5171e0d0fafe27186782db879e75b834df400497c2c77e9b21abd2fd4c82665b46618d827557f11294ab62227d82e0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbd9a6dc9a89cfedf58ef3da38cc2bfbf1a9d8edd94384e5fdb5f6d05842fa201f1e21118f296ba8f8781c14db941623444774044fe6c51a465992a9fa8b6ccedc1432323bf16c3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he58020e0301e1bc28ad4bda7fe18ace3e77181e4236a18d16d66ae6acdfdfdf33ac2ac1bdfbefce3da723d7bedd50e393f7164bb4298a1fc7c22ce74ff415bf4e1500d65ebea57bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he488482a30a9c15980717e64feb8f9aff0c787bca9fca14d5a409b1546093dadfb131137d7b4b03a5bc0dfa6deb9ba723f16dd4ad8520243549fb02b7029aa9835b79db394a3f9c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he922c2579c515a55120a626b50d407869c1aada8c93ddb2cc0f6a8f1ed497138f5a1b4abef211223559002f7803f8f7d0f5fe761c2794a0193948be45edc824d04a69bd7bc6b09c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee53832c1dd14c2e785d5e9b8eb6d70d84cbcc39ac716cb04f5a0ee2ca68e179290c31ffe8d107c4efc299002908a28fab972b48bb2832a5994a2cc1b0098f768e91db6c1a6f6acf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbca170e87aa96b24cd9d6b576d16d9ede88859b66019f0578801c8dd46373e5075fc815fc9b8c6ab160f95252883113e7181c36354bb0c2dba5b02250ade2909636dcd557aa8e397;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85a0427c4af7b71746ea9855aa1ee4e86a85e06b5130106d77c89031553bdfee6e865da09b120bf06c110d2ba1e20c212a7f146f7d389c6ffb4920dd34ed86e29d0f37a8c4aaddce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95885b82b06df6d4c87357fab92eee84fca7f92302cc038949bcabe13b4c2509bf4837c80cd0cd1fcb06f25c1ee410aadf8ba06c180d8b863d9e29a4338d040256c425f7e6c8a95c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h355d98037c5e98ad3faf623fa8665d354a3533c003881e2f765e4ce66a8bb8d549c5e45e9ed687027f7ac3dce2cea6a1b2854f2fd01edb759a88c5902ca6237798885420547fa3ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h479fccc89a8f51c1f5783a99a29cfbf6e29ba9b24a17eb4f2cc38d8b6a412659565c45f53faf8093cad72deda486a3f2bd5df8b0129e6fbe76b4a0a372a2e08ca6aa793b47fb0c4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb565b422d15dd125a678f4d1b00bffaf7f918a32424231f13b61fc260a9127857fa6306efbd8b2806434fffe53e1038ec50fb5b682e64b7e144511cba4895d7f64090df74ae9b726;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5f9ecfb56fb316b893b45dac0e8f8e2840b7e1a5cd14a65a22b978a80841a7855dd0dd91acc1082c7fc6fa5cbaa9adfe63d7eed6620cecd5602d86701c408ae26eeb19bf3a7ee38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc5ff8088e0abd6246a5993aba9d26bb8fce1351a9343d4fb3b287dc04c02873aec09cceb3b6b29f959cbf8d7d651a75d04cb8f030e324c812da869cf8510598a8f825e9a7da76ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h689381e1c0f37ca0923a1148fe8b49b0eae820610950ef307efaf7bab245baf897106e2e8492cf7add34dbb44bc06914c1fb54356b22b911d25b6da56d1edfc06855395078ab43d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4aabe7cf1c3f0c09ae8a9018bc22572d6a741232f1fe9df025ea0deb260e454ecafa8850761dfafdaf07799930124f9992be5ff8dd8eb8fd5e58c3971f0f4d293962e9616c9f239f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h828a6bcb287c55eed7499c524a52c7d17039968dfc6a6581dd7e8dfcea98ea92d54f638fdb09fef1317e534c79cacd1fcb78ac5f242001fcb20668bb928b9b10ba8a0d03dc59bf0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd13396bebd4af47a826f23e1621a9b6ec4922e95ea71382953aee6a688fdf92f790b01b84d2217367ce8596309a5230e329e51871223913a44a213258dcc5af6b233757197afc322;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86049e8a5b4acfbfe0ea05afb8ce288427363b0b728f3b518e8641c463d7bbbbd9924e06ed8a4ae364beaaada22843601c91966eea87c92427c9e8edf9d1a1fcd4bb7acadd0c2e0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c292aa8317bb6419566fb9b6df48879ecfe77f46c96fc5115678ea1f06de9c168bd31222835b32dec407ca6910e53b11421cf72d3bcfdebf727acc4cf194d58872fa95100f7f1bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49646fe6e8f36329d013581a8c619f62ee6d7c4b74a0e9f4be2256302c41744d9a86e7966fdc145aa52631eaeec9e0590bab52cfca50724eab9aa5d42599cd5eab064eca3c2d152;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8eb28da02dfc01230fdd584e30f75e99af0106262e45bae3d08087141a5223bb175567ffece4d1d8a22a2e73a237c02e101b44c7f47034a075411274408e2742753e31d3c1b16214;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14bec80dd89207dca66a5a8d5fed7233a63ec890757c9f5787121c2862dc442117bbdcec6bdbe9cc5e69b1a45e96c4bef3e855835ed770100e10a5cec34d6cb121932a76d672b62a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62b2301bdfd3c62a1ca7cdbfeae301e48b50e8fddf278b7916c3f0c4f2cc0e6b49b8a8e648a27fafe94bf9dac7484c1a05a016a2d85771adbdd03aac21b7b7cb79aef12a94705173;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha38b3198cb26910899115e38d5854dc61b1d433be9a46e5b26e6df760394e9a90c7f6f0c4c15748e6956ee7acbda8b0db5e1233cc05e4edda912a4f39bfb4f8879db9945092f6f87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e70163f0e72dc03d345108d9ae7a7a89994227a794222fc45de9158931a82a02c0323b8fbf49899002239a84409f594ff0666dc1961e9a4fb678a494af57917bf1650cfee26355a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46b6de60d4b2ae0e80b9be01b137a5e50ca6c9d7ffcbe571a077eb5e62348cfcd61c38de3e1b9866b11f2c28f7d83cf3a336725df5cead5dce1fa216daf7bca50e58cb243b7b6262;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ba67284eba32f11699a9df42dcdc1789a8f52235d874f30c8a28f13b6d8117e542261265b0aaffab585f679b6e8b72592a86638cfbe7e5914e9d879d7fc740275b107d9f6c69ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd21f4a70151e8ee1c3f7b41b6bf06bbbbc770146d8946cb9919d15659bc7ffb80b4e58fec7566952f88fd7fcbc049cbeaccc704e9b8fc757419c0c2c66a0f69b2745bd063e90fad4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23346bdd761ff5e4664758ee7642912989663b8ed7102cab7475cb3be86df0fdfdf30e05dfe82493365d01f7dcae5734c9f3b2fbfd1ad39828d62e47e7aa9658db3a4c231e78a503;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25d0050e1f10ed12f9859c5c87c10e1633bb93146907c977bf7bb35370e61767db5af47f66f673c985243a0a6eeb95027603815f0e7927d1d41f3cad48596f40dee654460f42296;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hece29de5eeba06234269507f0b923c8f318d1fe63b5fd4032c3cc047bfb9b0281c6d4319c4a7a6d19963bdc35a1dd5386109a628a7a5c748f0e2edc2ad71489e815368942460f378;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba608a7fd435d883eb559b3dbce1eb03f3d2f3c8ed474a3060ebb0b56bdc1a9d2ca38b3360398f70dd5c3c6602cf6f863f8681582163c986113ca2eb7b88ebb0fa7f3cbbe5e89223;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8ed63842527c45f5b05a474f9c3baf32d1d130ce889961d37ae84e64db71317af5812ec707569b374274972e2b26c4cea22017f034ccd5ffe581edf4b0a0298ac7a88043a1cc43e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed7c17d0c8e2403209ff75953dcfa4c1f69783f1a405eda1e6905e8220cb53cfa9e771b518271481d1a14f377fb77323438d058d657338c16c7118e80a11fb616fdde87821cccffb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4917cb41cd33b87548aa0552b5cae55bb22e1d3175f6939f36d4e073ceeaeb52e8add362bc29577c02c0262d22e094042b58659f8df6138ab6a82d42b23b487186d08a8221c9e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ec002516cf3356cedd7530c934bdee996a34f6fa479f9aec72aa9b0b68d225b08228efd2ba8fa7233ab3ef1fb9ca72c90243722fcc2128a528f5c735d439d1dd8bfb590719536d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc89c6b0f231b2bddfb45646099ef7b6c822a63e426462d33ca52f01e2efc3c222b0218f84f3598114c8a820d852fa4d62ec37ff72006aebc658dfbf11f73701f1e57a487ad9e525;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14740142606529775bd9d72344fd9c21098c45173c2bd0181b9796182d312391cf2fdcd2727acdf5e25cbb73aba45a8f3da20c815be6f570efd2e516b462a264b9356b3f9ae7980a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde02e33fc29866f92a56c474afbe8c8f3df170a7487fbbe15171e4282e7840771cdac74a7951b323034f128b69b990976202352808ac5988098ac4381f60fe952a67877646379d4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f57567d359aac6dd74ba2c96febf9ddba2bcbd010699dab8dc4a393102faec879d2cb6f3f397fe76731ef3d2a9d9eab712ef6aa1d14c67fb5baa971fd88bf9d054075af9b9dac28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa132ebc221f69a4f5360e7465f6afc695dbba7a1854b902860b5516ba669441785fa5d4ef48cd99fec8176938827025de29d0a553c60e64df66f9a2b7497a88c558f517cb2d6b98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21668795718e48ffcfc3ddd9e59841e85697404de392133d465c5cbe6799d44a3ab55f57686a4d9ca05c208d55ef15594673cc77ac48890dc10833fe626b50b9be2805092289bc6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd586d7f373ece14503ba0e579e1c693aaa002fa9ac8d544b375d48fa583274a13361ce4744835ca12adb40169ad036d7fd9307d80def815eb93adad9610dcc97bdd4f5feab085dc3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h623d672e044961b8bcb7ae6056048a5c120f41a4c29ae7c97cbd1125909acfadfbe1570498a75718b087dc5812eb4846a3bff347ea8799e8fa572d77230ecbffc5f291f07009efd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ccc4ee4534ca330ed29e6a41e4dc7684412fcc0b80d30ecace72c2ad00ff58a7ec93d4b0f00d34a6d9b6c6efbb0c36eed4b76ef97a9e7e3a013666cf70568c0a566e2df70313bf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a148b87a89876ddde04801a6100db3553a0d083a6a63e17d1b923325503d619d39fd15c1a23d6e0464b9a5eb30f39b611bd07c2dee97e9e245afc87b0cc2a33a66c82b3f1d1502;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ba995f907d32299c479a69d7f02bbc71be1427748d5bdb60e504cbdfa70623c65ec0a6d76e53044808a1c3487fe90962ba1f2fd3d084453e2650f84047fa6870e5df392bcfe360e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa526d379c27e64d73b2251705a6e16d0e9d0ce8c5808753411b40984496c2e9341d6ee563efc2a1bc253f40ed3610250b48238f4420f230e4694937972c70f0cca6dd05852a06ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3be332fed54aa464896532c030372ff4f1e1ec17d7a86477c74e9bbfdf338490fc597767d6e3bd6edbe5b33b6be2c8fd882d2fe969789baab6416f64905d17bfccc63da44627874;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h372c0db486d28f75f963def7a68026791e35463b8a0de259adf83d7b08bc5d04c0043a6523f05ae91fd929fab18596b114999f9cb0cc15cae0b07c592729bb690d8f1239009fed9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a0ed4ac83af9f228bb92bf5443c0fbd472bdb57155b34b611540ccbb832ec2877fc78a1e04151df9693704fbcc6d0f92841195c1a8ed159a82830c2baf94a0041d6e9590130517e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91d9b289397daaddc7d50f162a70582adbc50541000cf489487dbc1137bdec8aa42b025cf2a4f9eb48bb653b68b6522f3effcf47012fb47cf17968a3d87d26a1b0832377d9edf00e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he10ecc52566b3975c6687a653fe7352064460ebe8a5164df8e830dd1744a1bfdf1369335e11d9c9c90d9fd6c37ccec695bd12c335a3710122f2e43ac73ef39ba8f18370eb8c0eaa5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c519981f78c3479da9a50e3d927e4b01996580df2842782c951aa0ccde449ca807626a045736b106e4a0457f5e187748ceff9ee34b59dc5354d1d31947f55dcabfaaab290f38ba1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha256a77b7a4862afb1d8b36df78b3addda6efc7696218b0e4cb5a8ad5993d8392676294cf0faab1fe9668083e55c28d494d62c7f119d0b9352ca40d9779499399d605f4222ed8423;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64ca35c82b98b671289e97e21ac02cd2d01770dc6613b36a0bafba24cea30b05ea482222ddf9c1f677a2d7e9b59757dc0f87c560485f39b303c62b0138a8cd7ae05ccc16db58f130;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebb24402afc813e4041a6d5652f32acb688996ceacc12daad75cf229c027d7f432496398f0251f3ca91939095e4e328e3d4e1012415e2930dd3d1baa487fe4bdff3638ee9424a47a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2975aeabc5cc93a7fdc4b0561fa612d45c0efa3c0e6b2e87456d84466a195f508de6cc763936d691c88622cfc51ab2e5d7fdc60a4160430650410ea48ac5aa7682b7afc3d4d6e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb908903ad4300626d3ec699d20b67352feeac0ff429f1ae175d72ff2460a664eabdef55506aeae470d74e69a2a360bc942ebb4df5062def4a892fefbe8fa21c58e337f228ff9e9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6bb4b37dfef0322a8a039ea1e4f1d124162ae9df6162732a4c9cfec482bbeaf8e04abe83bf44e87122aea5232e369c7ab2946712d1d7a65a53d2f7dacec7d1e5f057d9e265c1555;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h216f4404d376223d7eff7471202abe47a493f34409453cd6ed5dbc0885e7bfdcea787de84a02ce19274fac2dc6fca309ca5a8929ac4069ad2cc78e22146ae2c9357bb9f900843e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb18b6cbbf604b4750976e295f82572287083cd02f5435b59cbf98de1e1c3511304b1b49de6a3c11b684fea8f09209a9630f641ae8d332a05fac969b3e4abe728dc7920bb6286e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h878e2b20bc25d2f9a2e45b13621b4bd4ff7b37658b53fed8ee6ef5da23357fe548fa34890a73dd129a7a82da2faa21a746d777bb42cfd7a338273498ea835f674afd543b4b309260;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf01fe528634529e616f274c1529d910364ea446698f07ca8b01ebdeafcb1d12643a5f0f68fbb0f1ad18af01e6786aa2a1c997a4e431192090e0bc1618fa7114d8c653e25d955257b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba5a9cf421369a90dbf387c758e899ae8c8f308b2a40122af350096ec3c63097e55982f18839f2f0130602911ccf318fce4ab815a3203a70ba77819c15c92eddbd53091051e97435;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2e16d9232bccc9110ad5b3c71f1205adad2142577cd19d085d42543de42aa538d3cb5f8f46088325ad9c0fb1d15dc1423b708af4dde1e086bdd1d8d52653c63b3dbb5993661a3b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5209b56ae15036da6ffc30fc4d45a9803da7e43a47266788c8f03d31ad8483a2e59893ba686057da6e4340110b9f5dd0782e033c36093b880cf1294d5806661ac855649f746ced2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73438e34d17cfda69922a03af1c64fe3b19330cd8c53ca024ad76f994370b0d4f7f5360ee96420a3977d0ff304da58ad97cc8ea1fd51c0865c9af75a8028c80f781e8188a01a4589;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he85a5101ee133412282331edb3cddb1d0f7a2a8f021af62d9def103bd3eb1d4b5daca20ff99d782245f3e7419c8d7f06fe43b2a3b4c22aef12cca151d644086297b20352366c52a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedd8cc61eb0bd2921a1198b29b283a11493a102883575b9cd01da6061c4f5edde4d03ece1cb05652a1d30ff937ee6cb3d7fbb1e06fb2657ccfad0e94bc901bdb0d7e495711a56c5c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb20239dc5cdc44e0c403892f2f1a567bae28967905e4263b4cfe761a8548d8824c45c5ddf5e3a03b5eddff6dfea54d58417572cd24c3739867ae0443759a53a832273883d20857db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h601f253a782eee553ff83d65c7cca0d3c361f216175fb91f17e6189be481a09788b479e4f69e3890f14a1eb6787b349d1499ce45824bab95bd4a9f13a468dc86cc3e84a7dd41e1a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h524924bf4c729b3e197fa8840d6ae9ebe3e89e9fea8534b485418c41f594caa46fab55ba5297ad9d28cebbebfc121d776860059ce65c1a572e7ae6abefe36b8bab83de65626bc93e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf51d8a6a61db930439f5e2b90db8d3146ec85e4ea3773f740c18a7830965a9935ae67bbe21b57316ceaf33cda96dc944769aa5349fcebe25129d93193feb9b304fec15d8be7979c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bb16991e67af967d6ee0e2274b265346c05ebd9664b88665cff804d39b71678ff85a72fc6d5ec39c121a3f8e6f4b8a99ac7189b3c180dc805658940da88841b0f96776039b82e4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h872bd5acfc5945c1fbb2880b345720db0e433e9973baa24ab5dabfe3fdb37945a72825349362ace3e11f373cd51fdc0dbba8f1fbcb05b0311de01cea40a041c82021571b9fc3f691;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h854274ac1b996ed4b9f058148da319ac8f6d1250ca70e0cff89f529f154c45aa3c1f0f350258037198dbac222c9e66dd65eb55a5c46c0783f7fd4c23b1debe4c9f81ba872a3cc4ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb43b1857beea4b7ee5475d85906d2692d883dfdfc6a63debc9ec43b98cb98ec901d2484b8b0745d8fac63d21b876f07249449664590f0191a09f38c98e4788d30191c9ce11d3498;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d4605340d5204fc73e3255a3e71ce1b6f9d8758c7de3f292895c91bd5d1eba0adaed36b22ddf19511256164ee6dca1b861780248332d748c13bd633026c9e6fa25dcb70383f77cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa6edb5a26f66efbe7cf303640cb0fe7068e6e45a91f797946715a77a789fa68297e86304c63804b3419a588707b8f0a393a2cbb3c0abbfc152459b76f71ffcced2a58c497020163;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4972e01d56d0114adcbd7ab82c99e110f6469b7fd4ee9e005001fe5aaca9a598f690f725eac6a5ec0b8893752df1e06826e4ef4c24d6ca73c3047378f2b6ac55bde5d19eba79c2ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43b32cb5ffa2aeb78859b161f8ebafa0b10bb5e84c5f210b2c84e677e7e94cd31e5003fa4d9bc71f33e1eefc2c72927f4c9402e60c7c79f5110d7f07441907b715999e410fe53def;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heba8021b988d40220bd273874dacb59a411c15dfc0466c05f0612400dd2ccc60c816b2bd16a1af4bef68e2ef1c38933b7b4d35b25c249c8a6021f4f6c151d860a9c528ebb82e1d5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc77a06eb9c630d0b95b8266fc6a2581ef789f238ec3d770d75f4dd18c664dc8effba27977486eb6b60dace1cfdf52fcde4d37d32d1d354c00eb72fc781144b3e2066d8fd835d5dbd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf97b863282d3f93f12af2dc0fedabb5aee0f7f0ee7c2b3eeb282678754c35a7de86fc2becd4ba7d8b4fafa479e40f7e4b5b5207532c19c72d5c85748cb8a37b9b232387e9bd97fb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9ed9d53b4a3e7c0c2cbb5560cab52ba1200f83dfede41ba58fb43e67e7ae489b0bf17da6e937587bdbf43bbd4d89eeb056faea04b98c6ac4232dc6ec15a17a790fc83da9ed16905;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba9be94d440db162961336d24a9c1b3867f18240816dc0f810125211a978f9ba20fc897a384dafc2e41b10971fb4f100587f5d1fdfcb11164457203bf933e8acf6400d5d66883237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3203a30eb2e991fe255a2be10d49c35ad8910a66953c0145da147c477dd2e34178547f41ac6b3173524db697697b8b4d7aff8381e11fda13f46f637e487da97cc0fc37ac77aac69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40c33b09d822fa3f5fdfbc369abcd991e7fb6a9a4ef577199e5bebb0ef2c60458e66811dad1e17820cabb9de0c0ebd6ec00877e99479d39adf36063ab2f5092ed57a7da9ae2bc6e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb62ac9a43c250d9f971c7f661a944f8daa060e8120fd93fdd0d5b9c47537a4c0b731c6b56e968123b76d64a384a99f5e85905a9c006034ef1d1434d92bd913a7de5049f2d8b06a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h718766fbdb7cd023f43593047cbf185df15131236421ffc0e2b2d6df3736a1170295b99565e2bf2998f3fd0a570d2e8f67e286295d7783cbe3b6c2f946969cf391b759a915140caa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98184aed1c207790fbf62444e4baff713bf35e88409d5eef8e86ba8f23544bd8b25e83ac1b0adb82281b56525f70f116559be5fe20c323d92443da346dec0c3a95954362a7a8ff4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78be5bb7f7a8bc5ec865ee066e2d6e5cf01481062c60d77de7e0ea7322c3afc87aed6fee5552edaf1409a8423514b7f7f23bca7f22906de0d2fe0c6d8d85ac914ee7b20f83ab95ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57ced75bb093a30a1bb78a9e6b6de72f0a2b04d193b16b0023129215efe3b6aa92a19e85d0d79ff29abff359f3bd0765b1947f830567079f470859e2a73c8e30ba6ed258f5f60520;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c203eed49dfeafde706c32bcfd709e6451167a83606c2253cc275f781c16506972232dbafc55f6519d55dcee4059fd2c296046e2cb742c7b3442d030fce4ae69710f4c2095971ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e1fd738a0a3689f36b3645f53921c0299f08b6299e2c329d87064af391b4c78d9613ed7c4a8c15dff486fe1840f28e179f3ebcee614a561b6219c55b2e237941fb4d29a7a7cb3e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35646d772255bac33f02b4fa68973c9375051e4c9f64fe5aba3b46626d5691857141284560361a90e08999ab27cb62b002578a5bda80abf4af92f87caf38b744c5a2c8523eab3346;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he326d560e4eac588d08b6dd80d24b8982528ec00937be943c487f273169329d99d60f27811c5672e307bfb12eb83a2a39056fcbbc7f04a0d34c3823ffd127994b3369f3b1be2269b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3f296f3262076a37223ce093714d31920959f68c01b48195a15315f9062654f9d458470ebf86e0268be2b3286a1ab5858d075725215bc2a513c2fac09588bd1c9921627ea33bae4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6480d4d37e84d215f9763b7278ba35eeb809e1dc4c6c1587f2f949c2294802c1041a9a680bb71886599860dfefa72e9e91f18c18e8c2ad9e4ad2426b1b45ed505831caa23f116102;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2026d6cc1686e43d05e9bb2ccb9dcc928192ff1e028219472bdfdeca9f535047cd16f97857f84ec5153c9fef2a1e0c1b1957e11f3eecdbb6f648b4c4e0b3e0cd12df4fc06c246f0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h302fdbf16c14cd7c2409ca2532fcbea83e3002ab46dbf5d0e7c2bd6c092ca5b8518715a907ab685d032cd99615884099de9205be3a78bef8c94fa97c81ae3b8630e8763d11ecda45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3694c41cfe4bccccb16ba8d7f38540d2abf01929be1e062cca77e09c6676ecb87176cce1f607ea91715e71ba0bfdbe40c1fe0f436b60c58385b8af4571d855f4097edee8f3f68bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha85dbfa2c647e819ad58224e64a79995e8e9565bda60f112f6017a00014bffe75a0025336c9203949ad94a3bba005cbcedf9ac927a38b57725aef74e02a9970f4306295fa47c489f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f639ba7d2e54372d9d04c84eda6bf0e3cdfd8910cf33e65b197de4647b74820a54123d3444fb5bbf8719cbe4143693c5de8275e71a6d4d7bc0a41dc182b04e98a8018fa61b49315;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb76be69dcd32aa03bdc558f439aca66a3ab069147e298e8eb1a2c2cb7e4c1497243b50af8491fd34f7472d13d971ce117bed5db6791a9e64516a604c065a912f7eccdcfab9b98ad2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2547564cb364a5662ddf537ffaa58841909005b68d66d6edd911cca477a1765fdb5caf65f403bef3399c9b9c1d7e84f74bf39aed26ed5b1c29c9e9fdcd9bd9903827f2dc95b13cc9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h212248c4727a1a6d503e6eb28d310b194dd6dc0d489e61ca96d1213601c7fb4738678f2d4aa3c1376cc9fcaa57a42c5648252767d876df48180426fc4831745ad9ecb653878b29ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h422d5dcd6f074cb0309f5fbec250d556727e43016e14d1a6ba1182f04798c2b608db1a3d0e6e5cd204422dd0b817925835a270a23343df2f86f2a547ef9fb380406716f995dd914c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h873c6c943275a6350fa8b7da1283b1d4aba7e5f27864a893f41ce3ce31c00df013be5a517a0b7f8c51f4e0bd6fb6475ab45dea77fef37f717034a696c2157c1f55a470e011f7abd7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb5ab69f719eb248a84d8b5d7295c9eed4d16f026e4023e046962045ce30a2fe53a54ad166bcac1c69bd14ea3b363f173dc333926d45974e6da1d94b59f610d3fbf4f5a542d72283;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23ba1fa32bb2c3230618b478ef8da84c4e4ba99d540436c67c032af641c98115d0337c1fbe3ef8c5907fb547fde92ddf6dbeeb4a1046c2804103eb2e393f93c4e358de37fb85bec9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbe8ad8649799505e891ba344e9ca99b1aa48d72228c908e731f862a445c4ffb8123b4d142a50852af4aca694a35a07e623698e2e4f41b2d7c2b5ed8c24ae9173a97dd99513a9cb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb554ce2a07377452563f962c396894c15cee4c13391be7e8045d953315f1cf6e769d33a48c0f12fbed29bec4b98339f0b048fe5a82c9691f719f54f7029efaa97115e3ce870a4880;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h796745f9249d5274a526b7245b8fd4fb49fa3d5419ac6ba85fe9cb1d0f825ec3467ce6c5c5893c0bf61b9da910284719ab8bec2d551550dcab1a306b6c81d16933f912aa8c474404;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51fd3f0aca16ee697fd646f493c4dca06a2e14e4f503cfb053b923cf2c9ff507a1da4f0915bac0ce4df86fbc7a80f204c5e9b9d19a29ab74f139fc045f3864fe7ec8c56964ee4bdd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3f634b0698d9eaf22863d4fbdae87f042885267603c009d6c5519e027ec9d5fcceef1ab48d1d8471fb3abd4e4ec4554c7e485ff0c5779c7c04896c4123fddc0105a541bf7970670;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h868a7e5b8be46976e020b22e75c0acb37329b3aa14823d555777fa5f825b61ca42bd6822d4a3734077a41e6f8c5c2a8f2aef8654bc891fd3a38e3bea51989e9c5b12f3a6803f79ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb12a69513f51f893c68941e67b72a441ad6383e3d5d63ae3cd234f683c956d366502f0aad0a82eb07ef22cdea0a18df0351283cbd8b12cadd6428e881b4316dd7a4cd5bd29283549;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60e5b90a9ebc4b8e2c2def37594f08b93d3ab3298dec00d3f7c7e15145b4ef215919986339657330adc7347b52608128c71aa375d8b47ac93a978041b7b0075a86b1503003e33c97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48a9c0692f0f4a354f28a59cf3cfd0b79686ac98fbe23b253d6fcb9ee62f1a339c9993fa51a2c1ad6c439fcb2731c39b0aa937a3c10c2c1434ba45f69d3f001524cbe0f759a720e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cb636d38b69cc6f0f1d0416967b3a0215cd898abc346037d8d805c917f2bde984aca6903e69b24dc331144df4fbe8c3a6289a93dc9576af04ce34605d8246ac9043c7c5403872b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef13b795021f49f1193b838edc1e57fc5ca801f2ec3bc6ed26ea11bcd7be7f474a865e90cdfdbc05ba47adb788d59b75bad437e0ae4805766883536183e1d4e0c7a7f4de6df8c51f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbb2ae8f7c9ed8d8e662204cdca7ffadd22ef23f43a2f5e2dfb9077d5f95667be33d53e851768598411f28edeea3626e04189dd979f00387f9cff9ce426060536f925db968ba4414;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbecf7d7d634e1397ec30460434be950cc516b8517a969e5530bcbb0f900eec1f3bfdf57f409207b2226cd719963c9c92e7002e4f3694ad74352ad1cbb178b9f37cc32297a0972008;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadf4a4b70a86c7ff60ac0c9a21bc2eac90e4fae1ec51514fe95862fa74b625d4150cb110a3bf1030da58c84e4d4f9b867164b3c60e3a249c1006aa8c1ea5be491764cd480c321b47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94423cfb1d125b3d3b4bc970655c9de882ebde0fc3de970db22949eced3e3818ed2fff17601fa4062f2477af445de1c432f585b7094c17445fcc99a60c6af1967fd8de7a21842a72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b091687455d16bf788a461afc681f57ac140294e7040de8dbec09da5b69ae81a356f0c97c30c3880068b4adbd214d3ad1b9012da3ad8a44317bb889003af8fb7f0f9267ce6988f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ffe980f9a5c2a0df68039e6c76eeb13962ba1e28c00d4026dd56803454d61b5072f5cb6a09787f1091706b5c57016e48dec35e31c35237411f41ded3081997dc4d424a5fc1f5a2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f94ab16e1bba4f4d0faceee4c4db69bb3a9111c6755979d06cfa30589b813f0a3bd0ffc65c4d31b1cd1a4905ac90f9bded39bc5b20215342591bbc7d97ae86321b117c58ca8a189;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6db9ee2602a16eeab62703c94adec526971a3a9c118d8ef7b1c1b21c8563440c84aa82762270685b792e0d765832ad8c4648bb41c4dcca6d45f27a26a9b880f491f70c9c757e7446;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf55b0069f1e4a9dfa11482a954c51cd3602a96cafe8fc6c27f34d49a29303db8b3916ff2290c7d88bd41151d1651ec6ce478df26c7b1a0697dfc1ace3831da8626567478c550b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6de699270dfaad11e8f3eb1e1d10f22abf459f352bb0c010481ef43f04a3d96961cfac469e0429ce8418aee854806e809e926abc8dd9e559e7bfae3f817430a3e9feed2fb71f0a3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd66b806517dc74781bcd033c3cab2cb693e0d25b73576ae266bf91ef5817ef8acfe48eb4d6f2560d94bc85eb4eacd07e0c108847996c0e3214aa26b9bb3be3645dc86a25cf68900d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6505692d9d9ec1cfe0612a5d287a42c9f29629225ee4385151a1812db0bef7dc143322d701c1666a992b55decc118dde0924c9926e1cf8bf0616837dec0c297c7cbc9891d4bc50e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e99013f5d5f80c2c42de14b2c58a947626af2812fc5f34dc24e1a1e67088d619e64a2bfb6d97ce4113770139583f3f9b3dbaf4b80ce31970a3596e6cf195ffc6f661b42237fd5d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h207b2b4344c925a532cafa75cb6f7ae105029a2ecd0bada395a5ca68f7e1498d6e06b03030e994fa146c6353f8669620c5011ff3412b6a6be4085f30f0e3616760fbc13b4402478;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h181fcba0f501b6ace75bc80e4b84584b2d93efe6fa89ddc1f31ef680706e8171b0a8ab1352bc2266a1be37099f0512b764aa39da0f7b48e690b6cda970cd9c6a5f75fbcd3cf40f3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd029ea8959559a33b03ad7f075a9a0e840ceb25300b9d8abb543cbbefcaaac30ae08b554b5c0cdcc4d44720bb860adef208b9c008a4c5cbfeae2f7c84c0c16d01712b2285cab3583;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49a395640801e936f07763f2f2c88b41119c031ab92a81df208adefddd2c98db73a8262eafc3fea9f8aec891ecac0c146ad41b58990a2f4a86905f45958040d29a80ecb6217581fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd54d5b76480eca76c3d772fbacf92a0d5063c245f84865df848237c420ca3ef4e7569accd797ace0bae76faa43eb91c08ba482c92a6bdfb6ff64c2904edf03773c1ead34085ea818;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a829313187cf395430f965ad9964d2a33fe9e1e0b95b5c008554c92e78d9ddfae1503850081961c7ab2e555f47f1d98e1e8decc22bca4fbaf409bc70106a0e034972f6b80345953;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9aa71366525b5eea401e883d39d48596064649979bc4746cd3671d58975cbb93ecb8819a71f72ce9cd09dede6cc0b58bcf8f6112b3ebe7f616827b964b8cbb013b0b06b48701539b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68bd81f51026f9994efe4b014872dbf0175feff92aeb00eddb0d4eb73cfc8d0787d37d9013c275fc4f6d3b6ea742124de6da43b54d314957fc5be71a27eae360b3cea62badf787d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a19d74abbe2d9b0d33c3404a8f46523d596a723672c3dfa9046327c2ee1ddd7373489e4c9c4edee7e686cbdcffdbe13a88ff7e2485c4715f69407b480ff7c86dc0d735c754508e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5ea0dbc18a9594d06029cb765a3a0a618e5a610b63485f287fba16e0fbe4865b12905a4664cf9839c3b64b03316ea3c87f78b6b23e6dd1094be787bc6748b8b4aced21afe932701;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23c85b389ef019cd9c246aabfdf5f3ee44d04aed6b3ad675856dd87b88c85b4d66d9509800a832f359c5c14830e82f8b37a20d5781dd96bae10aa6c121ef8b56405370e4a9279965;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb73de38affed4dc56b1ab63fd36594b6b28ab8920cae55c9873e6c8421e59925e11d17835b971259c642d8c6c4eb6faee0ba1c94390d132e624cc02f75366604785e5ae2c2b7d346;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedbcc3bb688b79b367b5d8330efc91042dc7fcccf61da4b872c4d13ca950e3a10a5f2d0bdfa71ae5883a042fe8c4c1fcc78cf7d1fb6c36df60864de4cc35de2fe44d38663d08d5ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f79ec93f5970eef32e3c91879cdea5f0c0b8ea667cebe21a54a82df91d249e0a097df63d8098a195ba40fde4106b9dd8b93bfb4062a4c123f8e1cfba7b96d432110f21cd83ccada;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h823d7164eecb4485307822b86838914e89bbfbfb8f4ec79b86dc75440e100b823c6337849ed60bdab2951d58344e88c1469e45b322d5f295d43b4a295cc95dae60fe84bcdc30c647;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd50faae10ed00d47c91d3ad5fd6af0c997d35efa56a76552399eb32e1248307daa11f49cf26441bb1881ad3b8a39032beb563d5bb641cb5994b3cc21f3a2ac18ba11a88c6fb51828;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87460251bb0dd9da9d57d96b4ae987fd739e7a9d90ae06621e22b1d0664c2ac665ea83b524c193496329d010dccf2aed32ebce8555d2c5bd91f9859ebba596aac6c84853c3c55f7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e61a81eddd81eeae0541b14b520b8115cfb2d90a5984d1fe532d468380ee3353f078b14fa14d395458343ba29038d34336cff3bc4dab36515bda89a146067584a385580eb31719f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba93bd2ea5cd00e7986f163b73b0f707d91ade12f3005b338c3b8de42f8cd4885c6937d980bb69b1d65964ea4da51418f6c10c22989bc6977a2368569d4200be3b036567cf11b842;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fe9a3846d7154896ef24da7a20c2b9e9f042a917f44207147008d9e505e1f143c2811b76151e4ab5e675f31a8fe6f2eb4233cd49642e064f4c3b38dd667819ede092d8b3cf78fe0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h625f8cae96b119e18a498466e04e8fcaa744a8adaf09555fbc84a83c60bd25e5fe2d00c53c2c19b89b9e3723f42cbe3ebde5527010ae0d57ef15489ab477c62084e19e8ddf8d4647;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h182443d490109f647e91bafc1745141f9c4d27c4141932198779ce95b132a59c7c4e70b2db34b40f09d051fa8411993bdeb08db9617a6044a7785398d93b4ece919d5c25d82afef8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e9e36403c9d4cd08f06c3116bc0e6f26a59def85dc942944cdba7ea3822cad38e8b7f889ba0a36921518fe1663e1c203373454a677d39113423e1f3f428248998f10422aab53f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h100f1977fac924f6ef689ed6be87014fe2f1972d2a3aef93994a425426bc5aca73566d9a00dfbca973743b3a983279dbe550c4cbf481939e7eb32c9b5f57735206cda162c40d401b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26ecfffe91ff1f65048e89391beffd2cf6c054dd9ef2a2ba32c09d742b8c7679b7c0592c47e4f6f95b2b21fa00d16280614233434c8cbc5d16976780debfe267389ea5366f9be18c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44b3768ad7f3714d3e4a98dd5c96b1f356ca0a1043066299ed99c7426a271d23108d2da8604f07a483b9cd3d02608da82bfe17738095f330f9fca73b7e5f4bcf643f6f8c2d53f3b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69801f2a59faf6c6ee193bff577e467f182ecc9d268f4e19032bb43defb8b191c4425d6f75c1999a91be649be5beeba041d741dfe2c5f8d3334f191790b680241965372a2e80d3d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65e66e5b90d8d70a5bae16bf81678f3c19e6799da2e6879d02ebac1e59d63db3b897d21ad4e80be43eda982bf1c3608178b659a0744150617bcb2d1e3aa64909ff193ba979c4eca8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5914706eabc8b844b77f5bfffd0ddd3149d2cee7c22ed21a153b7891619d8ea563029437bf3b523bee2286f8a06c33b859da641f1d491e2976371d444e1c2c84871486ae095a5fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9c33b840f9a78ddf2336ace9a1a540edc5d07665a9f205ad43a3f01a81aa662250e17ce3a05c090fc670db6aafaa5ecacc0c3ea3b92e9c338800d65d0d2331ed539ab6f2f16898c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92a879874f4fe74d713368454d975142e969068a48c4f4415fe184b27223f1e8b66b126e5a58fcce4012aa953ab05697d49933a26dc29261d31e25e4c58ed410c005991bc6fab6a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77008594d34ccc53846dca202bbba85c09df4d16dc93c91ee3ef1f41f054b151d018e575ba5baa260b8eb25793c1a58963241febcb05a2db70073448d70a253b5f7104b5ea74fd97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13b8ddd3326c523d7bf35a554a0dd7e3e0b8180d51ba565ba12abe4f40cf1619f5c0c169268dd99e8edbefa6b22055b6fa8c378e03b295347118ff5c8a5d776408f1aa268e73f240;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf87e880910390552b21964bdae9955461603720b400849a2c24a9bde35e68bf638ea24f37a82d03b685b12182dc8b8a38b059001b628dd397e4736f3f67c867991634d40bcb59093;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55dd8339a0bbd09e477cbc2304895178d6c3b072911a8f067b1bc6097ce042387259d0f1776ab71d8d9cf1e8c7fe39eca3031ced82360b30221be9cf380244c705884eff2af0cc39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31a962c48c1e1cc34f2ce28fa1f7364e57df81248d78c3d2cc7a642df7e255804ee9a054a2c70694a635772d9cb744eb7583ad5135ae0bfc415c298cb46b30bd0f30a622976bca04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd07a6671d1cf16a18ce2919c799a7fb9e3857d975e9325d40cd251d4ae309758f72b1ca13b9f9695028e85988e38f2a771afc39494fdd408d3e22822ae56a60b11bbb5d9f8d6522e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had34a59c4f8e7c10c1449a03003389f5b0012f4845606bac9bcbe2904d37a2214709b21b555efff7b4b8ac13fc5c615290ccf7c61e01cb6fc240075a03872d820e42c865dedf04fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc62eaa46de4543e61d9c57ba3c04293a156b24779525bd1e41f687cd12d27c5bec32b7f2cd3cd78e29ed0af81c7d53dc3abe81be2932eb093c78ceab2f3284552f38ef4d3a9cd254;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7df47b4e7383ceaaf2daa6f177f77894bbb5f05349997984f5b3860f82faff7877f924d9c9ec8c31e89c51626722be090502d5d1b9111d2033abbc07415e12af401efcb799a8c91b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc76032efcc280b8d119e90e3c3e2aa21a51a9f401b882c46162b40b0d72737e3edf0ae8b1175a77df58a642248b02ec6a33c3bb22c7938aa8cd7a42301af18b137654c9398c7e55b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45adc2a69ba2e18be1cd5b9ea02a8c25bb5009c7438888142f7a4612d01a0c7d7e4c9cf6ce51154e0d6f26ba5899cb1c8ad9c927bf265ab6374a1ad5f95fae08c39d6daabd8a3cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8718d3f95c1bac01794969a32d0139a3c0a5a147088d8b5f38c85182eafba29d10c5e8cc91d4bf87e9c84a8527f738d7bedb996ee003d1050557a07b012282a9ab095c3d2ca0341;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h583c6b304613ce36f0f00ac7ff47b68ea1a007630884059274afe30d0e9310ec250e4e3af6f6d2d0ba9da90fb6345c05e9e792d6f15f0e0f3c00ebfcafee074c30beaad7bfa01c2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b53d552954748f2e85f5d3106295cf548572f0650428af990bbb5d52bee52ca19fdd13727c37be7e0e0da0f86b7b3fc7df1709238cce0de825fb6e7e105756159b9cbdbd32c9210;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3488223bd49b86ca7675d87a66a9f6d3109d315d51112337640129388b68af8620d0217be891cc4d5e3bda77b9081f9769f9317d29f034353663b37a1331fbb0012bbc2c3b321cb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83b7d6e0a9840aba882c3ee7214db4a308a34e7c7586cc8b39f3d5b41ffc35c043733fec971daf9c77f2fd86bc258115e8e76f829560a7fb42c71b61a35455342fd5269e21f64a32;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ac769f380302fb7b8926b3d9669fa6f5aacd1575f772e10edfef8038fef44b8d0185b7bee52dfa4d76130011db03e9497ff8323d5964452cbf343c0bca28b1fe732781efa59d3ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1961faacfbd13f3ca48f2263a8a0683f7c849365a1f131277e783c41927f89edc149b5fa92ebb815bcac038d1d31b4594c3378545279ca7d5b7cd78e60092c4012eb8f7ddfc577;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c107380a1f04dd02bfc21857ef8dbd0ab14cb3c24f52a0b32020162335d4f6743b1cc3e7969ef87b2acf2edbf02b21e0df3dd7943eb75cbd53b8353efa0f8aebfdc0b53a2838756;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf27530462a5e4538b0cc01dc30efcbe50f2b1d3a09c084fc2456b2dfebba39a5e834661755cba6aee7aeff5ff0a4f9fa1e26ef9e861196fe2cd3efac898de827a84743e9dc6a6fd0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha318f228d304cbbc197f5aed0655bed32c54b135c302c5a6be461a43b749f43aadbfe92d4b8abd55ad9b61b9d172a19921f28860c2179be52d7f2f4f8701871e4f0c413db28decac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee2a6e127adecf905176f097dde4ac33aeb9cb39c946d7736f2fd20f7d1193d14cd12c097560e4fee358e651c35993afb3d0179bd1875bc1eb676c17bbdd6595b5b6b40e43082173;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54a27536f107b4e7613af276c29ccb0ee4edfb36bbe33d1514fd7ab3dd737f97a51085e2fa15000ce3f7e67e52611db54422bab32241432e74776d0631b7b05ea1da43a8987e696d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h496e1cf71b1771c7e1354c45bb8c2d07a5c3812c5fc3adabb0ab5afddea79a5dc83d226f6479dc3dfcc56ec20cb15838491ee5a64cdad8636ae1517468577144a3903831d97bfe5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89c48adb38003937127e806d97ce93c6a19cdbdd4403f6844a8724737e8c0ccc6dfc45ecba5d42d8c6e74e2a35c7336b5ee7ea5ffaea05fc95512157da2eee6fd5b55ee9f1c65ad7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c21f036bd157571db332ef15cac3f9bf5b26c08b64a9d20c89cdcf076d8cd4fc9f1983d80cfb6da3c86a29eae4b2bc9eafe3ce29dd2cc2ee05db982d35b054955c94b0c1e9a48a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15b03b125e28decfe86b4b462e4ca8aca01c591ab59028baa8771880250907ca775ffcb58261566cda924d1ce0b6490657378577ad56903a84fec5a5b4566ea3cc9e5e70fb76e54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8e4afb456de154c098b3630fb34a25708f39b9b53332d78221ce2b78e690ba5a856f0af06ecae206906b228df61834e54d440fa82a692ea64c79e97f280c2b8c6424552d85dd71f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c79b51cad5f0efb86a4de932bc897989f47dbb95cdac10f5e40ef4af39817698a82e46d448c9e60c5cf31effb83c65d0fedee150a087de11170842efad7d560cac78daef192048c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5ae9f0dd7e061f7b89d5138ab9607f8279781644c33cd02db7f9d14217b845e6d6d81daf18e14b48a53e0224ad74e7f19c211b2c6a707dd8c3767c2c846b5cfce3aff9192956917;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fe751ea0a278881c9b1f95ae8b5cfbfd7698f53f04c93dd6e8990d154a0d482e21f4e7a8250bb45e5e221eb350f88657636ac107a31587cc966622dedfe229c7237a4c4c35ee037;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde5917518c72aba02b6950295484ca6f19724f9546b015ef27b4300d251141ab44c1aea5d873a11479bfccad42703dc7736c5a66efe04fe18b94c3fa625a2f5196aa9544b1552505;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe9bdc520806a81621afbb9d490f60eb0767443543b03c664966039754613e38e6e1abe331808941556dbb2e94ed4b14f90bc9c017c078ad224e157397509bb1edd605524dc866f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a2a16e24d292aa6426e35e26d235043c05b6474f150fd0c252bde70a0c1044da14d64c22ee6a7d747b068672b6b2bb281ca5342e74431b429d6aef00a6dfbfae9f1825805933bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc43336df8e869ae1edb7804d43abf83f7a364e6650ecbdf0af3a67d07f9c8a121475523dce27a48c44ef4e4248436259764e3065eb6cd72ed8ad2b5b9d39231c18458a5057cba6f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h348aba23bd58157e7c58dfd3421095201f1dc256bf5be0e667103af33ebf53c20b1c198941e9779d2612769a98b948f0b44067b5ebf497f163d1f04bdcb3d6459839f1fffa50e0f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24e7d1de94338429ea0a532843f6accd1d20f45e0c4ed044aa8bbd9193ed21ced4e595853ccd9ce0177d537960d1175a66419fb368fc751abd1db2d9ef69447ab38bb037054b1395;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a86195722ce6a7e543431d46732486856c033efddc27062a57e5245f827a1e45a6968aaf3998d8ecb57d99d0e5cec5f5dca88fc1d963fb5b76d35601ae9d5b16e93358610e862e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c4c821b5aa6845ca867e8607c43d9df3215881eb1f7be0457a9bc4defaef83f1fb4aacb2c1c35b5b512832c906df9cec88c0b457ff210b161ecd38ff807039b0f6f387ccfb388fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e9deb647d67b57228d9201585f623f23794bdce314d2411ebe7599c17d3c61ecee8af9141d30ec5c8235e609451eeafd56a24576cf71bd50cd541b8c265e0b9f8f3130107e1cb1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12d35f6187ea15128e66a02ac6ab25a4d29ec609d998b2150205a98241bf93ce2141247cf689151f1ed1f21c9ae13ee10a73f1de134d70e5b2342f64ce09907a821fe30c47c64b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc871de65a61625a07339a7380928ae1715886c8aba576fedca4b16a6998ede465d36d4f8851be732f5d770e3e47e14cb938aef3fbefbd741facdce9d54877c4e2cab2fda0115be8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5df5814ee7c8b4e7435eeee476d0b16f57b72a38d898f6597f778702c5782a773071d6cbae29b8e14b11d88173c29ba0cb3b04d728032ebf82c088841f52ced80f7c042e5185ac92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf91572455d6fa45754437562211314e32ca8de24c98a799fb7fee3e9c469444addca12ace521e23f002a831f3513e062dc898ebf1d5e213b4ea5b60f411c769d8e4fa98d8abd48e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h506dd92bc234926f40d149063c761da3ba1ffc72c5689e422406fa79eede68e32afaf2ac64008934e241948ba16b43630bcc130c962fe81f0bb30973f7907a11eb2d6610fa751c91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b055248d867828cf6729fbb27981afdc99bfec0bb4017df4843d28a0e2d6e3ca832f066a4f51876759ec469ff232c267f43a4ea62df927d5f7830db0963336e144b79346d4e7bf2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98c3f4862fb14ca5d2bef93aa705e83f6e7fee715b740ffe25c2393adef35795a0940bf62494fc558f519cc7e4e5a93f4e7ac3a7d7e501bd3ce5c8f5076fba6bfa5519f23ddbb521;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d6a97eadf88dbe71541975172bd1e71f27fdc0542baa72310893777cc7c80a4f7d284aac9f8aa9dec80f08d17c7df33ba6364d19ed960f9cc9c7ba8c47c78a983a6732f6d9616c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99514e903277e9c8e1687d7d533a8d14cdae82053a7d591639e41fcc21631a2e86348b765b2aa4d231a38573fbaf74c469fb262ad22d67db3acba58683734882eedc317146e1e89d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67b47469fdfe5487072e1aa8ee26b3a8ef0f338d28d305a7419937d33db2ef39d6647f0f82bbd1d8e5b66f807010d0be5e2cf379931dae317b88d090be95b3bcb1241c95b0fe9f15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f4adda4179d25f05d568016b5069891f633bdbd1fd7fca6c07f6006c13489ad19a0b938dee57907556e19393994ef47113d44878c5a45d61b93d98fce1dcc627124be59e8ac5cb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7191ebea1e7d894718ee54b30cf9bf906b1f05decc1fd648e3441eb06e8003ffac592b864b68417a34005e9c895bab20f55c0b4c4831a20e04b6bde85c2ccf8092efc89716d16899;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed84fca7978a35a562f4db5cb3d71a7e4e4f3c98674ed18c6ceb052f9c24b72ab1b5c1f99313626e860f8fa9794aa92453a47bb2db3c5e92f6e2722522eff15f1a5d36d81d6a4ac1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f9c9da7bc1182bcddd4c9500b859413e2e41f41dd9207c0293a0720d5b5cea9d397d9344cb01d34477402c4fd5ff440a8bd0feb5b648c9cb809c9b7e463b3bbe8a85282ab78bc0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4741a42354748c2b8b7d7037d19a6d2726d3b4d6910550efd2ffa0350cfbda30fdb131ef0207172f19f022509a9ec3f50604e4da1c6ea81e06a2f2735b167adadbd9c9727d16fb38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69af575a0241a85ffb6b5f4308a76a9f5fd0248ddccba4745c26538c33d1fb0fca8436e2bd1efacd6953d8414bc610e1149b3c4401e120fdc011c80a84d32e59db6f82d7476afa7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51f983714057be52fab887b8d8c969cd295114a6e06326742b2102d6755e4d7e7628d6a9fcb95382d2151734deb6552ccbdd8e05c9d192f96f572fc1933bad9a3396431e1cbb7189;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f1a011cb928c9494f1196676ec18f9babc1422a605e4b3079ca7b53e3e914fb5488635b7f015e62de56376c88ec888e66dab7016fd591b3cb68d9745e5a0bdd3eca59caea5223ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4f6401ad0bab2410020dcff90684e74d862b187d3f87ff6cb0e51284b1a4fee7b4bb5b58f99dd40ebe59f7b99901e9f26e2dc47ad97134d26e0527111a2b2b03b2045ba5204cd6d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cc465d3033911353b78b7db3714335c73aefbdb2db4aeb4c635b364abdc72260d08ab65cd95fdfe8eca59c1093e8414f35c841fde619b18dad52e333a4bda8efbe4960b8af92f6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80ac0bded7f819b72b5326e1d20678d05d5ae38be6896ee732673a336ecd2c7d4e29c047b31da1932ff455c8a2dfc4f8ffa573d803841fd87892940f2cc38aada165781e26eadc13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h135a3fd2d850e066bee42791aded43fe9687dacdc79b546cc944412a032775c32f77354a305480e4c9ed96c59f57c7cd57d2dcd58635f60e47afdec26bf4aa90b9fdd6184a9eb0e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf889da307f178c58f2ca1ba83bd8ef29e85dd5edc26a118f362b5e04300aba805906065f09770d93a643fce653cc15eabeb2067c11ecdf6cd469257caea7f70f6e6b0bf1d6dedc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfadef2ec800ddadf0aa8e8b2c5af2b993561ba16c1eb4cbf586db56298f22b67102ab55b903e90aa7f722eddbb064da880cf591a533b515bb833c537c5fadc41616915888be6ed8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc11a8af57b397ceb4208832b9307c9d6ce1b6f64b4037fd5ea7fff90b4629ef79e2d9d9c1e5232d4f23f44af10cb4648a70060146bbeff83f8468352c469f734d5f414628889e9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e14724ee451f1ba097f1934bda00a06ed0e049a57c51da935056507ec42a59066db0ca681120a1d99b2eb82cad616bcdb8542b56258e9b71da8939decd2e88ba67b70f82e475e89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2eca89514664f8d0b88cd09d3d921a75c106ab8eef7b326e976cb4a73e455f5c1953b83087aa87a9220d962cd45b58a094b9d0d46e3889563ed19c43dde1bb1fc6eca0f3a0553f28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d5dd066636a667e359a52b9e8d1204c6c29ca57ca31be0e5a82f1aab28e07318de1435a5b26c7d7f6275b7c017eaa663ff213a0893f23770af38a79840fca8432a07aa8d54c78c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc69809d5796d1f7c3a4ec048d9c3eab7dbb6d4b6619f1b08a2067a5c8dfdbd03df71e8785d46096b144904ac70133f56e0747bc784428eaa9eccb28a008ab31b9e08963dbbf5ba4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h490dbe75d47cf1af21f0c9cc91e14a86c6cbf4dcd426d5f544a5b87f7bdf479eec68e5d5bbf2822126b4f1c176e7ba9da587dfc2420006b3cf3ed2809e0184b3b0ef78942d61d250;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6b491da39500845ab41a23c99524dc4ded27e2718b4dbfd9c6874cbf234e02b382e0e628c32ed70d7dc6a7166e87c4e3646d11f5e5b34488902b0c47f0b8f3d5e458b36e74f761e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d4b8b515304e864db7f8a438677bc19f39960d3bc0a7a5046df55859984badb14e701f09fbb4d7ad1b3ec07e96c85906c91f908bafb8a81eaa65f2fa4c6851b88048912125e9c4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h904067532f5d58270559de7eb0c9216372ef5207e5ee4a45f98f47211f671e142e5c6441c38367842c7ba038d3c225ecd62c6576e562527b9522ddec155fc22d2bf95ae9f7f3796c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b6e01781df908b60abb40f0f4d018a58f06e05030156858446fe908bde367032da7826796dd7112a68d80125a2051d6182046afd6674338f2ee1aa78f98d29ed3155221a3df5deb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ace26b6094992eb31ebb1ff8827af30ca9132d334e8a2220aab39ebb1527a0ede2b1157653d122d0a70dbdd46ac23a7a3612fb527a7ad26d199474a02bd7787cb1a14b4aed0e37b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d8e755820b36901ab45bee6ab447e1cad6919ba8f0cfbce57877fead681248ca442dc2a6adefb159b537d75afdda3206bde6068c0f72458ab9ca20f264f09d32105fe7ef486e1bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20a3134a6411dc59fe0581d2fe1e83c74389bd0f220de17164994988c01777e1ffa0d55a77fbfdbe07980c9a90e54524f1b7366dada9881a8eafe5bdcfc5fd11f461091138582734;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7372415f1810c56b53cdac6bba6e3ee7605baab2167fe9ce76964cb0d441c5ea3e712150f3e6fd979c9b031eaafedd23bc8622713e1eec079492353538fd2a888fd2111ffaa16ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48103516ece039679804cf75bf990d8f3321d415cba7df1fa63ce2ffed826902889d43b34dc81629435b65c5f27a1f7ece5df66997dd68cbf7a32767255b599536f6413c7a5dda96;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84b50e61ee704640be615574a49c0ab847f90a57824adf40de779656e319f0b9c0e53496d5225a5b47b82a006c4773e47ffb926ced0489fc803162824164b30a02a59ad7ce2b454;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h199c6415115124297a3ba15f2386e33632662f7af95bf48b9c0faddf052abbdb4b592f283f3180c8b00272e4bb4c2eaa2c197f48f9ca4c534771e528a72d46c9b94402b97be11784;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a9101f2d3da5a5bafd93c60129904265cb37685765ec50b2312284e41063101239653934d93f38886adace62859a3bfb75a91cb267e88838f60bf990f2101924c1e8ceec47150b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac907353cbc2ee01680d29f8c6e3bb02382e0f95c213744facf7e1514533604f1a7c6d066304be51bad04e24966c3757266535a3b97d388f4168613fd91b975ee38ebedc6e729e77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he510059a9cad526fa557bb29984db4b935c0957e915ab985a3fdad18ab7add2bc3473bbfc89d2296bb1dce407477196d2404b7b8b7adc7c2a12aca14671a486e30dfc8260abf2951;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9792f3dc646c043129b25b9cc516b53cb82833dc91e921e5f49fbba52103b9be6df4d80dad8dd1b95da169e75dba19566728e676d51694814825c64887bb8a7ba639548446565c34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fd8b57594fcc75c00178505d5105a2b9a3716664d6dfb6703b6e041c075fb0cde37208e7c157d610c75ffa50a00cae193dc225f0ef36f9a4d439f4b21c516ed3ad1adc69cbd4639;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7948997e43f5560952d06a6fd4b9f1e2e69ad6ccb924e036b1c8df8f82bf7d7cfc3575f7a8ffdf5e042ce18bc2489209d639543e068a8fbac3057b359d47047755bdd1aa6527124f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70e15ee30bed0423e8f4a1bd3dbbfdef3cda3b0358a0eda5c78fd7a4a3f2ff8f4ddcaa85269fe7fdf558a452e2415510914915493e1b9e6431057b776477660f1a739c3c325350f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a583e93c8ce3e72add3d75234b7a600d49fb03359e675cb97ff4aba3216c8bcec74bd97de1d7be030035cef6fc5e1442f4bc4f19954950a91c3fd118cb66a73aa71a719dbba9ea6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98d7a08773ac7d90fdc5f68b8cd866a2105c92a6656d49ca2d683e92ddef34d3b1ab913cbd8fd42a2586b7a1bf2ee4096b5ed37b1e45eeaab808cefe3c652d5f965c56e46b5ed2dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2824442d5a643bb290c1c59f89e0b192e3570c96e7e5d9742445accbd81c2ed7322a7881160c78187cbf474aee4c32a8367a1e2b21e705eb256709f57367af27b0ad0c3e7b904f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4edd3a1cd6640146c9099df2eeb4c64b498aa855cec0d789816383f44415f16d4baadcb0bbb28a90f4fade48eff3d8f152ebf5ca34b67bebae6031426aeb77978241f2e4d4647e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b7e6dea5578ba838cbba5adb5f24bd1d21c5b906985682d36190e53068c7a66ab2dbb252d77942733a73a137d48ec51f89eaf9f100637c019a7e4b8ef3c621a230346150e212d42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ec319468c0294f0da00a9c0127adf32b4941905541f6ff60faaf6119cf8d38093dde231818855f346dafb56cb42695eac9ff88377ee9a89138bb852f461345955941569947b18c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7a251e2c70533493e626281c368fbf61bec480425ec8fdea6dc2c9802a235d8c682da3904b585481495577deea6e272ffb187e81940eb263beb93892bc28ed1c77c20f2379a1c2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d7b6445ef9b2a256b1fc8946c8890c1b68410071fd4147181ae5d504bd64137b14c4ad85fb3a47ef3232786ecab6e355af436c9ced30708ea074c7e187031d18dccf4a230eae11e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23760def64b95139dbd5cf81cf496ff478f5696b6c63063729efbd0aaf29148b90f1efff03d423be34bf6e6355612eaacd40b1df689f299ed74212595aa0cc1fa748e29af489cc9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5f16a44be0917a85bbdc0815e1ee888c810d0b668deb7fc0a81182dd214c25c5e32748a2fa95cb86e787e8a4f3de36c9e907532384a2386ee532cb11ef20aa6f8458293640bbd56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5ee79095413a6b7eeedec215e83e2235f15bbf59e982f4c250e0e57727cb28525c1476b5184edbe93bd96028d5e01390bff33d5aa395b67c774b765ad27686fb051baeb66f1fc3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbee2dd23de41625ebaa19852fb9f4524f86bcb3f70007c1a46f08ebdceefd00f74f0a3066d5134a66c86ba13ca026d60fa3148c0656a55d6eae896e46dd5742051615e3c39287eba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b2451599e29ec8331dcc714bfb4e02916b786c8b395ef2c5d4fe218ab40c0923ddbb0cf9a17a7ea869db6d9885effe0638785a510282e4034069ccead393527846153c28b0b9603;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb753efb09ff388420e89ec89cd34e2ec51e7cf9526880643716492651d85c36e4c139916e07a88d352f06de017593d81490fb80dbd3bf2bc06eb05f55bad87b8c239902fa2b9120;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b719608694246ff5320e95f003cc1b31dbf0cda1aa22116fbdb15d3291ac3ea8a221dc69f7455df11390c9d95f456d8def7b1060c48c775bfa690363c5d9ea4e83c4bc95b8393c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h760915490637157aa035ba9b3037016943e5ba3881e624cba481a8eef1a47633bba8310bb085eb34094875d5e5d860b2b52d37e816637c4bfa7bfdaadb5c01c7004bf4a20cbae660;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38f0edcd72019a0c46e87c695453a6b04d6eaf4e27e1233e4842dcc32ad3597f443a1ff4a3fadff16d58128bd8ed5267a4186b57525a87ffea4c75b7adf2503c0d39537b976c10c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d34afd0b9304a532dba51022b0e703d723f1854c7a1285b7c477a97f61b9835df6662ecb250c96fc427be91948f853bd5fbc312dddc61269b2864f87aec6d41222538a449281c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5616ecd6c8e0af83d11788c38c32718b53340e976e182e8227a34c36574f550d05c93d39fedc08eda608bab919fa5d47c8f34e30a49295eaae683513b629be53939cbf5ea882f1cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25b4114c14cdb0e8f94565d94f20aca048aacdf62eff359430987d7a79fffffa856170aef0b9c60c850bb1fb3117e9e61837cefe62e3e2e36369ea20567cc6a1820b7fab6f21613d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf86e732a10d726e6b312a48b44511e1288e986ed812425117d6cd618598684edbbdc6da66c72f315db5d530f165ca8818a3c317192967ee27814b848139707b955d2a0aab51d69fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf64fe8898ca2fff6aacc4f015db86676c0d40bd4d5ebb389173e36f9f56494464ed012a197bb199d7a42656d4a2fb44708821d8dc70be8227db0291ecb7e158ad10edc1bbe093e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd08a9611777966161ac9c2b23b74ef205148c39400cf808b33266ff1e1b5dfa1f9b4df62c03d8a18c33a99fea1dc70179723791e53cb9aee3ba29414eae3ac860d62ae593e8f74e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1eb1bda117b17ec7d2ebd627e217340fabb6df6a7b0fde150e16c09435f81404afa9a7fa356d8b90f62afba41b94b802ab5ea7c80be73d6514644ccf3cd3b7af9087b2881491a51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86324742f3fd3e38ff953c8b905965f42501d55ad1569c991a04a6ccdf97f8e8d54b9a280924f280b1755401e56662f2c5fdaa02a3b21ad86475979f6e926cf73a2f117d2f9e6318;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7243912a7f0fbf56c2b013456a29dd20296a91d65c14adca4fb33f969a64d5f5e7a219de32d215486ec4191874e11b7ca295691a4b66f5460c7d8c71f50027985b212b73ad0c0d8a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h309d9f2636f61d13097855f331d5a3c50c3b9621409120ef78d4f1e8ae700e6e90d559dab67ff3c53f637cfd88fe3f4266dd892df8cecfb57db4e0d60af83e5664bab25fdfbbf2b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6cee8a8b8f1fbe777d0537cc38188a04046be254b8ee979c3e5b011beafa5d54879458a11612399dce569828f2db33c3e3093d8d051815a635b223e23f4862bc9421f8adc314134;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b368841ad5c106abe191223640021bd2e820436443116cbff219821d66695df875e3e11587feb8b45056187323bdb8b76fbeede15dde333697706571cb93b04e6de2a80fd52648f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9922ab529a0b9d08a49c440ea3756d15ea4d0a817fa2cd0d7b90bd10b05ea42b823ffa47ea93c59a7325d61428949267cb6e346cb31754921011423e4c6a1e4cb0867dfa7e26cbcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50962fe711da722df651449e1e209a3f21d01d04a60b6e303dd7e6cae287d6bd07eea50c50fd29ff9353347bb9a68bc046454327372be26d1ec8e2a1067257724d46e179ded1670a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h545b6bd1f63cbc1ef9e909293d4ffd7de9a6600b01d16b2afadd970cd88d36d91d6f387c8c2c1c76a70e5e9b7147bbea6db666e64278d1ce7f3e3ab78c67d35e5c3cae46706f1297;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbba0c8741fe42b64ba83a2406613e2eb267059f599f244c718eb79e5a7eba75303ecfd4fa1a0ee0f7f58aa78feaac530a8548b8defd3762edeb4d02915b3e8e08f4c89bbefc9777d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc01f465ec17da09976d48eb1c57d63e4c4c23aa5ca208db46790b3309527b9ffed9c1d2336fd0426d24542af312901981b62e94bccc179eee07638c6f5edbe5464ce1fbd34f3624e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h330802052982832885c243f441cdc673366b9b4c7e4275844ef49f1b945015e71c4e1d4bd308a841167142c55ef7f8f8b7aeb0c15cea86f3da97e20f2a7d1fe7f30d23a663199538;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9c0b0cdc4913ceabef51a1aaed597a55e7dbf523780c5fd45a782e9c6795a28720890d37137da9dc3952e08b421945e4412cd9adef501060d535d6f1842b6f1f825f5a549107525;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha54c1b79a3c5a36528c5ea60d240d2d8035bda8fdb555627aad08db668fb7fc90ef899606ca1974c04d83f20f7e84a28dc7efab5cb6ab560ae95951ee3506de58f9e8f87230e45fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2f97a99ef90fa2bfe45958fa2794584c457a9838eda7c6cf4ae3ecaf3df23b50bd4eda247c1234317b1ad04f9e1536c48472d8de2a9c00ea41e4f95aa3e9cd392ac1c99018503a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a11629e50669618f1d79282cbaf978d88c7d804e342f4739d9ee26cc4bf79ada24c07f9f1f9ba0a0a790ad5d51b81b5ef7ee13791e5f10c821b0a2e8b8f3b536afe646042c9c067;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82a5e9aeb10ac309df6b0e1999019595c0bbb1ecd2277b65ab7ebfb6c1a39a7d6e815ecc6a1c7d2a59c667a823c4f2add549ae155e74c9d6ae6d6c9778b98a36e9362c7a832d1e0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc561152eadbf21962a008ed8ef23f71dd8a2a1ae17850e1046f01f342b56ee744658e8352130974ca1f6a57a0285f856d1a36ed640d074765ed4556feeed8dada54d793084cd0d76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb333ff2e484302c4974096745266f57c9321ee94ab3d1d0182a825075aa741330c4d5bcef2e9a509435993d4fc0bb372741af79e26d9424ad71f633ae9d60b00abc6309db8c29446;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b5c6f0a7c6ba22068f1363f3e55ed2542deca777a400d4357e919667750a87c2e3204fc53f5ba977d88d78cbbc59a3745d7678efc9b90ed69ccc7c52f30583192220d7725ad82de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6d7908db6eb4ed2388f3c55b849d2b6afb45f38110922974da736a9caedf3e6887aa3292c0b46fd4d9b64c4d006e7d8d0bc4624dabfd173a8fdcd4fdb1f1cc9780e7015ca07bd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha249b0a6a8768809b5b23e251af667e2ce84c77d2769d80ace4bf4d550ee69b6dc5dffe46e0685be96600926fcf65efe5772a16dbd541663f15c77f1656c355db13da7eedc9890a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c3c1933041fac5b735d8ab150795c04a0d06f165c3c21eb43097fdaff619483591521c527b017d93080e6c2d309e9faa10d6d90a879bb183a61d51ca2fd0dc674fbd19806e61f7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57c71b7319c1f370d639432df3fe1e8ddcb473ef464f4dac72b2cbc237ae308d652e9b82fbe8b3e7fb2c8fcf60a36d09b5ddc9878251a8106111ede116b39cce91ffd68a5da31c16;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7f79334dc7917658296c0e7a9b3c8a9319aadd2d78bad8982ffd74b4030c8d67f2578994d2ef0f8060c279c759db727b8284c0fa77048cb320f3c1f3c8f576ddaaa0467299c315e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5de416d4bc17d0034d50708fcaeca23899e3473bde2ed5554825cd37265a869f82617a2ba12efe9e7c2f69e48265b558fc02a53e949c9b3cec02647477237713b97a5b6f9c5a7010;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d6fbea503d5858bb969e507b1b51156a279ea18aa8d059984169fce6d9b68cee609ccc107595e7c32adb6cda273e086d5f853722d94a2cf2b604fa0dc7a6c171e355d737878c38d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc437d2621cc9bc1df3b03aa9b80feacdb2419405ab3109ef8c9ced3fdfb44ba5329ef9851b9ace413322c2c8a5c40244ca0a8466bb879896e573f541cc261cd69d5747a190b24875;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfad318e2ccad04aa65b1e4f710e28423fc40df6c0785a1db5894f96f934bf1894624af9c39a7178d7e091a22025a0ad8a152394b5a6e3e2d9732f4cfc0b22cff132238aee224b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e5d44178fdb65d801ff52e7541a5cbc06dcbfc16d3ffaacf3f11466def58a08e5025e26696578e9d03201dd9b56f9182d759b06a9a16b76250b38f45fa02c375f84bd2fda576c5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ba1042ed7616092663286c6456616e0a70294892049a5f663c0e11be7c0eaee25d2f20ec8c7592809dcbc81ba92148a47424c9a0d4457d47418c07c3d80db65daeb594a2b96d85d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e201c05cc785807e5dbc82ce941dfeea5717f13eaaa4b11667d95bad67babfacf48b8d9e353b871e43a3aa18c8f3e040536061ea3085a3ab9613dffc42589d997e530fb36318104;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f988b29b3313db59ca55a01f4c620b151d90626837270b8ba631cc931472162fe398c05817df4c866d996d3fd02968e9b77643eeb11e02a495e4038bbed820500204554872581aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed6d5fdb08cfc0f6283f7ba8833fdfe19f8a227412b786fd088edfd223ed18b9eaf1e393ae15f6daffd4c9868aed2b94a3af5420b2d9eaf52ad02f588df163696c63c344712bf6fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbea3fd723104d30452a9e7403033f15847c79e01bfaa53812a1e129842814f299c050cb007a9bcc85e1a9ded6180b21c217b7aa0db66e120865ca1f552196890ad0d98079e2d37c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7b98d23012323fcc9aefc36c68b4362ebefe8fe555aaf18415f11eb6b73fe10a1f10c8d7a51e1aaf90593f2d47657d79d1a68e7c6979e6a95698e4a86d025c73c38fc66ae70839d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e840fc84592ad31edacc711e22b7cb4197aa6347082c0f0cb855b2fb564eb94bad1258087c9da37b0b9f95623381bf31037c06f38ff8b2331228442467b87858bb244cc0602613a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6703e33b464793a6398b29033b7608c066dce925993fc4e38bf374f9152df7c068f081dae3eac39bd6368e305d3ed342d1945a444ca5c964fb864c98cf74b64a9b281a356c4c05a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58be05a094191abd63e0345b40592cf83fb8f95ad0ca17728ee6b6b63d474503e5882e8c2c5c26efba5c52a5ad85f0bf79873b7673653b3f9cf0e8c2cef4d13a47886c6c8f560a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he987af2f8a48c36d9d463d56263bf5224c577d3b570a958f94cf16df7845f118b2358997d5ea0e91d429979a7461a0a9fd02187fe1efb52d5996917c97e59c75316dd251b2303bbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce95e5e4bc851916c44ea518cce58cd7387f08389b4fba97381098079c1ecf9380843bccd5df596754e7ea48ef2494f089c502de1915f2681d4e896476576ba7b7ccd67698113426;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0942b28fccb0a92b253bfdd068b44cb29bb2f2b6967e0b9d6dee9bf06f0c22adbd0363bb6bf1b2c1349ffbeb9d6c2d7ac52fab472734cddbc3ff1d4efaf4c7497162baf2a01e51f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1cbac4cdbffc4223b9ffd0c1366bfbeffa46151b58298fec3411ab674f2ff3c9b1a30c6f307957474c029694810fc26811f9f18b7f5f6036735749ec444d1d2b4fe92be1549377c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f21d587e43bb3627170f17e677cb83674a1ce144989b8a0135a6990e50c5db801686b27797c7cdd1300c8c3bffe0ef1e3146d17ada6b1f2342aa422f103e578051161e47ea86399;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ad882d16952eae7abd3a9be1dabd7f467234076ca039253b08093f53abd6b802b9845aa96bcc2bf25d7d9896c04b720bcae40694786302290ef1cb447bba463eaa40fd75121e663;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0c1b86b28882ce880b070729914176e32fe078b52cbc0c74bd5eb06863d5d6549f2d6f8e61dc53ae50a2d850934a53f637a89187c720eb6f7ae38edf1386ef57e9c2a94be54072d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbd096d611936cfc30d6adbcaa84a3abcf32ba393cff9389398a9748a204a4b75bda7cc1fd0b3b128dfbbf529b97b2fed8d6c53d9574bbab53c88e3ed05ab4916d0e7b1e727e65f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4be9b40c17ee828dd0f520a4ea8abe4e40edbbb0a246848915c78108d1ab910c0bca8399f3fb613d757c29c43083c07eece7afd628d7940440eb8d3f2af384013e0342aaab4f43f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61c9f00e1424bce89e46904506ad12830ed83190840476b8660fca251ebff5b6b8fdd02319c1191024ee51a2279e13d694bff42deea37221aa5af81a90b66a5666db62ae2f2ebb5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h185e6edefc8fbbdef018eb375052e3b4f43d7fd1824a5c47b5ed7cbb3073d097bf12f8e92967903d44f211dd57fe88eb8388dcdd12c3f09d3f0069fa1a5506042d09c523f9a8d8f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e7e7f8221de98e59db9dcad67385cf4e5809fe38f642438eceb40f059aaf75ff8a585096e5622f1e6ce226539a3d63e18d487cd35c9b32b92fb842db9abc3c799cfbdbaefd3d4a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba561c7a7f179f3104262a90e7095e472c40f44ea0d776007303707d9c5c6be72b92157e480c157302c45a32c0eab28df1ae8b27eef700d9ecdedec5599cd3b3345afbb30314d777;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h963cae08bc0528f82b38f4b76ed8fe53bbd48141dbab44b8c57c984a4b5e6f1611278c6c92c347ff56b5bb2ccf37544682dd21b91b17ee218bb4130cf1018752b674708e72088a6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64a87518a721ce0df76539494282034a829e201548efbdfc818242996b276bf913aecdce5801826fdccd2b422740532e1cf96662b694a6d3c395a03c7abd6edb609a06518e101218;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf89ed24591e9a0b95962681fb54ed0086eb037d220b98cb742f3d4a7bde27c4d0a58beae13a53e1097b8ce75b22d06d002386e27c3b8091cdf6a3a07fa92cf5df6199b2ab8b8f4cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ddd6d392a628ab1e94babbf8d7295c496f204221ac48e6684e649d97422e8ed1db33205dff0e931c0d9bc3cb2ac22cf3def7dc49eb50cd3f6522817c439d87ea306a345b91aad9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66cb8d6856ba7ea03a3683115fefcd7ea27da449f862ba0283516b52a7c4a7ffa7bc568cc86f9be885e692c59cd445e39275f4be1d01d257d79a7cc6984ce237f6107d3c0b72bb4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h908ce0f6c3a3e74c4e87ec6fb5c4192cf5d9b5d81f5d3e1c3cf7c757eb1a04365e3cc1b538f783792b4d62c4485a5679f86ffb7c7d9fe3172eae5e7c82d457cec638cb7c8a46cd81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71d33a0ffa6bc4b1f13752b28f13a768cc724e29000799664ce75f09b1220030b109be38b4f5bf99187157837bfc54248a5783d78cce1260a683099bc58c0ef336a2930965b0d0ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71d282427381a25be3e05ef4f8b57d61dcd5134cc4be8a43a8771f084b18f750c48ff8fe06d500c989897381bf61ee97c053fd51d0928ae60fae8f27cfec7e557219a8185139eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c34a08eba5234f8f057735e03b737f6c472cfbd42bf43478add743c97f07daaef20f460f5266900afb15aff8b057ff8086bb7539a6522880f4f1bbd8ec2611a45e78682b6d0be5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe120583b9b01b88fe4fda781be79d2ab33469d06869fdc505822c6a302dffa9ed1d500daa7f0d2194e7b69f58b6cd3fbb517e9909a27c5013c21b744d94656140b1b601b4fa8c17;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7235c28fe588d7a9673ce43e4db8576f24c74b852368de0249550d5ef9da98a439f16a2e6cfa6d2e55ef5b996d040024c3a240178c87b2ed3cd0ffc85c0afb86954ef9792d8f2096;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9f4ae8da1194c891d553c28a01b84bc9a7349fcd7324987f0c2a3ec656b9917ac913cf04588f5c8eb14cd33de42ea54f785367623e1d15feb473636a61e8ca732302ea1d59b948c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd14902a22692b2a92aaa9f09bd31bf79c840e14b63944f573e533428dbf01fd569ae2bf0e2f336b22a64d1d8ee65e67501dbf26398bbb6a03107f66fc1199d74a03fa959e8c7f258;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h704c147a9842785ee55ebd688151c2f6ca7b3df8d4a223f4f723ecd1fe5bb2794ff93f0daedd3b36600191627a7d4beac990e1b73de1782a9beeed883b94341b4b41ec53ed26f84e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd84339eeccfe89b7455e2598e91e646570ebc6cb7e52e8c0e262d8dfb7678ce6c94ee7fccfcc9ee71543bc5887d75e24887d252d4a4707fb275b1769efe6bcc18e1dfb2284f82a5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h592b5da00780191c79128327951ad11c8002794556e7f6e5b99a740f8ec0a0f9d58d59358ea2e858837f6ef5acf6eacc9ecfafde9819df630cb3545d657e3f5a04b3858fda226cef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h531e68ed58653ca308e0588e8c97c06514c8cdc2d66a65621a6c44b42862ef8790137be3c72eda994d4466ae4ef8724e3edea2e17d5b3d5e3320eb2cedc0af94c0e179ea6f189d33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd68dd32ee39c8b2b4e1f5ae7b0ad8f7415d1c97f4ec0ad95802e0a5196ebc60243d40656a6cf3c4ed731707b30b70ba137dcc35fafffcd7b4cdc7374e6f1fd580d562582bd40ac26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9279bdd444008b30355fa2514119d6048002b58871bc4492d422adb3f9d4c002fe738aeda13dc8997f54f3e1843a8b14011732ad6d485f239a9715753202dc04ae4a8a1fdbafff19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf411e0efd5cfedb23d83f4bcf27211ea842bd0d5fda3e50539a986c80ceddd63804607bda1b648b1e9213d44f3c35a8dd2379ee15716f2a5499d3f4bc7db1ee461baca3e7faeab27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h737e10a109197a49734337bc9e883cd1fb6d0a49d99ea0925ae4090ca0b2d58d789380c25120eb85eca1b68d3591937cf766818fafc69a63603c75ec0b1ad25edbd6ab3813b0b1fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb7562920cacaaac9fa784722e105f183831b33ca17ddae92b71f41ea8e0dc1b4348f3b31e3c5e7e2e25019f0748c88e8f0752b5c3d1d592d207912c8ddac3a359067bf999043b63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60e5fba4f2fc845032a37aa5ca69729a6c415b7bbca21740fa08309ec9222d25615c3e94adb01f9d2e3433ac00aee14b899616b7dc6b69591d6a3789dcdb1e9aaa98dac6886b80e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d35682a5c6bb4156cab09c0a3b366c64374479a7c4631bb35a10f6ae3193e452bb76a26517bf34f93d814f6e1abfcc75a775abebb2c300cfbe6680ca80ecdc0e0a6d583e4adb02b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bf4ea0e74a9b7a6e2a4be02cb89da660b683c3fc8bbbef0326e7bb28343080a02e7186721946af654ed5ee42c76fa1de72871ef45b4f62c387744abaf0cc6c117e92a02a5cf229f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8964cab1d8d034500e180c66b0267dceed168838d4867bf4bbbf7a39917b5502839a811b49f6465855b22b11e41b1dae8ee901c8181347b4246a8f4d7b78e936a95ea7bd40d85bf1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha38c45154fa3fa558ae377539e26392d59b123601503e7ee28bba0a018bcca8fe08c83548a21b41a4aabceafaf9ba20805f9279ccd7e699783a83ff43120ec547968085e456c4b08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fd119689be8c79b6c931e170fcfa0734f7f3264f564bb2770897d2614a7cd95e7744826362bcc007c47dad0d090de6815a2e89035105b53634ce3f9fea526b8ad36de6a1d9bf604;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd86a46773c66a87fc97479326c12cf8192b302428296bef2fa18e284df9fcc089783f0b0297857188d0b2f875c2bf0d0112b182b7805b0b88a410d2d98ba8ffe72343f8f6ee7cc81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha58614c1b7a8b57c7ad1b6d183aabd83605f98c5daae722d1e2ec62d21012fc080882a9d8050f60f1fd7e4fbda112d335917340e3344cbbe3b7a364c3964d3150a7b75a4ac0cf76c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcca19cf83b7a83e147388810b31f2cccf41014e8a1978a53d51421055e062683cf4b3519596b6e66102d2d807ca6b810d97858ef7dbcabe483edb740684dcf2998e90c149e2f9049;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcdbb52ee791b06be83c1f9a0d7e934239d4e510c086c55493e8a29f75187c7f3d264f5603e0e3af0dde693cf1c3d72aa8ee04fa9284261b206f9dcbd9cc96710af9fc1bb329d033;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d9028a603cf9815e58e4f66f88d438c0b23eb9aba864520dbdb1a4d139b36f7ee5d2079c38ec2385e7ad518feada6362b9892467bcdd457baabf8c48f40379ae646021807b5d0c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b7ff475c076f4b54bd7e5c9d13fb66c102a05b38d9a23246ce1f8392886a4d9dfb5c1044f94e01c95361e5b0703d5284ce468808bf93792e049962bac44b65de390e8cf13da116e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd009eaecd4b903abfa4bd5c2aa2c57298d0513421b7c83bc586a379db20ce984276f37927f80ccfcb9b4e097347cd440e12ee715e89f13702c3d457f299cad18192447a4b7aa6a08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e94d6b3a56e571960070cdbbf9a72a0858d6b88ff3a9af02a05c1ef8807655580a29beda2c3ad8059c3f72547834d9d19902664e2f332d62826666c14ff55e0ff57a818691084f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16cca4d270da20d6389e77e95ec2b69bc41df97179e6c32fb9903f100d53c8d172e630e860209a4898687ac434266f17d2b9a096a4a600606519bda7e872776a8cda054c58f4407b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f818f26f3b7c222dc671dc951ccc5c601ed87c44472205e046edb992ee093cd34e2e7fab6acd181c51db1d6f3f46252fe53f5335b8f16dd2763f4b568a9fd9e7ddae92c232c72f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89b9383f9116b3c751af6eec690be1046469071c8b9bb70e2dde9d3692153425e580681594cb37ac0dd46558152ca9efca8e40b363a073f37c64716f90250ef4c2e8d9cb5f38d99d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58a4a5014db8cd58e20f02cc98dd95cd9bab09ad0dec3e6dd1fd976a46a114ea638fb58e767fea1f03ae4b548d3af06b32625241ca963a21683e7d9ada36349adbd1d51bf30082fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba403b595775ab031710de3d64d64130a414f829019c87e14c5b2e43cd773d8a1ed6bf31fc2d73cc984575f174f83cae29ae4b4285c7e6b791b432cf3c018c332acf4db8e4ffd9a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee1aad4ae1b98fd7515c13ccc16af3ff8f6a1f5bbbb821b24375faec77bea3c8f56fe2faa0e64281a1577a22d5c9a2d10ad28821996400613dfb3144ddc973a7fb5795aa6637c4e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61d8453e0955bd619a314ba520f543578cdff0074081334b9f727a5e9d7097413f72a5af423528dcd989ddf9c7ee02467c270c386bf6e15eb66930ac532fe9abd96e30e75ceac5d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f3c4713dc6354e22ca081c485767b3bc5fd533ae5aa4a936360620f2ea9046aa877b45ac8682b370113afba3cddfa02c1ef0272a1edd755c88ec232247719b94a36f86b10bf24dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d8d7d2ec1eed8df8e9eefd582b534274917aa5144c1262b949eb26142101f618f119b0daab4fbce313f8d9e45abcc0d4ee49610661235b27f948d28eabba369066ad5ec6c15d76c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bc9e1af7a75c08883b2a7df264d8721cd518c75ccfbc6b451a3d4cb2dbd56f7c8c1c16328fbbafbd4fa4c6ef02a6a0584bfab2afa181261ebf7b2fb00aab9cba818a8176cd990da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dd3d1f330e0284c907c81b658e77df6adc735be47e712a96e9c7ea1a71350c015a6a99b9f40d6cc142133f2175c4483b06bfd51d72b7bd426ad6aa1d206e02f473df02b49d674b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd838176a9be1a3494d6ce400c7743415ca730e84ccfab0d3f41b06e7549671b0618c5016c01e5de08d65ee4a4b771f08c15bdaf53802c87899c956c4a5a0da1f6240b5dfd8c5ae50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd44bce24747d7dc102a480654f3da25c542475445ebfd538a2731eafe6bda612fb8ded32a8492928456461c1e59c3311c313e18b2ef0303710872355958bf1cd2e4b745f59c9e788;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb866161223baa5943f5453485c50c212716274bcd092f5ad2b2b0a7c228f0e26a8e35b4df8753fb2021aba0000e7bfd8fec209defb814fcba6eba8995a36e66715b8a70d3f765cbe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h695627820a4d71464d1c4f98e3ebe079cf16fe2675fd0817e42d009b1411df23b39d803acb2ddbba7c672aa74077960293c6a0a4b368d4b5396b8c462d1945d3960fe8bfe3595d15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35210c2e9bb5b7c89795b81dc46d3c42456921b5ae3c1545e727d64004576c79421e2dfe49b12acfeb0920e1e8ff09bec8517c3ac7ccaff793fe306ba0180eb074c0cf1ecede3fe2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf36ef59dad659617dae580003c2180ba4e69d824e8a3501fa7b60fd27b19c3267a328c237ac04813899ba81385a28b26b687341dc1610bc2c0dad38d97777b2c390d78411ff59a79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ac3722d55b8ca667ff903a6334392c93e49488b73b3ff1ac6de7e7bb8a244c01e3be2c475afdc1580980d62aed2fba3fb784ad0f70d87b3c44a5978eef4fcdd924cf12a72c3373;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb01a2040f266a5f1e9b089caaca090e33ea0b290dfb2b3215f74b52515e0362f545e019b21609edb670b6c9440d1f0c46fee2082fe9ec26206b7144e2963a574a3f9133613ad0464;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bf5333e08707e54326ae2b81acc20fc62ca28be10ca56e5e8e8c3aa00b3640904e84f8b6e6485afadd804f5b00ac22bc68cc3061152e1905c9a5629069fd8b99b803dff6821472;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89637cd8db4b8e5119e2cf111ce9352b1da64319d0b36f8f4ca5a59fc117f6a53a91ca4f91e36ac18023bbbab7bcf944d4b8aff079a86cf95972e9dff8063fe279792662c549c300;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d94cebcb1ebf311b7275675ff0763bfccc71c2ca320c036802be96a82df377c3423065a33918b3d8134427e1e4d62cddee1b3ca008d2406627c95ace65795dfec5cd18f84c4583;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63984b77c4a3d4925148eac11d1f21062c00a62d8210d4a62e8b1aedebb881bc16ad3ac06160cf02661dd54dcc225ded280f9f8f53bb218b44f68cb035d011a1cc0271198229704b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29489c843e89e858f8939b206925691cac86fd409a508a6669f55ba6eb8253a457e7dd3591da00972b25ff4ff095c1d1329c48965e8fad6d08da0fd56fab16d482cbea96b2ad1cde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd6dd79ce928dd76c704f5e8c2395996966ac42af8619988244c4b0a084734389c7a89af1714fc30e37228abf79a7091c3375b0284f05ea9962e1743ec892382af3eb1e93ca6573d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99bbb22c41b70f28b3ce11e76edf44e87c5b8130c3554cb9587fd0cfcb8cb1a115173ec60283c904eb03d8a9c68369f495d620cd70389e72dddeb1bb0a7934be52f87163ccf5607d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbaa4e4dc603c88cbfa9435429553c7192728fcf926eb8f52139fc4456af9cb191c01c8bd050f8245214108879aa026cbd9aa3489a533ae8d34f30365a24fcf6817cbe794edd3df2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bf32754abb556ef50327a3905f3682851a759220bfc0663d3593bbff43d5b4d2a1c0ac59f0a00cea1ed41898bf1ead7572508bbcb2a1df53e7bad3973f2eeb456878c3af399d302;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dd57e020bad937245d8f82ef5ed35b32b1f044c47a7ae4b7c290effca7e0120b9ce5d16ebff4ea4b744c587e5567c460e8fd682bb017c5c0366df1ea503a049fa1f4a2f80f92044;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he067399aa7ed743ebfedeb6c72ffa6da23dcd2e3e27c963ad1cba38c5bfea753a9edb98187ef9e700972a7bfca7c6f18af1d584cb43dbaf451b7facbb116964318099797a9c22dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d6d84479e57514b6624220b4de5a504b5de8dd82b82b8ced9aa3858856c0e848ab5fb660918a7688b691d11d7ed33fdc82ed1878664a87eda586b5b57bd57ec7134e4dadefaaf5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda5c5e48bb1d917c7773aed0ecf562d76ec82e3e0acc472adc6bfe96cc7433dc28576696a410a959050ab0fafa1aaec58ae869339317fa763033da638f5d8cfc66ec5ddc3e3f97f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dad46b3ed02554d9b79d3d3c6e514fb65549310ece79e30b49ea70b41f3d7093a6423094bc010cb9bf9d7e6716a2ca396f567961512fb38e5bce89b4f217d091ea6092176fac434;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc010e8ef9eeefb43ddecf9f918ae1a5925e1d10fa8e814e0a839bd1fc9a03d4db1d8c8226553386ad927d0f97c9e4c2c72e298b202c514a76bd46e2acf8c47edbe7f7e45a0e3d06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha308610766cbe7394e971cf1f6c0011d45556e87ca1759ea276937d5d0673d99338a7d986065c43d05501b84aac1989b47e2b262788cd218720f902ee5f9420830b801fd92495a14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87cc6a3d98b31eb189212e1dd9dee43dbd3c400167aacdde5b561607b81507929a2e5daac8d9c4186d86dc822ed9dbcb577471274f0bb19674b2311af9186f4235c6e1e5c2f18629;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h122096be68ac2c6cb3a2f33a219efa0f85a4ba696a593bae7cdabfb506e61059039dc7f31e0f38264bbeffcebbaff3385084af24e68fece29647140904571b0233a3177683a79e65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38c0eebb80beb7dd54760a2d3850ad0088689b1a97c72ad4f1c7ad2249022ec2acbe1bbaea9866749f9b95fed43ae456b33547da6477fe4f9e724b1b79a01a88e42e0bf23a6a4112;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99cc4e4329c2e3a01d9bdc14aaca0ce2f12364bbba1dcd030ac9cfc42091256a23321b75d2f8b8d915543dd7f0b7a980f02f87d7ef276eff0987655a1899396f3522be136208767;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e91fbfbd74db4ba022bc0838f0dfb93e048baab224e0d5da33829d7bc4832e958c4bb69c38db2d6030ec7988173beb08b3be65e4164cec67d15bb3aac3a7ae88c6e34a165ad9a84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2489d704f31bcd4d30ca65ddc5622c49ebd10c9dcd0e31bf3254132ceb9517fe5cca10f81a78771532169414be2c1d17cc5a2a756d3873392e7a1647baf7e2d3ee43267a240e70f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha577991627deac20c01fbebf6c5c0adb21305969f05708d379ed0e9dd0e17c1ea85c1c416efa18552066f813697ddcefc6cd64ed64b950d004c81bec693a6d98fbf03b05816b1b32;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he86db3771b40c3ff1aa528dbf14aeab68d3c8a8ee4c128d615ad09dfd3a29cd749bf310ec915cf44295f88b0365648f70051a187cf0ef446a6d2330509c923b66e845a9d842ddbbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74c59150f4fd79f01a4be2db7540367197dded3118c2b823e58c7a3ccadc3f7ef8825f0620558fbf52d5c33b0ce5b75dde4f82065dfb0c32b62567b21b8f43b8cd2a8a0196086fc2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9af15ad9a11ad16f6b4e0ea721f5b02f5644b65256ba15a5d933a08841ae841ad9d4289741db5c3fd1668984a00bcaba0eb8be8d71a6950ea4d27724d55f00905d97c05b83f95f8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h603f8a122501bb5476239412a4649f60f7c1602782df6903a93409d1bfbe1751224550f38fc9f7e339936805342621823a586824764376dff3fb9cc5dd0b944630e092b91eaa1979;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9950c591f23af3fcb06394ad2f8938d7b49897dbbc4785e08bd3f5489d82a445b930ac3fd521969383cea34a385297c574718ca605e6aa3f398b073319e64c16cae9c559b9c488af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcffd928731f8abe86519c740d2aad78b1a115d44797fcc9726591ce9d4a945d31c1bede129751d8605b9770172d50d0c0e7cc266d7390c5fbc78d57ca7775cc686eb222aeb6c727d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71d8822838ce44b402e93480d18c8a04f29690f29cc89631f973ecc8bbf7df077af34ea47d3aa1249f1e6ebba218ce58406d35b3bc395a5e272f0133e5ff3545ebf1d69155685b68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1fef1ca2dfa10a4ef5d9843af86c2fa02a9e24094bf1066d5194b7ac13ca78ee6a8986777ddc020574304061159234f41678d744dbef294c4a2d83eed653d8fbefa34d1b3741e07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11b021e46adb6852d3a491d30d3af0809afd07a273f6f4337e515f0cf500aeaad39ba36d338e05951e14963819a0e2bd6911face0b7ccd0994231899b1a7b95c6e24b532d59274b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b71e40f84babe21784c59cd74cc07b1213c11b69b8544e04977a0ce4948e34df0f66dcf105f691cca6ba8f1ee655bb7864ff78742dda1022d3c5ae1007c626c1109fe8e6f56fee0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5a76098aa2adab5bf2ef23f971e8d143e71e4451e9aab1d58d227036376d809898c006df3f30c4b705226904b9a0fa5f1c9022280cd9c5419b9c4ed3e0dd7a7d0d4f78fec407b84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc0eac6f40ab349c18c3206d933377701fdbfb4d466d4c1fb4acffe8ec22bb66c9d2dfea897150a005214a0a4cd8f4e9512730cf68a7b9f44e542267397a426e831aafdc0bd49f3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habb66b422e7512a3521e158aa768eb2fcc6aa973082742301ea7eede1f6fe66c1e3bab778ea8a04d17cd0b61f0a557accba53855758e544b0dafb08774686c333475c84e87ed9176;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf127f25217a164b8bb60ab589bcc8bb0196258795072b3ae71fa883a441c1967726a0f7bf2691f4ce6860cf1e2157ab66504c6091a9b5fc3026b5be520f709bca02bcaeb4d492ea0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbeb1b125dde4121a0554261cdf6d266fa6b5328982312cc0717170fc27bfec849e7862681b38a52c522346a0e38ce19a342aeaffa868a218f23349f45b2e456e79365da47a1368f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4bb3e0e3324183e6dc824d781e7d513faa8dc8cbc3411d6c969de3587d7e656215776b00ea6d08c9b52b1df55931cc0baf2c75003c0c876dfda062ea54e4ce7b854c466181d3de6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50f51171308d1a4894b24cf8419744bb789d90a51acfb8846bc75334d7630bc618690af7793a651f536857ad26ae865961b13497076368f7e543a61e1518c8e87f70387290b582b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7c75484c4f9977edfce50484cad1be24e4573a1d63c53d87804e0ffaa420660b6d36285af4ccdb118232ee78d394f78f418e33863e14f1af0673fcd39be09fda9c9e50852610b72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9fd3da1204580183b76182ce4121104cb6b8d94e628c2438738005755ed662b705ef188731176add148e530b11888eca39755c1f865f2e402b46c14f89d532523a9bad2fe59b73a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc400d96f9f099d8a184f2cf884b2b27963dd875b67d272fd195c4862ef4ee128fc1d97a9ce067121130d0c821ada4f8cdc4f9691b1a7b30a40361ef9d3b8c7a82352357bf18000b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd6c0cdd428700cc8ca366950974c04d895078cc45775eae4763189383db422595115ef204a2788366e3a0b36b35a5979cc09489433fc52b5b6b2f7ce90df746fc4e8ef2ffd92a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h340e82a4669d46f67a6adf93328e23073693301c6988f76f6c76fee0e33359328dd935eb11d413d957cd6c626f228ef00c46d51045e3356e84097a4c214efe5509a004af61584690;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae59e3e440d79b664ba952d9587efced7a3f83189674ee9c0562240b79af5b4a7c9d7d4a6ea3328d57362888d565ff8dfefa146fdc392d766981a94c658c5a1fdef736e91af2f530;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hada7c4cd1cab92d5fb2bd7eb29d4d60ba98969ed48921dd4508cda1c75edb972134235d34c6aa36013a78820c5dfc06efd8304a1a4da8dee21548bf9d32d49a6370068342f16755f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb67b3c09d723e85a2aaa15eb6b24072903028402c9eee1e8f5ab2efd470774c7e1210bda6cf2fbdcedd1cfa489507474d6b87be8e058f57c6a8457ae8398a3b8d3541c37804860a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f8f8751d57ed6e822b938595b17a8c9d7694dc24f15fcfbd2f6c4388662795ced00d85ef1c51be73a00f72e1ef0df65f73e2516522d4ad30e1fe379dee3a18d577e758d82f753b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a39f869d8ea2b9c6bc338b500159d4118bcdcbbf969d3b348545f0e467e9ac1bf7a00d9618eb5e0e10fe7695b00c617aa9a6ef196a2184ebf7ea081b5c90028335033b8ba4f82d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he89dee5cacebebd501d105da21bb82dd2e6966bb8f6038bf203e27646bebcb6ebf6130459e4593aac36f7d81a090ec859a9995fed3c42ddf248b5e0afec95797289811c0bdf62f24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f10bca62e1c19694c842e1f4f693ee6346a70db2ea5971972b5d15357f5165075ce97aeadedf73cab06833cea9b0a71f7f261dcae77d72f84ea31ca10cebc5dedcc47aba1b89dce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9844cd3e9af09906021608045952ab595942c0171488e458b878ded5b78aa49c200f27ce8e1b9f5f6544c00dee19fe8a6ee301875f79b6780fd69a46ea727ff9e2f4178adb8ce50e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7d8fd95f3311a1f265bae70749f5912feed74807d02b0559268d7ae223c0af80a7b35eab4f8ac5c5b482da87d6e782691af9250b5badcc31a937d014676fa11017dc97e90d80fde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h623fcd8b2b30bbf95be7ed5f57f88f163d83ed2c410e35c7e9b0f4ecdcdaa8d87b7f7125e22a48fd784aa323e2321eaf5d9f1916c098a849c43a3911c6fd5e1472663fa857556e66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc010a6eb01d351e06762a1a4e3d659da75f578735afa0242ab3f36361abcb5289e9c9ad8bf8957f748c630806b26a73616a6fcd18635d81b3a9a9510b614a5b662dfd67475328be8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93bc82be564a8d555e22cab2d6ddb8b049fd92679b6df40944308265153837689742b5297f6f1f165876f456b9407476bcf47824030f15a43d1caebfdd579904f67c1bb05b260c3d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1e2cf903bd3c716c671aa565b8118d8e00e760e9bf0eaa2f1e57747a7d3f1d5cf69335fb161bb4afafe57346a347f619ffa27651c583a0d839314f5cf112e74bc31d41b1b813063;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab9ae0c49f0998165451c4a7630f0ca140a6f6216fb863b98d638ae9a1878bf164d4aa201e23da70f7b52d9c668491fd4793f40b0cfac8dc1642518218f38adea68339d3d3615335;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7f076970ee312b5ca6c50ed36a34806fdacb410174cef3b5a2d7595db32e767dec8822066d4f2cc6fad5c7d2282a8c616b96d0993f9877aeef092fa091368b595d476d1f582dc91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h110a64cb1b44ee59c8b7ac5beea8b3b98a2aa380c8abda80f633a581b2f94abe902d9e495578aacc678c5510c84a355a554845b167810a4942922d49a95d14c88477427edac2dad9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffd5a1e60095455bf24d16b08fca61f4c7c25c9e7cdab2a66bc26b0b423fac8c11ef8e141c115ccb9d77076cfad9e6a2ea99d4a2e693ab9377493da869bd6691e1d0860fb06bf16a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf1e2aa924c367f1f5bde5b9683534efcdefef36ea910d51a76898deea15371aede97315245a0148f4b19f9912ec43a99ccdb5c089daf0504319d0a98d3c21540595e05963640576;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e381e65c8e1c7b2d0c33ffc4cc1b2d94cc2152a0c52a0b0904410fc675e12eaa9a171134e11959c43118796555494b191f3ddb2ab777298c580554bd7156370a1b743ac2059d85c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd78a30a903324f371329e19d16193df8b8dffe497a79e4bb9c910728c419de9fb709e22e36ac08806ef8281e9f0c0c9d4b112f9ee49b7ab9cad1d863a7b737c262b5e01cf39da139;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93ab44b13cf546b7293c9b814a983c2f7f5f3701baf1f44089a50afbc9362ab75b000ad6a406869c8be39fc206d0612973525a32f937790514befe395e599c1e6a02c0066bddca5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9d911462c480d53b4fe09c83b63188bc6c96ff0d31f031c60a38136f49f45240c18c15069f763358f1a9790ae38db6a15a1e1f3a540ad2f623175472b54b3c0d914630ff3f80ca5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haea35011fe3d2b759b23fa2cc54377af1b0c595b1fe1b324891eec2c639ff88f2e37d75848ef2eea83ba3d21611499e9544e3d7bb1c28633e083d3e9907fa3d0093f57a0b5a14c68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c5f55462dfd8eee7c18f7a280615c7a7c98756ca6055e0aa6d0d156d1b12ef649ea8db14889088358b2a2519f4b7fdce8ec2f1de03957e78b3b14c247b829285da36d8d7929d138;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed47b63c47e3112b00bf80b943b35b2ab27b1b0f0d310fb208cc65ece584ecc8663b92000786887070c66fdd964d7eb8364fe1d9c8a40c5e0c8065baa690ff1e859bd4e3334936f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56ecf1f8001ef507b3482bafb4f7381162a4ebd742295d8cb401916f27996fb29b0d8cf54a37d1fc80cf2b32e3b3660c9b9ba544a9bf608b80860c2d4e198e997d67f1bd2ba8d45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e83a6db8c4cfa1df3066d4439683358e4e3f29566f4946f1f8b93e0c0ea7574bc00bca9045f058e92d7b561184a8072fb903fe16bb24651f333df2abd267027af70bc50a47d6b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1acc06d9a808aab1d494b79bdf92a9a51fb45d83cc57c7ea088575e341b72533f38bb8e83d26641c66138c623f114120e1a4910a791a7afb66b670c056723b5f608d273aa3bc036a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9261a86d166cdd0a38dfbf6d64dc50a17fc5a22047f3af2df8b848ef7fd226d7fbe7a6dc29b16eb1d8250801f1336b24def6d96d0eee37921a4c657d276f8a884b0d10ae33232c75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a39857fb4f7dc37993b4d0bc753505f721cd2c49a7611748175a0828552abbc5bfc1d20db1074e6f936c0519c6783f761f1c107e36d69924cea3d3612c8162df9c6497b896a7e85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5470ef79ab978af9af6c51caee65f4b38f29b02e07f5bbcfcdf63396a8ab934573d7ddeda48c1eac4bcc92549e6c98d4e4c02424fcb3903a24ff10b8d21cad2db5a97b134c00ce3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcef2f25e575df219af4c7e150e0fd5bae49491e6915ca3b70c00ddebcadbbd69fdc27a45acfe12704e9206998ae09e2e44c236a25a8399fa28337a2901a7388291c4f8ca6068164f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h963a00a06125311b8a25fa291288847e4411a087117e3ef5251e13b42f32bd8f90ce23a444eb052546af6304d1b55ce982cbbdb6c0c6942e4bfff4d5852046b463b96fb413a99db3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f23c87cf27c4ba2b5726f23af4d583c18a7a86c358bd601987cd512baaf39a0234a3d891f1c5f188084a6328be0d1578df27570dad971d5fa3db5c2c784de61dc31fc37a265d614;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb99fc569f4128e88b1ed80ad03dbccd2ba5be73d9974dc18938eb30c6f39e02e0535fc3cbe0f2be1a4bffcddbaa84329bcb1f71be7162cdba178d0ab7db04b7264614869f1578b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc68d4a8615863d71b5fee55ca89a2b4d5d64453016d15672791c476142a0f41cad3dfb84805ab12d78750960a8e1c0ea079f118676de4d152606640d52bf554c66f90d783eb4c6ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5771d39fa5a3cfefcbefa1e48e9f5be28be13e3937e70a9734fe54f86e43ca2fe4d5095d3d9d7c0da1c1251faa9b8dc5cb05a28f88cf3199436b8e2861eac6f8846b4e2c77b84077;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda42725e54cfa62b533cc82923af64f3b01516b935cf64106aeff4b9271d26e99099a4e1dc91fa414e1a9d6fc5c4d92b9847ca416b1bd21241309d1fda5faadbef7d29b0454dd383;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a3c75960e3d9296b84e3c7b05e7150028355d37c152fda57191107599bfbe94d00768c6e9afe05e427917b4a5f3475b2ef3d670eb2be6ee1d70ca51c639465c7c21fcbcabbd517c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19ef9c680e64b852e23459c5ae67abc8d8465c7c08c2e553078b81b32f88b4c8c2cc78d855e027bf826aceb72cbebe583ec620501adfd7b6730ca89bb9b57562bd7dd07891c7d0c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d89f9316a19df309ba7f737d97dd3c642931ec38a4858b2840a5597a587828f9291bd40415a5056c7d1f3b433513880fe1bf974fc9b36b3155a8fed628d6126bdc7ec2716706434;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f78eea59756e2b74a46c55b10f0d9c40a13923e93730aa8ef4b3e3d882f24a81f53df6ee41102eda0da22ba8db8eaad526abcdd5a4520a5511fcc14b10e3beaf212f589d3c0e6ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60c39c75c5117f68c0c16ecf627d947c39bd26b2abe96da3ff778629ef455bd2a091ccbe45c676c346c86c1af1f35773e283e6449e906447a8d713084c0471073c8cc39d7a74e8c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2172bd9479adf4d9c1401dc3b467d71386541154ff20f29c652859b3f48ccc5f6cdcf24f8b2954c9989f7d573ae40b8b3ceaf9077fd88ad78d6ffbb560031add488a875f064bf99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb03c4b7238b3ebf08ae72f824bb4a6e4e5e9fe2610830c6383da2ee13ac0805cac3ea9d0e758edf107145981cd4632e592dba002145665cc53bfc9500200eb2274efaf40590b65e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h221b43bc9eae05f8e6583f502949c435b3d27828cb0032a6f17de8f41103b9c9b128eb2832da26ea02f0323ca439a2e004aee8d5b06caa7d5d5da0aaf4f22b10979876172a113f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf7d0fe1272a1d4e17ed60cb9078843dd6cae0137eb0314e2c52baf26a00e2c3d5b3117eecec9deb38c0009f726ab95a28b9644642072d05520c8faed391e7545d206c1c7b893a3d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fb80eeec7e13f69b65d17b5b6e8b6c7e59d95ddb24c189f1d3f267da0b993cf5d2a89e83f8bfc53a6dace7c152158881bc064a17156ef6ac0d248b2f1fe332220f4b385022120f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f0584fa3eb502b54b30a2e6f0cfe2f140a1c7dc95f618c02ef188b551b10dbff705c5c3994322567538be0c2936c94de2eec0f6172b74e1733eefbb4826be7678caf3b6821a9bf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d322143dcfcec0a165c47f3e6001876045cca9ec9bc893fdcbe8dfb6c694c7378353267362fbe98a6577e0a2f80b092e25ef0f8a7e6c04ce99c24fc6dd9b4d6248a8c9efd59c118;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h751aa00dd334b9607af52a2708dd405e76549294716965d26f656c2c5dc1b57fc22dab0ddba887a478a86b0ee475196b584e6f0e552964271e1e519cb041a3c2e5dad23cb17b780b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4379ce2b00c05e6b9ca7f5ef8d5ef1bee610f15d14f0e4a9db5944470656603181d81cfa3d5061c5f9ed42a3ab3cd1ca962061ca4a2f80bfbda41db4a9ee2c165794bb95011aed30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcb9c4bfdbceba7f735e7b22e29507529503b421668922b26d202f85d2deefc4a6111db14a5de0ce349d5b8accc8f378ff67379b0302926cb28a8bb254119fd9801a1be288f99fc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h569819e95e1d6bfc6e8d2821ed23ca33f8d3bacc696311602d6cae313205b1dec30f915997ea7921e41b9d62db59ebfee692be3a62d73bbffc14df575200cc8f9004c8c0a34f74e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc19d5bf53787c7497b8a3fba5a9dacf4593f67cedaa3ae10b0d15ca990de0e2c30936955a85f0ba45b5923b5a27ac89811cebb02207e388ff45f89190b434a5a26005761462c7996;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe37f04df37051c9b515d423835ce93bef8592925fe1a5f4f58c424e84d12d9cca2f82ff61020e92cdf1222789d9701d33e7dd61822e28be0d0df4aa8e31768dbeb4caa2bc3398eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b6c35394fcc72b26d004b8286317f0ebb365bcc2fcc3b0dd534588fb64e99341da0d2bfa9f872cde45939c451d15cef011ff7e29def07b14720be28cd6e58b5aea9f695cf53b7b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c39c3870b9d2335edcefec19ea091c44ec477dea7adc5f40a58f07490b1d880cb71511d81362318b857c142673e4a5043ae88c641f291f794fca1b8958271f3a4a9977645e21533;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97685b7a0998e0bbf7d6ab6954c2f604429b8e124acdf0ab5dd1b105fa5af175492d91fd9c8a2d2304d4134a2810ab1d0131d855079e40d84ec06467131c74ff976511480f4f5a17;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha500ad6d0bc12c52c8c46c46dc888b766053d3f50fb3e6d4a588d7316ff9a395dd006325457576f1381ca23fb223d54a110a9b978a23ad29fb1bcc41caa26677ad1fccd3607de184;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb64aca2e5e7082b6bd973fd1f4a82bffa1a4e862b91bc5f1249eaf054470f5190bfab009a57e036b27922429a69002b4e248547bfdd38e3f168c45e7a633726ec0cbefd8fdd77f03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h123593f657ab22ce03375d76a408a99aa8bed1462bcd390186fb691638182f4cd3811ef81d1edd084aa40ff0fd477e319691f33d73271df219fa3a4bd5ef06a82e0f70ac53640ad5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd60ccf61fced84e8a212f1f7408974791ff452abe8a9fcc2c5bf29e23f20f1407b4c4062f3140edf39d7b83698dcf9207dd1e650f497c0febbec8d44f661bc489551f14d6f579c6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h871710556f1695aa71b326566157cfc9a9d456104b7206d9ddc309496e0fbae5058ff63effa4c777dd8f6f9aa2e0663f214b130d7fbf717b86de846a63517d7304014eb90722e2e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed7f0dd5468099df68bc7d8a9562686b13d856adaec6d06511d3896c64f9c91e258f662c4fb417788ba7c3b9a0159261c30b36068222b2c36520f9160e1b99b585c19b2bdcbc2345;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd83afad4e5f6220451d4f9e458376d783423cba3404a825c7246f27e145e0c16a27a976fbe830e05ea1c28b692c01f0cab4b1e5de55f926532dfa8bb7b5d22048f59c115a9c6d051;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4e8eb48c6a8fecb37318d17fc93ce675fc28e68764d5f17d2acadf44f31aca9bb48a833ca1c6ec605105c8252284247f2d5378c8ea32f52d80354e3d118bf19665cf36731990f77;
        #1
        $finish();
    end
endmodule
