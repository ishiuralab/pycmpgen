module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [8:0] src10;
    reg [7:0] src11;
    reg [6:0] src12;
    reg [5:0] src13;
    reg [4:0] src14;
    reg [3:0] src15;
    reg [2:0] src16;
    reg [1:0] src17;
    reg [0:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3])<<15) + ((src16[0] + src16[1] + src16[2])<<16) + ((src17[0] + src17[1])<<17) + ((src18[0])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8de713e020ed6dde8a257c1c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h450521b7ba218897e86287d96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ed0f7c581dba60f529f1a6c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha055a58c0932977299740d4b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c8c6995c1899f38402be732e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f24637e900d8a4c9a99032c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3beb806234db35a1f85117f1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9daee54faf88c52960b0c4036;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac055acc9c646c1226a67b680;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f0042cad154e060adb14a292;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd05d0d1c8c25ba788eaf48890;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d98b83ae36d458b0c3333328;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3494c6176a5d85172104ad07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he078439dc3cab10478a682287;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60e0abd26d63ba5436de945b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9ab97517fd58722c1ba963c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82236046f0b189489a53b53ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8e188e2bae3d0d560933e31f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ac15107146e49f8ae4ac57d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef14e64de7e8f201457ac4ae8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64030bd01aaa0add078b0c5d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14ae1003269aba8332be636ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he25f1c794b3f1c0457445c4c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88fa4397d5575f53aa31543f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17c932b4d78ce97bc68e01d64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefdf3eb41e95a4880448bb3db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d43f7c3bf81943f54e4233bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h881d93b2cf3a06e5ab37fc960;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc069b8e40e9785e0c25372a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee054a4093e63131afc2ffd82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd14b9d9abef50326c9370362b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42b32058953c54feded48c56c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a103034f95777f97a0c80f44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fd792a88d1574f56c6cf5a52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec8adb8e1dba202430f8dc700;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcea8802056bddbe79d8a29e59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a04ca7d5a1c9cee40d9d2b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h766bb34a16eb9612c247cfcae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48c531bd320d93b39fe09684e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fb8c9a8272ae9b4b08928062;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a7dfb600d39c1b63b537d44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd5252f03495a01598403ce7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9acf14b5abfa28ca81b8786a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3a420478a63ac80bad75dcf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83c777ef41f57041842216348;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c34ceb7902fe3e345adfdcc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc85e91d6aedd1f189c64a9362;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33f2dc3af35f838d2d5d8c096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h422593f64aca18a4d502f809d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef8c426869588b6556fd40197;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fbf5a31020c7382b7239340f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99fc8801af1cc20d573a8f96c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8ca28fd3a67b050ea6ad27f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f680c7c968f991a118111350;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50bdf864a81efcc89301f2982;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86ad2611899ebadeb7a4dd7ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda0ed6f790e399396fa5d0664;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92a0ceb0ff042bca6c3f388c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36832a75427ec4a2ea35b3088;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d3d783706739a161a38ceb81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc28937d150212c1dcbb7bfe3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h868d2bf5c9b6d83cd945f2e57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h432bafbed6296b9b946d53877;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24900cc053925d289ac903f55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59086e23306b91da5119e9ca6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd22cb722d7fb5202329601349;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6fad1c0922a1d29574cd990c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39d50c815c262bafa2cced8ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb9e957f4e6467f9a5137503e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaa55b4c8c9f23ae37f6d1945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89a786f963a775bbd5839a2f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fc6240b61e04c3ec5e706b2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43d07cf0509f7dc962b5b7ee9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a47fbe82c2fcbb9ba9463624;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96e6b4fdc6abd4afa22e9d9b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90303aa6a4ead18c1d416524a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19763074feacac05a1aeb4fc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cb173deb411c8fdf8b7e50c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65ed7dab95e92613f04afce32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b4c4790368adb53b32d2c9fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h934f2454897a68c8a73ac8bf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cb383b1d477721240597dcc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h819dd98ee5fc714277062d09f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d2f679f8a40ac5305febd4b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h756e12ce1fd390e8f82e81310;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c3343ec00613d0810d10c9b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2684296c842dd5420113073e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5eb61a4f5236c5a3f4241b1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29de66b64c2c3cbb6629a2057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11acaa820566a68b4797691dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc80f0fff36b17a3a25884d2b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab3b5625dfc30b46da9b991bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2222006da96294c88a5a43b4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc4f3d48bd689aca9617dc789;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99f543de05f6fef3834d3be91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77c63118d996a4ff79172c505;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70617299f6e35d6b025935475;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27118e78d9444011fe0e8cda9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h434ffcb009326ae7c957bb906;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0b4749496775491995f77dc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha835d2efbdb075f404401f7ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc68147d0c3d86736d8366b97f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2231db9652c0304af0eb6d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cbe28aa6fd5af542f473345f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha153c6d15cbdff0c454f98f8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd67794682ee2b9a78e3c3c922;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h712829935e5e0e587e5e9b7e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9feecffa68a66af86698e65e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a34dcd23915dacd7101a743d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf870e49fe0be5b2c7d6009db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2f1607f4f23362e69adb1091;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86000db674efbe09dab5c086f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6393ce51b276eab766f79fcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31068c695429194b4f506cfe1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2286649374a64ffd42551b32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb26fb78695bb4bbb6c3f5c1b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h161537b489b622a1d6b1b5b28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97d434883961c73d67b1e397f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7293328727fa01b2a6b6ec42b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d7e0f79d3658ff9ee2e3f1d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3389ca47a27f7f64fdb7cd0b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69dea6f1ff35299e800a3a603;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8adaaf00cff1ad2c2685a05cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h436c091cead05777639d97cfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h319f663594406896cf2adf93b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc120fe32fc98cb59b9dadd1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9917a7e903a1fa266298b261d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf500d91cb1d2d421b621eddbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0617bcff398b0cea82792132;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h179d3f61283c45dd58d678c2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb848e4b91502ccac8075021ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3de43e3be22d529caeda9de31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61f1dc6871fc33f7998581e3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3234c546a6bf0b600a8d0ad9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb37afa5a0a6402a3506dd745;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h780d86029953078dad55dcdfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc979e36e61722faa0d278cd6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e8510819fb443071cc8659e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h963896d71e8230ae281774477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2ea55307f13adc951abd2e56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb70fda3e84230b3e5043b9885;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ea42ad0a61354a350f7597c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99a26a83394477a5e65a0ef78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d07ab0313663de1dfc2485b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3213ba1d7a0712578e493f2e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2060f9eb7cd524173a7b6197b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78076dc1ca7535059d5e1c4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bee3984fd99d21c4856520fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67d6e43244506c58cfda0e706;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a3d47e367c74e791374f313;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab3360afd1175c4656c82dde8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8260b4e33a68914089a7f9421;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2199c6c135ea58c1daefda328;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3d2bba0c3589c20b5eb3817f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f5b168df55f1913c54a23bd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2eae86ea1e66709ee58d6a37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d720a5e7b39585ecf370a402;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a07c7bd79807a6924368c6cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23421f58d2341cb525c5385fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b4e1e476e5a883449953fde6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2418e4c6ba34d8008c2e6a0d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2091e1a784d0781e155755bdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha32f6d3cbd08ab4a20593ce4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c5b7d31cb5ad943eea6e09cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f0d5c1645814716a096e94e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcca0e1034e355baf20e80a87d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h150c1d3bf9b83a4dd501f2b35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d22261be649375dedc0f24af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h735b1a772c6afcbb8c40519b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8032548b09fa2601e7167276;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha60575f1bbc3d1dfc766e497b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf986fed1d4a2f806d91a7d6bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h653df3fe3ca45b7372d5c4d97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88076cbdc6485323a90bad8ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac30e0417f2760c81cf10ce46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h314aa5211661d64c7776103c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c08d595d0fe9c4eeb862ebbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda18f984d62545360ea9b51fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3866e651a8796489255e8f51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86eed3d6af777af7398e613fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h270684d31280423dbfdf9490f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63c88a54586cb2234dbd46e66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha59df6f42fe472e0da79627b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49ccd19a20ec5778324f373ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h751b3ec557d4ca2bf2f5aa86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h658036535d090631088d6a427;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b15ec9fea7b9f567f86c7fb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30f5d3896ce1707909cc56eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfba2bb8d47f83deae7c51499;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f02af12189c1965b17b16b9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd48cf6f846e4c4879e9b8970;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef3d9f6204f53268c77313726;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd3eab424d02f9e7c2cdef35e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aca6f825d8bd13358158c110;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h484f42cd39d76c51d6ac0b384;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63de9024bc64bebe1984490d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4172a6ce72bffea471241fc93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21467d8da48de32940fb7c7b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf63f8880cd992bd60754fe777;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfff4143be9dff16c1f63ae00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80f770333c6bb7e08100c226e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6dc78d0927e95dba2c18f45a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38bce77223083b4666f91bd87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h648be51622c68ec1503392b65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92cec60a31ef3c96ce942f608;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8336bed9cac92c2e2392db34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h896b7b71e6aabc7204ca2b94a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he69e9af5a561158e7cd95c12d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6087f80dcab6f4559db0616f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba0619f5b3aa4434a39824273;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcb185912bda6bb4dd8c97308;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd457ba9a48494acecddc64869;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83272e28bea046618001196cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5f16c7600077f1be40d16984;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9b63877a82d613d5ca18cc1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e593f07ccffe6e374522252c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbc61589cdad7d1ff620a31aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hece74ec6e8c3bb676dc017f38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0e33b7c02fed9e3f49ba6cb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87213cafecc50d1bdef7d17f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27ffe47150d5a0c331c456836;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbcace7ac3a2b9084bae8c9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h743afe1e55b07e9df92a3428c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94e05351b0f60eafc1502fed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hade66a7c5db0151c3074b2a02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd28676a2c02b326cc102d77cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb31ba4bae6897ad826e657bc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b0bab3889a31ad3fcdfe1a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h738f699ba5b62706b7f0844a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0348902ce242ade0c10ef2c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c1217c8802b4bf08677a3b55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he367cfa019b782340b27cac47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb85d5ea1baefb3350561fb68b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb43d081259d76ee194f7dee89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h207816e87c0045618163e6ebe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e9fe9debdcb6ae9cdb30cc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38fedeb22265f8e9296de93fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h510a24174f09e0171d94ab1ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89aaffc58a05f2ecf517d92ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc76e90dc021432e5c746e0eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he195bf69ca5efe3d2fa8f2fda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f78da1e301f850292a8eb178;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8710a24255abf74ada51fd8c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc8fa672223f623c949469c36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15685d9201cb49b02696ca996;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f7653f5c35da79d00426d510;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5d062a59f1bba816ab803036;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55c669e5f2fca8ff0dbcaf4df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2ebd2353ee5a445c25560c4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b067d1d0386c9c23d10a1f1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd419e50747d604f7c04301a64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27b51bd213307be2878c07707;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39d9bd9ddbb0513f6d6e1a025;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1783396d9bc41f7b6f2cdfe23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha66d670fd0151fcfb3e9d88e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbae381a47e4acb294fb132ad9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h857f22933ac2fd036b01269b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4d9c4251235c31071099c07c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e4954960128de1d92fa4b4c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1b34f14f1c5fa574465e50f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5794c45912fadb88a6f4637f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9de80f1a7acdc33747621235b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc754b056ded9468dcba12233d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf007f8ba46c9772947e74e9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9be390190243d0fe3e7972946;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5d46b497f081ceabe5026677;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h415405c80ea76bb413eff7aac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habea9922cb0ab5479200cf6ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h919455e997bf9c5f8cdb1eb33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4549a858b0495dc6435414a19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf8a640746bc5a7c708b76dd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13df2fc588b2ff934789f1ddb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b3661b95cac5684590735adc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b90b1c318614443451ccaa2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb965432372f56893c380e4c6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7065ce9593bb5e91765899e5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c2196bfaf818b2349a25e6f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11d2b7013cba3ccfa26f176d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9ab4d1e85ec6bc3ee075d9c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11a54c984235c1e81eddddea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b7234053b7bac51eab570c9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h279131fcd25089c755a8c6cc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8c853fbbeaa38abd80ab80bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95139d6fd421bae93c79dc7a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cf609609b2107386fb84f9e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h637dc5c7265211b4004709f4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75ba2e477d7bca1cadc7c295;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec30d0dc73ff7bab18ec4ae2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39fabd014ac518898f1e3b842;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19a953e223c1a55ad60400094;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb7629d8b1bbf86ab3816a16d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb882090f930b979c2023f0c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4852c00ffcf05a593f00aaadc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b4d56aeeacd4ccdbbff8d688;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d78ac5734687090413193101;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9c4983c7db7baaec1ef34530;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4772941e49465f3c87ccc856d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d573c80e3a1300d0a476b897;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfaf1d6ddad9083355c9ec7fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f03c987dd73a7454f4bb241e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf65311871b7d6d19f7422fc1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26dd74af21e8fe822275f061b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fae80a441aacc859f43bafc7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8296f720922ef6085a64581d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e2f401c90dfa5b347ae7901;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8f3567707924fa6b42de9c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6921aa342924c0ee62eb6e75a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h299f649b5fa2adb761ce5e9c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4d03c0126495963a8d8fcb34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef60dab5a953ba48e297a317b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cd9c285d99db626ccf911fe2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e7c7668b28e70ab422699caf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d1f90229a8b5a36d6cd66db2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e4532bdfa4ac30f13e9e5d41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4e9c11285b612edf5abb442f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2cb5ee2db6b6ece1163129ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0a46417893332a28b09a3209;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9de42d017dd2b3f31914e5997;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he46e145218c6c97a10b4233bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c517b713ecd80529ce51a5ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4ca9151134dc16baf743b44d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h278dbebff02755ba97ca1e7c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb98780ae528914ba591294a15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd68818fedbc5db932f8219ab8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9521dc3b69c1a64d723e9a7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c91098d01164ab9b8b7e42f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4b690eaa4f4e4352f31411f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h914a1973eeaa0b997d9eb48f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec9496f57386828b33b90ffe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fbe6978056f1fe64cc3e3641;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa193f14ae317b9e3a9f407ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4d59936cdcc381757e01b78c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h932c51d6738c5d55cd4bffa68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cbd7b722ec21c64a920a1b1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb108dc3366923f4d7199684d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2d47f6b91cf6c0303042f569;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9698bc21e467eeebca80a55d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e085797f17dbfb6721d97026;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93d6c36fbb574c8231a923c0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69a09ece11d0e49ce9c9f4403;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b91531436dc69fc95ecb0e3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9702f2f31e54bc9849326bf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb57059eefe52a49bb19946456;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92a38c22711fa645672664241;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd142ce20e804078f8ebf57352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15a74b902cb0739ada2d13adf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f087ecc09f1fbeb9fa8b2fbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8201a8ca4a1276523762757fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11dcc438148e5890d97c69e15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdfe15c122931731e45a70a72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf09fd499e2020c55deb86598;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ec5bc7d02f398d66cabbba80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had175b61fa1f5a7a2f1a8b503;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha53c6c7ce792a2e730b56b056;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9dcf6c39f357a56565122439;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fa8aab7c3cb04652a07be7c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d912c754ded47d3fcde6e0a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19a186c82316f698d741ef085;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd590229d5f8c69a0bbcba6d48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb447d9c20c4a8cbdee10b61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3c7f3593d65f3610f2581676;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h962055107d87641d0fc77d954;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1780d5179bd31c2621471ed6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5481d923488d91f4947d444af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb312a3931d72214bdf6e49e89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4397f2fd56f893e97acfca35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0b49439d6792f8a07a0925d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf43bc0283663c433321e10692;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he558ba9e268a7432e624f7ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6710d619a01ea6c4ef9203108;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80a115ac56a9b0fa64338c71e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51b0951f7772f3e5d38f2cb25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73d11533e64089ad5602e31b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca0d0cb9199478458fb95abd8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heaf0e78f075fdd863c014b26b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ee5f6f97bff55467ae3bce74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d78792e8fa1dd11e556cee18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b899aad8a1547b8dc5513bd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9ffddac8ab6bd15597c1ed11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cf891f6e3ead382287d4a0ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e18a7ba29bd3cf2275c70454;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f45804bd5b1e8333763e7923;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c8b2f8e67d74b0b70fee721a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf78a862f2f419028511068581;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67b9d33d391c82441d3d244c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fc8197d26888c8f392626b2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69982a8272962f17eb1d1a566;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h969db83fa0be9ac1d6cba61bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3341cff0222592b9a18c6dcbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4c48c0be9e48797a8cec33dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71f71efec8c87f0c387951a16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca67c8bd026b6c4ed68a6253c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2b305a9d3811c8d6529721a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d63a6f064a3a23c6c5607d6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a476dc242762660da38d6ea8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea900c3249862bc8be1a9eca3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd78866723d7da1986bd457a1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cc9e35ea161196a601b15f37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf274019a5bf47b6e06602f70f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5762606ec2775e035c20ad54f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac60e8e4119352da098d8bd36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde856a5b7c02b26cc2ddca5e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5926ad68e9f3d43eb77a3b3af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb850294eee4cd3894ce3d88d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba235ea9ab811aff9caa47249;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bc9a550d55bbac7a50bc6bdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b20ce10c4cb362921c72775a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd5fa1790443cccf5c7b8c80e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b59ba502888c788c338a58ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb6ee6efda5cde0cb4af24a47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecae6c8af2a29411685676631;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf280115c1c2629bc39078232a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e7ae236ac7e825dd78d581e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h148c25f590e46b6581dd2ef21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc85da400b565cbde4080a21c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6f4fa850322521e4b6ba495;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7e71020e6245f51de7d73149;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54053b18be57989e4e5ead262;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a7b44b3fa35cbc430e707717;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h354d13766ffdf52aa2221df7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfff03fe55c3e42f43fb8e734b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h935bc75a7ff8971911d2f8ced;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51217275e190d55290cf7df2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bb8def37c4eed5353461a1bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d78d42b8b9bb1040d2bedb8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e82e91cd054df7fef27a3f12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeceee3aa79ab53cfa98d3d2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba458ad5a9846298343de6a3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56df0d74024eb9c49248f66d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1addf5e29c2f7464de9b1a55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf296617d8fb1b72edce3a79c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h446fbbb49375b8185c1d0fdef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h551b1406a7263740fe35c98f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb81d855b1a23f2b471d46e6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha26f203ecef5249765d268439;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f8106e15f04c0f8f7ade368b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h969d15d6ba15355fd7b4ecbec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35d2f74a4edc52fa4a23a8823;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9121f544e787171a912225a5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2700ec1f86a08ef6e4cc9238d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2876cabba947ec44a293d1cfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21cffbccb30d15efb9a8c645c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0ffc3427c49ee8dbf413588;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9735d647f7eee6902adb354fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d2191639764c6db4569c7819;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c32b02cf049f1a179181961f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he56218d4a5512b8f77af4a953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30dba3019eac44762053a3d99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7394203031374f7b777122fd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h809d12df1f3f20a3b49d96451;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf09f2ee82ecaf7b3ae1905e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6be61daa56a49eee23568d9e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbe9fe52d83d0aefa5bd9fa02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc19552d2a850a95311d5ea24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b148e06f8b4e4e66e6164b3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h892b5ce12043d908cbb2dd439;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42c477a540ce91305087b2477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9d23d5f652a1bb9df205803;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f9570b34596060bf7f789e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5b6797f14d97bf8cfcc120a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bdcb09651a4e8bf292db4630;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52b76fc5118717b5798520e1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45eada5cb81a5063ece91c257;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h859412b1ca27da73d207b5fb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h480070a7ff15f503e60d4e5f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fc2430d9b6d27e2af52e54e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70c5712d24849b242442df539;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d347b3274d4d1447abc710f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83dc93e1926d4353d4ff5cd65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd092d8ac3b8296a73f1e6f83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6be7de9a1337793522266a0bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8946e32391c93b5838cdc24fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14b24c4e3714a7424548785a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ee0611c6d45db4c06e47523;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3309742b3e3b4ec39d2646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8233875090e4efe27eab33563;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafdd28f43923328b43b56320b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7201355dd3b055308c880df16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h339207e49fd4212b6875ea98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h483e14bf11c6e32fa0665bfcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf26713568ca8a05c6550318a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63021c8ceb13efd3abf855784;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc0593530e00e38dfd8c797d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7566d7cd432b91132a87141c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h622503b309924ff76392b046;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9d17679b08aafd16f31a945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb753aaaf94dcd8e1dfee32787;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1531f44dbace781c07bcf31ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5f9acb615acf4d6fb1ac914;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a1569a07c45f584b42b1a463;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h732d146590b10ba4d2cfdd94c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb6a492c3a9e058b72e7959fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41dd652d3fc6de0075eb3df6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c3a80e30f967b2645cfd3bff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea1274264a4dfaa4560ab62ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98d3f97549beb6daa81924710;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ca421b8234a7d19f5f4a34a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60aa16e78ddd1f0223514b132;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfba8cae2f2b41138bf881861;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a9af2cb504a86b36c2a925c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf59d1eb8a9918282d54626b1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed8b49fa4c978337aa5d69b1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfc57bd10d77a0a628526ba29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3413ef1b42a7183e644bb7f0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30b7e1e2fe2937135faa2d854;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8d702a1823696b6e8b640b42;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81ac9c2448a11e7971e6a2418;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4901c8c4cef5bf11f773e9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b9bf01ee1162258bd2f93e1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ac6e7c3818a5bf8e98fc0de5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b2f8c4339931044c983f4566;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf704ec7bad8279d42151c3575;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29d88e9f8de5631fbe0bfafaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heef67e59e480b2e1c4b15fcc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21172308c9328e771a71008ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68e78068bc8eeb6772e663964;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52cb2ffd922a446238df1bf93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h903170f0853e637c347493736;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7452169685879c4d93dbaadac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36628169757b0128cc25c12c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47b998694e53cd8dcb6c2a5fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ad734bd51861eb9ab9620bde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94262ac399a11f799c35afd47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hada66a99d32433616b440dea6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9b47778e20d8f82e1be9a2d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3754d3c730465df4a9a2787f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4a32be0c8ed03338b99a7397;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21890846025b72c48c027fbc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ae2b73731dea4b553db9676a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h642a87b9e74a8739300e0c00c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fdb2e35acc1022c79252e34d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3810e1d1caddeba944739f973;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ab622f00fa14064a73dc17e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd13c2ddadbbe456f2be63c044;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4a88772a291562b8391c343a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h793e1ef0f16bbb669c4754fb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cf424c539091566cfc4ec6b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3882a4706d6525e82a405eb07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f4b40bfa56e46323c6212892;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he73a2208c5498a53dec8dd8c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha55a091cd9f845c3c8705c42f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dfcd9003a07feb869ddc2f53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a3b9b241c5424e03dc03a860;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb941a7034e142714fd20d5ab5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h773de2b2674def17e87d8a65d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcee767f3da2c2e14423bb8ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83c8529d321937d5e95f0ec5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3dd670bc78ba49d59b2f7d45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc282355b7647b7ccbb5f2f9a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha266bc6ba648fd6cfdf33d46b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heec1b333f54e4e9b1993fff3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9ea401df135e0682ee173ce3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca62265cc0bae9a534a052593;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b5b88095d0f63f006a3c69ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeacd38daaf457afb869ace91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca458f3b1ff8c38f8f6eab041;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8e14b9c71bf6397005b9ad7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0718d53b4e807dc2925b0976;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56709937508bdb38628e19500;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h592f59c227a32fe79a2e760b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc53acbeaf0726137325f9b370;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53f2d9a4e69b68f7c7f8b11c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c9c45c470b1a1dbc17dd61c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9146a9c2ee44e5a31f2b894e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h433462e647b0e99b50905da33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84d31f34825b868b706b493c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20df5831b5b613ee88d302417;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h779941ff397f8b740c209dc68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he79c6abb476c9560849b5b143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5711a58c30cfcdf293106b2a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd835f54460da541a65f88bf66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h607a71c20d1026ab929a6de46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d1207fe6739f4573c425cfc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha190470c002e2edb38d40ca6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50d36342c4a90426de41a1ae6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18ce69673ce45ae5a8c476352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0352d7ed8339c737a08c590b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h179f38b7bc8f740006d0e6108;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e7ffff33b74244d0436c86d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h919f6da3d80319eafd2fb734c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe2d023a50de58ef025840d02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf11abfe6e9a226b312d6ba7f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6a33ba95288624754213d993;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60626718c8757a333f3e9b6e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb88b376397ce186557ec2721;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff57feced2566b456a28aa5aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd999891d4bcabae752119bafe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd1976511ad4231094c0646c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f5a1054ddb46a16a6fea0a4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16f01ab07dbfd53ffd66c5baf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd09f0bfa2566bf357e8284841;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e7637f1d2fb1706d9a73b494;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6ca8356d494b8751fe5c6d2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96a81f4bbacfa5f58db248cd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54af75a267320a725877699d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b915b3747d02b788fcb48937;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h373efdbd0ba626d0542ae0610;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99571abe5eafff6b497c9906c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b13334f3ce0f5af3d0c4ec5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b77492e55a7ba9386a0ace08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e52b57fe4dd64ecff96b9c19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haebd1a57563d9de5e30e5ae5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3464c6f7b138acbd0c71a5f9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ff86572019146007c3390744;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33b4096a49ce7d528406ebfa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h426c3b453383cb907754fed50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc562e2d6ceb076801bda36e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a68ee13968b16a976848c2e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he53dc6c05371e17aa6d9d18fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ca073637973afb0d51482d62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28f45e0f1202010c6b2381d60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb77327495f74a751f7137d82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebf221a6242c262b2c5fd2b19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff5f4638b95c28f5699f7455f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf754c47e7ec8c36fbb136ae3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66d4d34374152affcb464c6d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2760de29eee481615ec2003e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a1b006ee1fae0f172069e539;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b988e1672ab9823a617fee59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h671b27f25cf355c6889cc6d3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7606145f760bf9d8be5a101af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83f94702e6f66054d00b09019;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a0992b7d8203ce41cf15b419;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a5e3856c3d69dccf4a930195;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa0dd24d327447c1d6b5fb28d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha66049445fb20a2a6d32cb29f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7dd279580ff0db7ad626495dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d943137d04244622369e2772;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3101d0b2beaffa8a3fe40cda1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d36dfb21c85b4245c7b8cab6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12274a53369455d517f9c5061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1215452178fb5277a31518e00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed51b6fc4a2457426d9c8984a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f4ccb4db0edadac9b0d09e27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c485d5536c1fa4a3e63cb3cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a7b198c80a90efe4c1dc5b0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb7286b079e7b64b039684e59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a70dae06c533e601ad6a4dfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55486da7d8c0db70b0d38aa80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h513cc15d371bf577578c8c34a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ddb34dd1a014eeb9961c3f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa5d118340a8a7c6ca6dc7ced;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d1a913e578e240c6cf16c50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed928321233ec79fde5521843;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7976b23cdb0fe634f3315655d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6aef1717b518605ead99a2dc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h150d11ec916d72b4b24321afc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4eafcdb41c94316bfc2a0cb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h180cb15a5ae165c1e7161609;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc19f5aa452b67b1e7b83e95d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7ca2152207a6e72bac85b56a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98789ad6105ed5db44e0c51c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9532bc9d64fea57f783700c89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59f26d6d11d150109a8fc9e32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca6bb09a93f335952776643ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb86372c0805121c8669a50ed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac4b4b1f667812518d7b714c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dec5fff98c620d816cf6cabf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20e5749af3a4939abaf8194e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h108e5e50ac79ebb296b7a2b86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c8e41332b2182476c8770fbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84b41c2110702cbe4aa7f4fed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd00c11a0149a6c18d31383747;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18597954de56e421ca7eefa0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c9a4c0eeb316ba4c2a37aec9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21b2bd7767fbf125e5d0d2432;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa460d6e76b8af902c610024d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78e0d86f847a75516e5f41a87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22f0d9c4492e1abd6660a7d65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c19bf912ee9a7b988c31edf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73bdfc6c0c9fcdd79f7844194;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11845825a2e0cb2882237fe6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab77b271489c6847d08059c3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e8d41298dc6a2d946c48e88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8748953874d1eb04988b6b7f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba32da35019896d73589f63b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38880819ed0c2067f63039298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h300e6c82f05144b2b0b61541d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f9e8625c018233db27568e70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf666dd5cc015271e6fa5321cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fc5677ead5a70019801c83eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc3f09fb30c336a267236c6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83d7de121cbbdf2e058235307;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32819ac92daaf5c73fd6974b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7d65e32fa66287e22b9f5a4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3dd92edf339f9261826b5280;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h459533e6baf126415476998e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a9bda8de4c407f08dc8fef55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37ab9cbafab73753253f51e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h269e5b3d15bc9956a57d7a6bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc157cd5585d9a25a9cf890ffb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96e9458cb488c5979b6f2b8b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h208df745b23d2003c6f311103;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h813e130540c195f9cbecaeb6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b88e877e9b1ddc899ce7f770;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bfe5c10db1fa1079902ad0e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a80cc443db73b0fd25b4d4d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1ba08e9ab83df2a1bb3ef445;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41745ad3ea72792485cc75e62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79ee5fd4c8b61b833f50eb15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3307361af1bbbce094443479;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0f69a8915753e65ff12c54bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16bb14d3b2ead35208044a461;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74d46eb621175dc3b908143ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e8b1853e57d7b383abad7250;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51eb1878c9281736564c22d50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he66645621a3cc16e5aa4d79c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4aa9e908261f270aaad6d1a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbbc8be75816f6820524d88f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h314132baffca09dc9be822c19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h246aad3900df0389ccf8b1a18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37f515a8383e0344745c8e364;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b508ce20447d7c83627708d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1e81372a852474dd979fb9b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd11a21567d58971ef8adf8298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha75a7b1e470d7d2a410ca9f37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h192ac1dbc3238c35669349f98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9690ad9fe9dcb6cebf1928df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h343482d4b5ce4436da4dd54ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a45f1e4c9d8696a4b0a79184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2504d33fa4c6a3101a1186d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5ce12baf61cc02bb51992c0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5702d38e5c4e1ee5be0a3aac8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc7d0fd2d80e535d824b37859;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33d0b5bad0b4b46963323fe02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb64eed912e21ac8155a86bb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e69d268fce3721fdefbbd846;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e71b2f899988ea03b7ed5e05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b386ffff9d506d172baf8625;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55358b06998fee9c51dc2c540;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he602b60aebf9398b3c25926aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9430b47cfbec10dc29321c6cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35c4fb2e135941a5ba1f06a08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fb1c09e039118f778620c11c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1231f86565bed189721b3ec65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda0564e9064702692b45d2595;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d0ebce3c79c190c6e8c5a426;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15b17d16de796f7a47a654336;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f177ec0ff48369f8f4a3ffb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c841efe552b8a855a49cc450;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h974a058efe977fceaa763500b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h388d01c78051094976a2c80f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc793acb4b4c4474ca59113eff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4acb1bc8a2dde1eb7f40e366d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b18922091cfa2f907a502281;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2602a26d47be85e4a03b048c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6283917b3e12e722efc59ad6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ccf8e3d5d9092925068e23ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bae91ba4f2979bcdd13f9364;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h734c5fda4f1a3b47aaa848c21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha66c7af82a87a85ab9847069f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce33a604eec65660732c9c2f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefdf96f6c7f7084b19f4a17f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83a86a656575dbab6630e4761;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7942d65c38bc6b19a991f7412;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6a81ea4b5b22defd5cc3a3bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3997e26790fec46a3bba0d8f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65dbd446a2ddf52ff431a8b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10379c58e3cacfe7a6f1c01aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83788a1f6cc032b1fcb713b11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b986cb68c9ba0187335c13b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f33ef39dff5b1bb04dc3e8ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cb3aa4c7011ad06e1fac55d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h525c434fbd2bb6bb2c88b3d1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde9c9eeae2a2960777e2b816e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he533474b17a0c4d03e5e7c455;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e5b766792409a9bc222f7e49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he24d8f0c54dc6ed4ae5268945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd61891501980d3a80be020ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51c447b38ec0b4cef12bede79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c61273d0ebf54de000c44826;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d3af669f1d54b1f56293919d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8a71679faa75134f4ae39ded;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63aa22cd7c5097d8399a4cdc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2f073c7a77636bba22d539ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e3110fdd1f7bafebdc70e654;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habcbfb3ef05b5e946200ecb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30f9a7a8b549c4faa6cdd57ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7aba5c06de7190953665609b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc55aa2d974a7158810ee4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h476aa4cf5812e49335d36f07d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fa00f6ef11c8001639fe67ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h887dcea0b8764449f71aba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h438283e2e3a7556d82c449025;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d936ecdef78c336b4b579a4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf199727487e44837d3e0a076e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c9b6dd21d019663b60907e8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h559da9e6c637c7ac77e19ece4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6a30981abb23c700429a08d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e9fa89112c17bca2d2cc267c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69dd80e98aea63beca83cf514;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38732c8b4945330d6481f28f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecd10801eb1d09e82481ff02b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba73840fd329bc4f549abc4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e55a83079e4c01df69565733;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95e96e53a7c0320c5f8468205;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69dadde4f253d8875f9db8e6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h408a3203c712e04ff030f0ee1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9807b515ecfd925a2f57089da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b13b6d75e1705b572e7f04dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f3be4ae9cd19f90609bbdef7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he19973e76a10df19c2cb6941d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6785d8c8848dc5b6c4d607ab4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf043e5eab8dad977f3c315dcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15c4ce94cebd6ab3d74aa3780;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb352e21ec947b022b3d43c1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h549ab6e0977bf235a51c8649e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eb5b859642fded7c0d2ea161;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h630dea1149ed592274d65eb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha260976bf66c4d1cf535f7dea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h608b3e38900b564560b7355a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6087813241c317c34d9776b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f36adc4eb77ffc335f77541;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41fa87b911aeaf0ff074511b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96457cc168d050c65f71c92ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha834e39cb9c3177a242288b27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd56686832d41011974076a492;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e92f29a60fe83cc5e9cb999a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d6a618d21ec745058eec0d62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h863959daad2ab2e720f92224a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h865d6cd4df9fab88cfe05a17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a2282ab68408dba0c57395a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8682ff7c44bd3b008d5c39de9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h255f8adba01465ea591f94edb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47a640837bbcb9e6b729e6542;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9405012ebc06715be6402f9e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32d905fff47606fb1b3c60be9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h790b0acb55d0f71c6de67220a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h309bbee2473d87f343255cb89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfce3038ad5ab3145dcda6c352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4caacd8616cdad8d3563cb30e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7db37ec5c95d5d2bac744a6e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c4eed43f511c0c58e4c79d7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0a411c83b7d5d29144a1adf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14b81551d7a24dbdc2594e30a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62fb97defef18478656f25448;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c1d1c1e1a2a606f5f109111e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ae6cf71e068ad03c58b84aa4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6c8f5045b1e86dee72a7bc77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4319c36d475ab9960f0def84c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b45237188c866a6b6d5d2427;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd92ba8a11b8ab2f3abc8b0203;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e4cf81cd7c8b75f5d1f12012;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12c164e23e7e9d6fe5e80ca13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99d77b8fca29482f8802e8dc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10fc2fcc8e11686f6adf92740;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1cfb4408b68bc558a4857151;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha40a6ff941fa105f86457714e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32727fb7edc0fa48279461cf0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a7f31a9b0c3d37b5d5ffb0fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8eef76027ac4a95db48eddffb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba675c5f4111395d62d0811f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f4de227e36c2954dd2d4ecd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h933e5d8ba439a9dc092167dd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h225e4fa0bc2f41ff0fa7cc6ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcd655d733a433e2c744edee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16b1102b23eee514bef688b6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4904fb2b64a7df2663d87bb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7691f4636bfc83b81a4d0166f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h728c1ece1d20c0a0da5a8d1fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46d60eec5e2f5240f063d7af9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc16e069dac421f86dd48e425;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4dabb2b4d27f3f2fe388cff9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25e5222ee31c809e925fa6445;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9db6d8526fa155f05406d97e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b323f968cb0e6188acc653df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26cc0b6e3011a180d2cbc9827;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8bd97c23dcb354f8e859e096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41ed8663c121bb7c959e59a00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h724caf8ce115b285ae5372cc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf786d2e621ceae4b8291f06b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a93ee35b4c41ad6443b28979;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf48a8eb71cabb3fc9c1fa11f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfc3b8237c9e96c0bdca812ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habcf3761f2ad16462e46b3cd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h257c86b3347f68f4ab558bded;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dcec76b696d0f72f03871fd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7633bce55b531d8121feef91d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4838a6921d03aa241aecc5e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf350587cc58c4ee423bbe847d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4eacdb1b82b1a6f9748236f1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h253efff82bc2515b78be347c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75f40485a4a0c803c7683e511;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a7e0e900a46dd343f2942586;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h222a24d87c4c54f0352eb8512;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h164360ebfa98979de3ccfb794;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heae9b175e7d22e5d7a25f61bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd8f186afe423f6988462be8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bc0f69fd9e162dc355967847;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82e4228e101eac98b05d50e51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12e832e65dfc2797a74d7de04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc838bb83f1ccbdd1936e25ed5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd561ed364cd43a899c12c1d17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he22db6b876deb5ecd4c77824a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd723d511bde617da2e125cf0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81811b7c59a0ede042b6b6048;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb44c1946552bf63552e04791;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82f5eed7efd3436a879ae4a5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7962560c2886dd2c371620dca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12661b2a26daea153caf4dae4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa4618a5e57dbb382b31abdbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60a9be759c04cb21863b9ee34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dc2e8a0bac06b00c604bc26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0630f674ae0f3557a260cfbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a4a5db4fcb2a2b909c4654f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha886016ec8396d980cf66baf6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc33292f5942781a2bb67fe51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcf1f8e0500352282c96006bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbc59d2b627100449c086365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c8ee5c020b58f1c26be1a1c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28ffdd85d125c81c7429de1f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdbe2be70ba39043f496cebd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce723683b667a4ac1dc9b4361;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23721b295af596639b25c7d2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9182d410c2f1654c3d0b88f0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd552925f74a7253a7a017b7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4f83543dc134fea9ce71b3b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b7a2e3bd9b094bbad9eb04e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c41e1e7cd6b1fbcba493f08b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3d4c51c27b872b7c24fed29b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf7b8f9771a807b0b7c7baaf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9c1ad294c351b3c57bba98ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h988fa07a6ad1d586e1126e864;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4793d0b493114d0b2bc197d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95e23d35792eb76d1d4786c57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hacd7f43c5535cfe6951c1035;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc284cd0d0936929787090166;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f5d501b8bd16caacb171b558;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ab26651d8acea8699cf6c85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31be2214fbbda63155781dca3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4478e014a2a12beda5c9293ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d7a29ae2c22e14a5c62a11b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9739ce2db3ba83201d54a7178;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21d598ad5669a1b784a718042;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2785492b16bd68b600acfb087;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha910b811bf96353bcb5c24dbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd4484504f32008b737b8a6b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h829e93df8228858f21b5fd365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda6f494ec9e3bbc43e7d9a9e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eda6772920c0e284e7c68d72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38d47d663c798490471695e11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2ca62f0ecf5437d588f36cb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfefd87504f8486ec95813f037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a68d76c5280dc6eae32569a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b78e36f50522eff9db6b2de6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbece9bcda751859346e0e1a9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbdd566fe9bbd4837855629c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha75d5d35a586d61dacc0d8903;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c3ba12deb7e5bede16b0135b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57aa9d8e5b5ed52901c9938ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7b010ced62028e32a47bd133;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc9d2ef78d8468515c4d038de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92f7fc6c337f0f3356ad8235;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc28c1a5bc78ba036b4b068cc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafc7fb2ee98ac7862b6f8c399;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha75cd01a6e171b72ac2dca94c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21f288bed66dba794dd5edce4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70eeefc77a9cd8750a0da8eff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4500dc18a145b99f5cbb759ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f60e74e8f709f0408cfc3a4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfde99faced7d81f5cd7c13fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3e016d39bd0e6e362b7a73ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a6ebc8cc17e9bad85dcbefe8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a6aecbd3ebc7a8ca7dd4dd8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ae1e684d18d2053621e4525c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd27358c7add4987cd5ad40b75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1862b9ae6b71e365f3b9f454f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c576d73cf8797d9873d57ea7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h148af5144bfac72985001b4a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c58cb0908a727f43aaa7acdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a571e21d826daba8a446a64c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18ad37503ce37db5cbc007b8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cd4349e30df509f3fac5e6b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3b0907ffd5cfab99df30a4f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb902b05164855ffd92657a5db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dd9b776353b50da0dd68c7a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaed21ede0b78f6d6193e3f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29ac6168a5cbc043649404897;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6e63ed297d8f4471dde03f77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f8fad23bbb35304c40174111;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h158f0c69f9f8a456d40e9c99e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h679ea44fb632434fd0c28813f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h400722ac479b784964363f5db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4be6090b57546f5c0c4ae342;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h584980d657508de5a56a162c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82a09013fb5e010ec857afd20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc385a5fa3aa21fba9174a409c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d3ef4c291d224118dc0e98c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96072feda4297980747c0405;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee2999c60bc2c5bc08d264325;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78ab19900f868a4bec428f40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4f4621ac33d74b81d08d16ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12ffe126e8b6fb66f39de98d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1449f4d4d6dea866671c55da4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd591b44c694e801a48b0196a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd19be8f7aada33431f8483415;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93eadef120a62ae22d5c6874d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f0280a53c52b0ec6f88ecb53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94fb2a0dcdd21ac0c7a907bab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a75e6382ec655df04c0dad45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac53559cb36575c23f4ff9579;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaa9bb649cade96e8d42e0ef2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h109e7593f261ea993d18e2a33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf980c124edcf93e7eddf17d31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b1685d7af8735fcafac8ad72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h938b41f173533e7d6e7051730;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h818b6da9033b8ab66eee086c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa3cb10807e99b483b91c093;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5a73549565e23987ea808ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h596eab8e6c785415169a0a0dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1c6813c7d3d46d884832924c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddf3a79f64f2017e3e4839a3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62c2902ecfed7d76182109003;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc27121ca6f11ad8b06c149cc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6254c8e8734b5944f86f28124;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4299216ddaa5f3ac749ceb24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd160f07257eca5750e63c977b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3a29bce5a611a5998fa9271c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc78b6f4ccc9bcc9f73100681c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90d74715496804a83e6acf5ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha89a97b57bec8b38203c53aeb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b7c1803933a409ce6529e598;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94a44302d575562647954d7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h643ff180d8a2e4be09b59908;
        #1
        $finish();
    end
endmodule
