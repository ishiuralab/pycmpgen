module testbench();
    reg [17:0] src0;
    reg [17:0] src1;
    reg [17:0] src2;
    reg [17:0] src3;
    reg [17:0] src4;
    reg [17:0] src5;
    reg [17:0] src6;
    reg [17:0] src7;
    reg [17:0] src8;
    reg [17:0] src9;
    reg [17:0] src10;
    reg [17:0] src11;
    reg [17:0] src12;
    reg [17:0] src13;
    reg [17:0] src14;
    reg [17:0] src15;
    reg [17:0] src16;
    reg [17:0] src17;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98e0d5b486e6c9b05c216785b6416beb16ffe57b657f40a0d47a6470fea77496a9e01fda240d8ceae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc3116976d33d924db33a6de2a27e67f40bd7bcbafaa9e3bf64968a5f3b6b07e195ba47226dd3f05c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h294aaf6c521d7424782860b31a83d1bbb9fff6acabfe002fb4054532066ce2971a61af676fa81b8a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h404c9c9152bd0948fa75b06c6fe7e7eb8aff641c8e137914f774eddaf426d3ca3bf383dc2d9eaa06d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfa8d72c8491f882900e06447fc230260d021193015cee9c52bc7740e1842a86fe8ac4bd697fb07f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hface14abeacc0524164fe25015029b0a7f92210848f18a9543a7d42be8b02510afd98ecb4badd029;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2afc5b168f080b2ff700bc3e8600e674a6e794be15df073fea29723b838a98dc873de915637b3f285;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11188f858b2e11d42f5372ec0c3039a7143d0d64e57bf9aecf1b840815583740c9d5d353ad4777b7d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ebb3a03fc4591d64f82f4dfe7120f6d4cd3041258ab335ce08bf2338151ed3995c4ded10ac3490e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c1513b4ec7c9c6583ec6d83a00f08fc2fc8468b83eaa7c91d818f91daebf0f90229af67b85800a47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d7438f642bfe3ad0d8371947dabe7da680fac2201880a4edbee1c13ae3c4e58075ec995f5035332;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d5041de7055884b99a2648bb45586c9a627fe9fd83a727915824ac8e91adefbf411d731d5aec1ab1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a997a75cbcb50d44c1f995a98f9cdf5b8acbe13033a376c84fe6f16af7bdc49bf6c541ccf215db1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3bba29665bafa1c6232194ec7567715e047183fb0b8fde7e0de806e3276cc884f1b38c9d89ce36e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a02846b3c19b46f5f16298b051fa1718aab48a0999977c1a03d041491df0b8b470e3e5d6f9552676;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb77e40a44aa36e86ade202734a7f4b7e64a13ab7c2c1840e164879bf72cf5e3cc254d9ba39f27d04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he27f99d9cf4290bca24bc1b8a9f44a80b94109a967d96ed6ee056d44f4b63738a046cc4dbf7a04a5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27fafb6889e02e842f07a0ad8863fb6add237c3e52d9270b4b954608282fb9b3d146039cf04ff0366;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2505c75dd2accbc5c46030709c6cdd31ea8a7e676bbadc52908e02f4656e6022bf57b159a56ea3f18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b68517c9a2a314bea3dfa309a3a993b18da174dc1e9097f03f26571ac7088cdf33b787ad4eb15841;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9774ea6963304325d4d8d01df5ff4efb7297dc01372bdf31cfa163e07f078956c7d3bd8ce86fec67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe433dfa5fa578392d226495be0d2d3c236e9a07d302e51e850a6cb94944bc435cc61669140b7da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1119760229f20e25309a1d03e8d7f072a19526d86881c37c105076346c2178b7f5373a17062ffdab4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5ebf42d9c01db1902cfe9cab4e843bf9f2f3d3819f4607d358a108de72844783481b8fa5c0cf176f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34544a9a5b7d53e0378e2a7fc73ff3e3b0ae254480fe611529cc5ae933cf160b71bf43ce3d89fe2c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h754c01db0c42afd1d04d002b3c76067f2ae3df6b19e29e3c7710c759dc42e1368535f9b5beb1f8646;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd702eb50b4e3fd4ad2ae8d83e6b937db1abfb32a73e6814dffd115db877b020865fa058332964f07b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bca8965d0a0be7865b30cd15a0bd14b0650a265034fa37ef3503755922101b40e78e2aea9f15758c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5feaab55b7085102e4c0a8f5e3b982cb82ed8ff386df7a8310c2e04d15f2e621ff982b5822c70c076;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27bdd307473f2681ac58343bdf0b29332034cd05ce96190551a96218cf336407c90dd1072d6c9e8d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0d97b8a0707962bfb20b2a1251c66cf6ff8e703aa39dd8179f1b5a4471efb111c498b5a75a40615b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10d98bd10395891d6d50f203f296986c4b3fa00933b5fd5f48a18d69984b9ce10ffaaf050ae538c99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb25d33836401c94a58e0fda474b7e10b2f0d33ff305ceb1af25bf2aa24b7b85e170e66bef164a36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h211530550b426fb6bfbac7c67cb17f1585adb786801b1aa53b05745a205a3fdc4b0a48346cb75a85c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c2d5e2c012a0e02d1eead1a4745158ebce417cc89446e898b89836b5ef33780a04f99b12cd7fc859;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1349ca4858321e15f5acb0443119c41a9f38708feeb6647c9f9f8302b913800baf059500b6f15befa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57cd25f8387e28dd99e93a52492fd1eef3722a5107090b7d5cdd8a0c24889d1874d4729da642c6a64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a8bbd6dff4600d80f17d200eaf9b0ab65d5aae6f5623de41b927471b5bf94201a4da629d861b3683;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18c5e53c5f1e7e977e7daf9d7124116576639f29e7f76b935b813a9552ac1e8b52e4f60b9da7c67a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e89125479eb6a2064e3438c412ade91344cc5dbde6b4fa004f4903e4a67ebbb56d390027fc1aad5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec2f16305b47a55c45e9967639bec0ebe2f89a0a8b60b3c653cf3a0d656a86af35758371bf466556c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb19e02dbbaf24d0d5b83c5297722a6d6d3d21fa5d0d9bb1232138b1855e93abae6b7bdd0b27f16cca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c13d0e770309c80798449ba1a6a9784f5ba0e256d7a83be202438cbe29ca3f2b8c6371bdbbc7ae67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c78cfba289cdd253cf803adb85ec9c6bb15d18e2bb80d332aa9dee9dc543ece56ff8017f7b4b1659;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd57353229e782b1e086ce13468b81f496bd69acffac2a7af4be5dd43bc579276f5fa24efdd200301f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bc1e3fd06d12529dc46750435dfb765109a1a5e149dfa38ad58065b783f0a1eb6c3d782bfd7eab27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a615df5023062490a5f423f5c35d37e20233d4b36e6c0197e5f999010f88014e69f71d74ae1b7ad0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8f904b699d22af0f7708eb21e3b6e106cc8da34fb2fb43bdea420d758367eb8517ae6d5c38f68129;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76a7d95189524fff05b1afce0c292527f5fb8ece7e4d37785300a104171f0db08aa04a8f1089f4562;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf68f1e75feea050ea240273c52d841356abfbfc91eb6a9b5d81317ac3d8c0beebd13dc1d4e6caf512;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf628b05f05ab6dd5c5df112cf54120fd6e6263a4d127332845e360a7e2c4e8a3bf1eb84a3b56e6196;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3ae451d690d13354669294a4f268a4fc6608f01f7b9f4ac61edcdd95fb585f64a60b7b3d41b749ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb87e345e08207bca959e74e15bcc717f5736416b62b521292c81815d29113debad83d712d7dc87b0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeef5abb34bd61e75e93f50a42412e3fff9846982ef22de437edf2f98d7f6b6924897e1e1ac6b12d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he907a76b892d08b77b6352d67986e12a11ae516692c507c82228c3e113fa3c7dcd25414c7094c3a12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h393ac93a75f8afd21a597ec3f71e38369844c9a1d293a02e7ea3c527004d08ae97afff7b901cc6f54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbe0da3472c05269b27a48827e63618ce70a06d66cb469cdc1e63c9c61aa37fa4f8b129a92bcaf526;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'head82dec93d4210d6c98c91847324d9914587e6a9dbcb5ea5e5f0738a778180e39e181a69f296fbaf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c5d36bad2b8915a5ce0ef547c84a87d43c3cb6804337b73da55516e0b2636dc33f70a64378f18505;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39e5869447b34c3acfdefc7db73a906934833acfaedd2b3fc270e26f4900670fed5226da8bb8f4eeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aefac5c02cf0b8b8dff6c9f642d05a6455c4080d7bb8cbda70b42fa6fd76a54bde39ce6d995b2532;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20cb0aed52b4bcfff11c0398aa03fd4759bb7ac4d5d97261ddbf3e4f1fa6e12cf15d7fc8e97a943ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83aca36825ed974031ef05f83ef28160b06eb4148fc667552baa6d4cea95c72c7e6642a3a733151d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b3dc19667351bcbe885e70238ecb2ffaa710cfc1dfed8b80a7c26eef9c3e5223e3734ca212979071;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f2afca6a7981da4d7876989387759e12343a7ea4736646bad845f5b84bd1f934b27258de26ec0c39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4cb408731dbdb1724df839446d8085934128bf111e49d1d759992ba9665b71cdcd7ff5dc04e95934;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ed31ca802d33a42d4973e1ee11bc7b6d3bdf4fbdac46b8c6e8d80f14e0bdeb4d1fa78044e8f74b36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54a7cffdbdcbdb60ab1dd31e2ef5c489efff5d910c8f6d4cb6330cb3311a9dd549d4351ba1736ddae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1cf209adf0db9017f2d90d8abf2935ecab8647e31b5b64735ba8c5b8f76d9876d89b201a0e58c0ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfed5f71c0cccff94f7dcbae19850325a86f000ad8e1dc03d5ee8000140d808da80f22db2592251248;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44138e72b27f45c1dc0c0d4bdf09d164ee1212058697f9cfea3c96ebb97fcb75b70b2822efc375402;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb23e08608e7c884f11cdad945e7c01daa67bc025dca75caa57e798f63cb71322de327c46cd15cb6b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h848ce993f8f8993d369c47bfe0b18fe1971766d80762fbe841b51481b6e5fa48a4af218e13e5fd173;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h860cea9330e758fa986f971f3130b6bc96a8c88e1e3b76c892d95e7ec3b8a0423df95e09e9cf89670;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0854bb147b76bb867b797d3275a17757f12b35c375b0611bf0fd0b2cd208b83459de7c3ff2276dfe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34136b5c2a20fd8e49ee9978e98355f89c3d3478d65d44f2ed9fcd37c0418e0babc84cc767b11a1aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h626373e26b08d227d9d1bfeffb0a68b1de8ddec2d89cc63aeb3af84d97993dd7faa8878c6da5370d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha32cee11bb0d5a8396b3da98e4ec600abdc30d58f1cab9d130147fb7e24b25054e7ae69d74fa4ed8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7cfae449e68614c450c462c9bf89babb61579b58bb3d5e10bdd9e978cfff4730c99685c44ffa0447;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb572d7a9d6eeef8ba8fa1d4bb9c9f73065d269b68e9a53de729f33f3a1c8b210a3cc469d50b1e557;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heaf7553ad22e0d6a88f5cd78d35367c1e230c420ccf7b8ae9296f82c25ff5a777e44d31fde47736c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcca48e00399d25a06e69b260fce6c02d838e60fc80f814330c6d21bd80cd620fa9bbbee47757935be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6feab6cc9e7f1d0cee195901f0131d47a7f741531a84ed281a116dfa9013007703fea4971d1f357;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h536df2fb991ec3982000d6eee3f711f94a539a8e45909169b01fbd7dcf8c0bc6ece335e5608877873;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea57870c3cbd1ef3e919a30961ae4fcae5db7f14e70147b953eda098bb57f4f6a185d3042530fe27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3b70bee5ef9e79e07432dd6032f4db1f7e678882e1ca731f4b6eaadc9f9b68ce3907279573611e21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fb40b370ebab2c1a2714c34cae31e396c533df07ae4e21a3972c538895cc776c41b88bce8ae152b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h828af75aa06234993478532a15fe5b8b1391a000a39219093f9012e0c48139be3c41d1be6b012fd4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0636d5cc1e28d5af61cd8fb784e55a6a8557bedec6277959b8380d462f8d38e91b82e202b2745b62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6f1d2d407def2941d548780e8f787c7f6d2ed2064f9b98b30aa99094deabac74170609644f4c5fb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cb0ae678d2072dfb0a5f64cbdd1106c47815d19b772dfdc245b99300c7318c480db5ff0b11603cd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a0b611f20d1e411dacc2223d1dfccd0b8b96f0624ef30aecafd526b57e21707a647609c33755e6f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd75a1e569d29c4d312ec4099f4432c8da511027201cea8599d4f22b69120be23d71725c535d42b954;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd616e38be6286703524b592cdd59757bdbef73d729e81c17291d25aa275e7a80b36e914cb029a9e0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h824ca42ae1c5ef86e78e169d37052e3daa48802189610f272ded11726356eeab3f73eaea5c8404324;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefb385bc2d17d168a65a6eb0a326dece4fb6312620810069288d78d6b514f8811c725469b755c7b12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13c2d68bb9e0d705ebccd1c5cbd4d5d3a852634d4cadcd70e7f33050a9234b5f21d36835b01095b74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73ed82f1e998cbb297600fcb3902f08491cfdda505152a9960bc8630eeb43fc74458e8397fc169f79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3666ec0d5a16bfd53c41c8208a131449a7ecf9f79e866b9efc350c4fdd9d3b39bdb07805cb26b6922;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e6f15f129472f736345bd76e1d79ee6c9468b1bbd35562d1bb6f6f5cbb1c0fa8367087ccb2c772d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d1851e8e2e548da695f7b15ad69fafa4b5d42f870b582c60c4b1da4c5c7fcf2e5cb5726e7d0849c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38505e89352f46b2e42117cf4ba3192cb441b7b2e0ccc9af90f3ddbca8563d4b1e08ed402cae2708f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6640f66a0eb5fa226b72d7f25fc1f468b7831ab0188477f82985a7e21f8518c94dd04b245feaec1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34500be8eb2ed4eef827302e155c7b8efeffd8522e82aef3709144393ace7b96d4a0ed26f5aa2d2b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h883e8fa0f7398e0b0bda1b2fe3d8c48d697d073c426959b3bd3d8b0689a092cb0d6b86793f6ee4f04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h326f826c1a08e6a6bab3c08853306392a0c082e69797a30d16e351d1d5e3a9eddf445134b55464f5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h424fdc5798c70647c15fcf15c073ee3c8b89076bf602ff3c8952f52f3d663179466e5f57f2cbec334;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fe82c582d461cb6988fa9918e8641eeb10c3b2297eeb7a89712a9bfcc39bce03b3ee3a854e5cb7e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7996d79366831ae969e240109ab1947bc8c9c24a89d4db5f242583c34dcea213b60884f63c4e83193;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfef85b8bdb868453060747372e869334a5fe281bae92ecbe297544f3e2c6a7562d897bc9beb4b9b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb09258fae6c59d5653641b8ed148a32e4eecb36545078c75af41e4c22e88162d1b5991310e084dad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f55ea6db097dbfa9aa0d863a7f6315c86909a08a9647823bedd58b9270a2dd8ebcc2230fdee07ed5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6274440cfb2ee792de4233eedf9021b76bef4d40018adb541402daf389afa992fccb81932bf73a05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dd82bc8840fd0eae8a2c7dcaa34234811b44c1d55ae4c2e60e9e7d3197fba7f5805300db3f1c5047;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6596994eb669d6cf7da11fe8b9a3b38da47be88f04f0ac33d32f5366de796db6e936e725aa7b3b7e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf149618ac9995a23dbf2c9c0dbf9de9a0725156cacccdd4a95f66f94243d40740d3c3aae5a82d1af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7537358e49a4ef6a49cfbb594523319cff6d3bea46d4ee77a79e63d041051061aabf973812641d439;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84968bc34c33fbdd5af1c15df8a0b8fa560c5bc26fca2364b4b61cb1fc56c7cc2bdb64c86db01588d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f4eea8b454add2fce57d6cf01a726a1bacaaaaf3bc4b5a9ab226ad3d4441e7d3e293b357b090caf8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb49ee7ecbf3bfee33948f852fcd4c37f276626b273d97757caa7f64e3a4a721e0029ee8b0a169d392;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h810000cc4f0980b612e7b9932a604c995cae76e58298acb76a1b389ea47c2b9224067129b74878083;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h941cf9511db19a33ee826848e35ded5570c19553b41e4603eb0b31b045cbf2eea41d5f5d78ee06cfd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cdab003aec429686c82f8be79295d95a9fecd6cc3199285587b57d5ac560e2f30c6ef590e7e01b85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5516157a8dcff1c45db67ced9fba7b995cde519e7f7d314674c46fec0a9d8e9000edcca5c8ab25d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa3ac8f533670157907c8517fd03fb2056ceafd6347cd17711c4138c6f4864f9d28d0b0ebf9855a9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha043136140f4ded798aa1ace70ac01fa3eb38069fc8e8bfb337a8cd393e74d3c10d47fd5adb5fac5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2effefe98e3808eb2652c30a59e46dee05689a5ee90bb1d7637aff88f42dd3e657382b153253e162d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1b0ccdd22583a81aa4047658cc838ae6e8f0c05584432531790fac1ef07bfd23189d4c0a5f089ffd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3e35020bceee4ed1548fd85a04a787d234d3233f16c2291cc2d6218ba7153618880dfe3b96928369;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93317f8c784a1f2bd6992661082942f885f3d5d18114ba7ed44231d7ab6ef4f1cc2938c3546b8b920;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcac25f153fa4886247b01656b3a21745d0ce37bc6a4bca08a05f4389adff7b973798cb0d3d402cd92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf1552ce2be3db12d90cf2d519da1561ada2855acd27b1a8aade32d283414feaf67c673c4fd45924c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d1ee69cfcad2eff0223012b6f4f3f08b11b6390ca6ee7097e17772d6dd34cbc4eec4d19411c7b096;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79edd47b870aea547f09fbab9e25b4239518787e9fbc38557b7b1801363dbcbf0ca393cf5e020c262;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82dcb19678e5103bfe18997f5ac42bc5d40f2749522a07d3a3e14cc4975dffcc8c462e52ff9f25446;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf01b19c90477276a43702638ead18e50dc65e7f4945adb9b34a00a3158dd07167dcb517184c03c4e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1f249c8536012d7e8a89c747f3dca84ff782b978773b27c5061c20421f923de268c000c4649a40b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e24d4ed8f12ebcd416c46c3aef3c75f6ae661beb2cb6fd4f2d9399fd3207655b26d7d075f3d54fb6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8dfc305de00b7ada93db633c2ffae0becf1392277262bb2eadc0f23cf8d67f83760a609933e8e003;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h354e0a85ee27963a7e152cd4f80269899438f0f149872fb57c4f562616ee925cde58cc7a36f6c364;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h978fe4605eda2a0c42b4eb4d0c3a69c4de4f641817fe235b5ac71ebf520629ddedde4964d8ee11641;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b5c04ca06d39f78c9d00382990868e8e745a894a635b9ee797a6003aea5b97c668c0aa7333fea6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39e0b791841f3b543da54b7d5a52562a543cf7e0ad1b1ff563527f3173737aa8c08345d98aa319a42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50cf20c12c1ce05510783ff4d92fccaf9c1f5b1886fb0f4aeacb5eda35554deb78a3ac5929c763d86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1c1402ae7a8ae98b0774784638ce2f0e878a07b58dca39962b09c980144af35c03362f26e57510ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63f430b5b89966206472877bd5f0ccf9abeb438e664e57a0b86595671e9ac80d6bf018afad4200206;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5561394836fd93f9c7b05cc3f87b7cbda540d744d302b75c1cce6f4bd2f0091392154ebc6b98c320;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7521ac8a14e260266fbc2b6dcb861a094c4555d2780271f376e2f8b67352db50bd23a1e73578a6797;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3833f4c342aa566ecadd96fb0cffc914a7033c36e77e728fe24add38c39bee9038c11c7cce3408bc3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32efc70d4f1607767fab33f97e539017325904bd60079d14d8d5a7b46b9dad7be2d87511362206a94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38c32e4f3fd8ac437e90ea35ce479601ca584683a4186c4d7c8ec1def3e15ecf366a200447ea233be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h597e691eb7f6dd28f99fedc01a707982d5adb930198cd503fb5ab1c55fd63926fe2166765b8912c16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h578203e8e02384f37c1bb2beeb477257b246d5e511e54d1f94f5e009c575fa07582fdf84ff18b0cd7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc75181187decf2ebf413ea1ac13c7f1bcd0f4657fe70225ea50aa3f5e7da2677d173f649f43b7000;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e931102953805b5a4321b0cc3aa44e6fa3eef85961bd27d1caa03ae2585d4751b37f8742a9c6c3b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd08057406f0e0f93c1f508aabb989637a3894d283766f4013e922913769a019af89e983ab64edfdf2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4d775852ac858e48ad5a70e8404ac5fea910f58480ad3f5d85d7f44ad326a5de831328478e92747e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5679ef31d9d99d8b2607254c2012145110b7735be0359d139405d104f2f619cca8b2515fbc34eaeaa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18e258f22f6c5038513abbb672d8f390bedce93abec17fb26ba79ba7c8c5a789e6e32253326d2730b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1298ce2e8a3b6fb70f980cf554283ce0ea60c589f6f92ab2b3510fb77ef0a94b91404f50ecc5ae3d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h392dc028c6f8173efc979e4dea4539509c6f322828337d1e6692ee4935dacd0d860b2133d361890b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2de0fa5d07469dd05bb9d1c19760ba92ebc938de8087b4748effd8eb8a4b7f887069c3018a63b4901;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a255e6eff73f64e8a9b09dd8e7048856160191f0faf1bf303ac45ed5ad3d63209faac7d93f9696c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17a9a4d447f255fc4acbf0185caadee3cb0ea74940089c58f4aa9df86807003d491f318e8065405f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bf0ceda04751fe958ee30a10225cd60746ead81448f316235499a4afafd11c539dc08e0b975c33be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1dde4e727f4c31d27d404d9b50b3c96aba93693c34b684aa3f09521d7c4deca2bb639fc1d75bb192;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64577037daee1694d3201ead1c46c31a161a1bd5b351927ec4d133b31e3cc744a0aaaa299c6416d3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14b7ae7a4bb603fab076e5ea6f19b7f6389f93b67b9e9d0e452fcbc7b07dadeacea473bc857112fb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h882207b60d59033bedb64633a88780f0da765b7226b0765bf6b4530f7f3034d931d47d2d62c65d61a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h778a5a964ae436ecf76a2645f54fa92363d7b57a54c98d45e9d09c9ce9d65540fa99efa3dc43cb3e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h340c4753325fb428664e9aed6aea5c8f2d8b65668b553635ac0a23e84da760ccdfcdeace6324c4223;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1977718a71af99a500147496d3f8fb642f1f2568d3c2c111c9711039ed166636efaaf6da861c1e4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefbb930efa6a13eb1e98baea5a87dd6f887293d4ce1946d204707819d28a47f9b0851985d39db98b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6f56a371514b776772aadc685ee7504f9359a6365867cbc6480fe20f39b8bddefbda5233b7e28f4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd30706f227e1e8f5fc1bf229096f0c66aad9bd8aff5225d3eaba658fd4dbfa99d3b079790076c6fe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3196a55869a9246bc9489b435d9201cd5af75a8a757ea45c6901f4c051e59fa84bdbd6b43b4b622b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfab8697845f61e39f560803fbe6882be9b2ad6a65cb5345ebf6b0d95f82025b79970539ab7505b9d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c6bcabdd180eaa3139612b69c1afc109550fad52c67d27e8cd39bc5bfcbde53c3148af1d6a8570c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cdbe7ab3c9511e7b0dc3ffe1c8c674eb46a5f3570513cad3f921bd68591cb78591a129d1190ef373;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ad9bbbf55ce5ff8868c8498482386a3022c05fd2f24cc9cf88d3743424ceb34ecfb1695e5d09f665;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d526b958cc806b35b8325ffa4d7ad563f6c401df5d847ebbf094bf0f48821d4f2932169d15e40a6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91b6d6b9c2cd201b96acb4961ee9d447c1873e69d8bdfaa107decbd3ee452e670f6e6cb6eed21d460;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8c8f4ff849745563780459f00f5f3c36e9ea5d25967e56972fd1d96090df5d51ed25376ea9b5fb72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5e363e7176941e761088eed44bd3f3ebc55778873d53497a42c9c9630ac9cd5a2d55ad4ab0df7e24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6797dab5ca494d6269a29b82b7e7ab4617fa740411604af822f1cc26feadc173f133084d75a80cb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f6e073b870fc4794f828bcda3e735f75e318f027e0bb48883d2a28cf5ea332a5baf97357a602ca18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h570264d20325f3d4d7ebfd6f414981d0e5485da1c2c594cc1f27f9a7c5f332f9c6fc7333af8a903a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f3fcf179fd8520048dd008bb1f84d663f6ae504893f04c0e83f998a68a4ee40f3d6c0d054e7bd130;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h668cab2bf92fd4cd8d17dbc78c8a338e63d1c79bd0814cbc2ea5cf18575cef7f912c74c7efeebfce6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62a4c13b2af2eb8bf523b0da4bfc39aaec7a6e7184186dda90cd72543371c0319a169a30591718f55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6223b0860c0850c99823f89a71cb4d55231c36ebf5c0f13a55f00c3d8b8cccfa9b9ffd5c3137160a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h725b4ccaeedfff629975e3c6b1d4134a5a68a55eb66376cbdb21eea4235316161a3f1d79d5d5198c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h798c7c7da7a44d560202be98a2370dfea5a8978be9b6f38408416ffe75b52b2214119043d668ce886;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dfbad37b03a92a7b74fce347518ba10b2a406d97e811ef20f3c530cf9b189813e004ea7b8d0a4dd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habe822ffc66ef8acd9bd0c9e2d3f2e8bcff3db7ff87da0eab68fa305b2e512c5ca8441e4d9d5b28df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d7213fdc6d3e276ea7fe1c3142bfab9d043a075ed2d2baff3651ac8bbe3883437ad093db75f59fac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d0e6919ec06991414799093d76357489c786a61d8875d2e02b35d8d109c196b215f140d8b3a86c53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2de141a12dd21b9548a84e813007002b99978af003eb4a0e152961fd0013c7e7a954284dc144c03b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5ce1c2a5df456dc654cf920dbd516f73f3668e9d5381bb81590ab61da84fb803e1e9faf9371d798;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h267cb74fa63f502117e5a8bedf6f41a7fc533f7024943f2cb47659766ce5570af8811a2d98cda1c73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc3075539e21b496821163e4caaed4453cc3ee42dee19848eb34410846be1c6fbbf57e992d16cc220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd99a79f07e9aca1c50fac7fd3ba5ced3c4c61c038c5d399ad9d0dd9976b33e6ff9864d3aaad447ebf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ed5b7e5a3024a09a2e2cc1b28cec1f0220136ddcebd72b795e548b814fd7fe7b273e8cf6f3d3f2eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b779bee3141b72a639ddd7f2bca5066ee8aa825151740ac066529fee19a376467b0131b3f8e61b4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b5372e1590c241327c0dac3be2645b85cbf21552cb366a58475f1cf497711530d29dfb3989b6db6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4becb8c2401de5f7a784a7e3102f019443a267882c081fc44b60c95ef5df3ca873a7c30b9106edff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a07da302932b9a9325773963f1709b07a9da044ac125b69a7807123c857d9aad122161f9b7aac860;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h340cf2d7e7bb9515270666055323b61ed55cff0a32b90b35da1458c799cae0ff6f899ff7ab0b4f83c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he284f4d61ff0e4feaea5f675f3f8068884be61db990ba3788be312bc557ec7c672f12ca3d40e7b0cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f47bd7af6b6e677ee751a572e6e660df4390cd056611ee4ca59bb3b0f1660e3aa9f0dd0d5089e352;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3e70e77065f92b768f6e7dc54ebea214926d5349b4d158dcd0102a6d0442519ca200daeb67357b76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf815e3f7d29f52003897a5e38a514b87c950c8eff86a39cfe2a64adfd849afb063253eeecfc419304;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8ac5ac8ddbd575e83545c0b52974d406370d426146feeb35c1eb965fdc1b9258dcb86a73975344bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h581c703c4e29e1f640080eefb58b9fbc0615d3535ae163c7cfb50a498c494af23d6b61f0329f67a1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94b1ca6c5daa70b0e8fdc2bd5d01c5f6569d0d46cd4b0152eefaf753d49743c7a0f61266cc2059c0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8614d8d97d0601157892a99a36107983ecac0e15da9a44ea2b4ae0f9e69a6e5324dc2d8eb8a9c368a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc44513ba15d4ebe017851ef40aa5727ab5d253a592d02420bb959a992859c3704f11192894b8b160a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h232ccd55d2021ca71d33d17414c238d4b31e4fa92413474de1f1f4b53ab1317cae7a1419099fb233c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha482fd1ded6db242745ac5bb4b974b98f3276f788c6a83aee7c4a38acb635c0ad57f165acdd356b7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32c75410f4ffc6e9c6bbf684e606408a783af029a60ffc3f74b63291463650bc55db0063516db7e32;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90bdb0b68cf8ea5c9051e5b0ec63aa33cc7bf2bb9c065778aff234f1e698329a5db412d3e083d2dbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2b50444c039b2f470d25c0fe2f0b3000f7e07d9e8a9dc5d732788c9ed0eacaaa94cc89266e46d16c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec2943603eb749a20331e775865ddb7a23591e1f1933049374c0178c65929943b4873265e25056644;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dc0dbb5ff58e260b62a94218f67188b4ff3a580f573dbc82e2e88502e4f93fc6e644e4b0f443943e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ed78463dfda99541befbc3dd989df312ae3d8e7874b62da981848763643f29bad18e082eaaf8eea8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc115a4a87f6f4c1b7b0a6a9e7df23b4934f0b440b158a4181334e831ec268303d0e6ecf1f2fd3b1ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6e5b65aba6c4859075c236407c9f1c952682585d94021ea8c5e0a50dd3ea6bb259b79085425e61e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf813dc425a1e94a4fdcfab856c2fed288a6a5357b07c502caa72384fae50de09bedb9fbda8603435;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcb9403a60206cdc933b948113d5ee0407e3beb354129e46df724eb350568c9428048a75046251ea7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2de4b913d1b1a77a166d9757d03505815800b8db79e869282567e760b6c32ae42073283558dcff70;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac11603e60e508f0b61713eb091d0aac6d862a9a691d2fe5f7d9df85ac5dc800e8da77b4f7f4c3858;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9086b102c95fb553fe85d3193db326fc0b8ca768b41be89da829e28b7ec84a0f12f67d5b7087b518;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41354227c5b6b1eaf812008f8b90bba6b5595d597f9500e69c2385c7f5bec0d396496c5c8a0809859;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h338867ce925cfcfe3fac95090f87f0f7b709a2a1a3632728c17ce07bb55550347a1d93527eb5f32e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85f53288cb8ee62023b31265d0112bac0879bd83d3aadfeaf94403f743db59d287150618be8e344dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78ec46e0518bb0475fb56542983e218aa734ed83b48d1eca7590ea5464500617efd124d86a158ca13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf451c4f02323d96327355a2ce94f5df01ac32dfffec5730a9af3d5a40d5e58a53934c96535952ba4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642f7f8b0f922a7b99801ef8153f999ee6ce27870242a634ab7d719c97311e13b17654b8c087ac84c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b2b01e99189b94a0ba057b9934881559cf7e968c9bab2c767ea9acefa6062e373ff346ef2c552944;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa869b3e0fe74abbc074360419469d8042998b815d9af09295f374ce02cd31890c524fd12530e1f6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31f6a2d6939076ab0ee3f1c74e29d4a86e7039814629bf8ccda0ac0d873a13811f9e45df9dcfa810c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c9b812ca1d1a267fa56128a57771b76d16c73fc1ccf7fc8319f09674d9c737b4588e47ac3c75828a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e09168494e68a45c5c8d3634ea55ed813bba72c6f444373e128c20825bc83aa3a7438a2edf48176e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd76098b042b066b6ca3b2a594d43ce2c902ec8401a187073f77b9e582c7fba3cc65750579ae07f920;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h715fc26ceaf469b03df05adc270eb52c165cbccdc86f223ced9d4246ae30ecb8e4945d178a29a8250;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c12802ec4ae8601640f17f83870c05fcdb5eccb5e6a4bd3ba9e29427308b1c03ef2d7ed16b90911d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ba1edc3d228da791a16d9f32ea46145925a9110b25437704a22f1f81e1055104c93b767cfc842645;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a874d4ca5acfa2db411219a37aac6dc5ad9507de8f7fb8c9c4ec576d74db4032725d012adb32ac37;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcee9a83f147bb50798300d294525965ba0c54e51355c01014ba4de3ea280179482d0b4844ed69383;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4ff738fe1294e08769915d72593a6450e27fb4f0588771d88e8ebfca6d4e09bca26ed470d085610b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec7a0ac2de76c9531f3c33d8ed59c1767a53a85ce27c09ea98b3dce7cc543796318a8de4d45d441f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h732881a0cf24e0a62c369e0c26e0ac526d531725dcb0f0d8d64fcd0fe08ef79c13ebaedf3e10877d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f5afbee9cfae8f1c0638ebf5fa5e60ebefc40759804e2b8ab83b6c3db7c92ec2e3ae08ae6c0267f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fe5cd7f7a86e3ec7a7939286e0dc1c87d2e626a0b0ed3f91125f44053d2e271b2fb2af620fa4ba2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf26017078dac25bd7306b10ad17be2bf3057bd28953d453090f4bab54dba776353e71d53743978e18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a51bf4d60803d635cd468b227f6ebd32366d16cd7f88044d21089630feabce13b5b89c6275c6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae01b87e57225c7a233f96c2d7f1b1347a1bc55d68ac724def37bc460604e5680dc903bf756ccada5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d50cee9b06a45f981074396af7574fb6d5a442514b4a4d16fca61e6af98652d1d5056e452b209a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19f857d66852e9eb3ffb5abcf44dd3a8914b1bfb74776017d70dac3fe1b68c0ce02c8647dc4b617bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb653793e5e08899b0bebaf446b2f427905902356d3047f2e9e26e46653a17ae32962d7cde4e1676c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee2200c740ad71da6ad57755d6f544f70f8124d2314a3215f94e6944178300ac662f5e3febf77c470;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79b4dd6d03f82a08ed50a52e4d2b4dbf1e367b12099092fb1d247aeadb2dc859e56e9b0a262335bd3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a62b90386ee4bb15365588dd1f042d9f3803338d7aa7a4deddbeaf4ba16630e8bf98b7025cfbb266;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h615742c6a4a087568fa6ee9a9f4b277f349c0f23e37d1c3a8bacfeb177cb1f7f8e20a3b76bf6707b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62e42d9d796557da7c2ddd9211615e2fd254d66619edd9673a2bd0958c5b0d0d7365f4b0baed666cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h936c7b01c27a6d72ef5e14af9ee84bff8f866bb46131a33f2bed9e954a876bb56655f199dd8c2394f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb8b9ff0610bc51f5d3a15fbed28566db727231413420829a63f3fa7ee4295954e6645f23bbbe7e97;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18ea912eaedc47b1c844ff2e62249f11895ff2654360ea472ca01a2f287acc83edc67c360a824c252;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96d2a5de18ae0443eebf3fd571faf4b35d96d81adedc9e539ba3cb552db9dad98c5d43033033fe4c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1569276e68e5f8e05a39417eb5b33ec79b20bc607ed2a7a730ffe3e39db3a807d25cf2ba28598bee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ac1e3b761a3225b0ffbf351b43dcf1f260678e1430d287135cae6a4684bc9b98219ed905b9bf309b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7d978059cdc0c4ada8d7789834674fe726c7381f6e91b3af4e78ca8d87e8a0cd20fcbc5f5e19475c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b3354d904bfa8db99758826f581a50ac08912933b54428a95c4a35e33b0991a31afa432a043d4505;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf75e4558a8bdb0be0a10518621845d933a834afdbd003ffc81cfe23d4e9ff991c5a8203e8c7fec35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha05d4729c15436489b2548f2a065239d58b2187e8993be56642db321de23d58cbf235f24d91a9ea74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86de06c393ab4f7083bc44b7bcf8a0f57f8e5bf4e4854b6685a88b1eb99b41a4d709b8502f1668c4f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86e047a4a15c3fe728028dad6d0361d0e3ae0569baf78a1dd7a3233ab7483fbe9db440e3554654b06;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f03a281a0fb5e1560cc5b2c5fb02c4f7d804b0563eddf30b322948baa760a2411f92d9707c0e9fb6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7f9706ff674ce1f1d974a15393bca9230d34204edb6dda34e59d3dcf6b292ae5557c2994b157b675;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c4def4e2f69bd4ec5db38b00658c6a02a1c40dfa8894907a936edbebaccd5751c8299806ab7754c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3110d6a095c549ab59972a2e566f54a2cbb858c7a967a58dffdc623b5fb27aa69fa681a0afd1d4f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h835c288f20d902b0e34c2784dd6e6c29a3ae6fad4fef167b6572a5297bdc1d628578a3475e971f042;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc264c4309a1d4b019e387522d349c42ebda298058fc85482e1353ebe79682d1a54db204d8bb76621;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fde0b94429ecf336a8ea0ec39500905c6dde093e6591c1e089184ae3c0f4ef71f525c137c5701738;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7545c16bc6d6f49cafc3cf103ae2427c60407c95cd5043a567b4f46d601349d8595b056ec448577ab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4bac62d6956d366b043b52978279e31b3798ada82b084b2d32ebd0a2417eb24a22bed44e707501d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5da4631d7d5c12a6c2eabce0761d2939d14083a83c484bcf6c7a6b50021f9050002609a25d6f51431;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbbd22dd0d9b48ec9f716660ac8be327804f7fbebf6e1ed68903509f7f863c2bfc595a4205d219fd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3a01768eaae9c3f8a51580e2c1731a304223f5fc33e507acfb4944e3e653d681b1e72a4582ca4b6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10fd2ee43a53cfcb747543e68cd1f4364918c67fea46c3f3f5640f788449dbf5e761241a194a942;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a0f8a2220a09357e078439910c8aa7c9c8dc94980ef210fab8b9057b5a7e470a5e413fb189608956;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45daa3cc5ddba0d6c820c460a945f2376418441a8cffe46e51d6d2839704aca7534364de2c19580a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc61550535cfb1a55b0f45a2e152c602c7273921f0b0766c4fc48a8172ac1cb4a749e47c5f911d21fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ade4de181deeb18645b4219f5a0f80186182210e0d942030ff9c6ecf2d4009c0ee1afe9cf700d1af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf417fbc2447f39e5e311d1f2114df28ed23f84b9c49c4915a69157431faf29d86447e1172bc7cba3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d5f99521867127fd1ca0fcebbd603e5209e3c19cec41c8a9f94c4b72c7293b35bcd517729c9d7544;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacefb040baa0dff05a56ef700e48054986fb244eebb8617a159db5c446f47ea78db0ade12eedee50b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9dfa3f3ad7f62e1664f2dcde5245a4a83e16de90e1550e1c681fbeffde901215885c3f00aab07a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1c1259c13294efffb95a6a97af0b226c075d23d87157a44e9286db1a4385452282f0a71dd0043222;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf54721ef1a14679abc44470b80a6ac5a20c2bc2ca721ec2efa4b5b28ef49d0f788483ddb9d5c994f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29af651bd0eba778b4b1b04cd61623508f52862cab02ab6cb8410ecf0e7115cd56427e551896d9184;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7879eea96f59e4976f54871d183c10dbe753d6febb6a1e8e401f00e969fc9c3f9cc2f0548d8e80e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h179c1e27ff79e0e2c8cccab9a8a5062a42cb535cc4d8315798c74d23ba2ae7569e36404e6b7df9725;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94b9327a7a338981a1477ea5c9d9f7e185259458f8ef02f64931db67b3e1c1950eac15063bc859435;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaa6eb749fef1d7c8981815979dcd8bd4cad0793e78a99929041f2fe0149e77076329989bb1afe9f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d1a1a1c4ce03f0ed4a56acd0c869704d7efb7aa43aeb62e1f0d7c0ecca9a4fb0d7b153b171e0be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47c513297a842ff4ab64982261e17ce7730073e954eb3a41bfd44634b874f37cbe9cf3399f06e52b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1a889da82ab7bb70e213ce7079b8cc58c152d57bd1cbb05c135db1d04781361181693e7bff93b388;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e424743fb5c31a8ba6ba28858760ab6bebed28748424cc51aa7d7851653d07117bc5c432ce7e8ce5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ca43a86357abbc78630659c83393c1ed978092d8fc5bdb0e1062f74af9c08448c9545ac0bb4eebd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fdce3c1820aaeb9f885deef10bf81d6b2a4b233e5b5b9ed03da0093f88f9f65715f187ca8f345120;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfacca0a960e8bf9bac8995f57e53426854fb4ffba45f0bdf6e25df5e902cf326d1b57603101e157fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec81db4faa05b5437b49c663352fd069bbf351f6daa74c50d8af553f99586467efff69170839f6984;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc45ee28c02e425c44774041ef45f0a80fd7bc4e8aed79c21bbe080cbd543b488a6504ad69ef19fbbd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1403b1bb704aeae55822cd679f7d04eb9d85afd8c75d6696eca970f4d9d97ed3c741463136afa3ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6733322650e1e010bb646c2073d989dff13fc23c99b5615c86bf12a25d5c6bbfe8155db8b29e61888;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c0a27f18c822475274c0cb57997eb75eaded4cf8a2135d9341719c6dd2f10a0760a00c6084b16605;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3633423942edbd2dd20a9df75c524d4167a93824cc2c843c1f119f6b831da24fbe31dfd1e0bf5008f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4ca844e30e34c403c206d97e195232f5de8328243cd8329b4ec644ab55a2bd3ba4993a71956ceae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc316e4750af858996f27d23ceefe753880a18d87b19059c64585d826f601e9fbb013038aabb7c47ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ddfa5fe25ff98691b34d3ea338fe46adda2371967cdbaa429b821e3a048dd7f4af2001b024eaf389;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92c85c3f75e98c9cccfa84eda3d2d71ea04f9d3d7aedd29d10c7d5cbfe9f687aef8c2d19a3b110284;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h811266133d0787c16e741d09e4c61e859c5603af0c05b1876001d8fffe58d6c998f664cbe04bf9c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcae31be5c1fa28ab6bcd83815013c43f17bc79afc90becb793fadb54fed3ee6e615a8a5b4f53c637c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86c61d2696ced1f3d02727c7ef3fa4caac830340314fe28f3808fac2fd0f6ba6a9487f23cffebefea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedcf06b05fa80c35722e40201bf628b162985f79c9e93c0a686829389cc5227f4781ba1d0c5da82cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96e8d69b9e2185830c347677840def6983f794b1120a2336d7319f48ef64fed50500624e5f903f9b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b10037d720cf79dab0fff9d7673834b5cc24ebb2928997c379d367954b6680d3705c74eb3bdbe674;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h784c4612ea1fe829fd8ab460f86508c24f88665db47e1ce1fa6c86363a60ed557cd1231680ac1abde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h175f8226e53c538fe98661cfe0ee1f81e08493da917ed6cb7abbda66e2c331e05718c6c61dc00b2a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbc6f11477561acc58b4bf520d1c850dc90cf8746b2c23f39457075ebd30e1556a2c4ed573d777001;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haec21703add31e084f202d585485f0d01380911b61a686604898b868670af943c0cf957429a165674;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeaed683efdbbdd1a50b896314a1e64463e3ebee479d7147feef92c07d74804dc1d754425c6545767;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb43bc9719d78b02b8bca7d5d2f0c9909d24d84987ffc3b75664ee0950d0ed22b9c8a30d5e850cb69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19da3feb5114ada225cda42e437c4edcd872b03e32be051dd85ba5b4e072fa88bbee528e73a43a3c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c4eef9474d36989c2c10bc7464df383fbd7a6edbe0aad378b1197f039444b43136ff853b82c7c891;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47c2193cbfff5f176f89d6167c0801027a47c7eabe2ef11f7674b590b0bf69b10500b9fd0cf026191;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae735fa847d16283424910fd8a2da338e73952948a08440664772410f2d136dddb6f379cef3707dd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffb4aeac0b305d2e0e0e82335663de2db76c3cba346b2401a860da896c00a0d9dab4c26c59f12b0a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914ae8cc741a6631fe938fe29c5b9839912e9bd805133c75dbfe1b7d0945b543db0344036915b44e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c14e47fd3d89b55c5f777b9a972fdd5c2ceaa388b32454d499e6eefe134a19f5ce51f1197666602;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c1df9e22b280ec0741be21385d971794e9ca7ff38849dc64f0521eebf3d5b0d4784856ec1201468a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d44f3923cd4f279c43e702c6c3fbf54a5bad361c14fc7e0e8bb2bd1820dc09ed6ae5ae46ba52ca97;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb89b60a2b8c9d727f034671f00b9d038f8e276b3a062a5cf88336a73c181308d8f68557f3cf277fd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71ffa591cc855e88590b0c5b821633c3aa3a02f0bf07aa1774814f214f72c88acbf1668f5be4bb236;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h976f63c648899881bdbbfd8431921663c0fff9b9e66bacc952b686b3c8bc6f6c9a0af2d5c8da29091;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he23fb9d3b5dae954ac6c1dfa08f6e54df433d1325db343b95683a8e8d2160e3d9308950ad708fcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfab3f850d06681a14b838410ad40bac33521102c620da37a2cecada9430e79f53453fa75c9e6ae89a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf674e4449c9098aaaa1a2255af9b58c6a4e6bf76dc243c273f93d3e92ffdbda77ee742f8f78c109b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66fc13c1802a4d03961f8bfec4f84501da575d3121843124e10f70d7f676ace93d86e012a79b2e365;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ab22ebf0381fe8268d5c52cdd2c71ed61931fab86c580a6a6a780e3d22a5fccd73ad5701316ed48a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23d6d2fb8abcf1419ae01eed53cd9ebe0fbd046be36905acd4e59d5bf4a3ff9f3b596525c668e6cd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c61d55aaa9aef0fcb37a0491dd4ca2d949b486d3b2216b5e897bb6bd74edb96dd431b4b6426c5a12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec7148cd3e095b18d7b6fd41a2a5d68a1aa9fea749c7175c45800c6984e32b9a200eaef845fe594ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d314509c9061f9a2c8620c324ea652b8e78b261f6adb91b30a6d71b3a0ee069249942f16e78f66f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c87588b1edb8899494bdd623a8fc344959d269ca79217c13e1ebaefc77a47f414a3173703cf1bcb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff9c7e48be71b4f6f7940322ab2287b9872af7f620c275a3e0915643f679adec3973bba0bd3eb8590;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91cbe41959e00d01650938a5998f84954ad6dc0bf4684a4b9b7497ab994435aa2c8f8445021ee7883;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h283d5536fa0d676c50e74892569d20a48ca6907d917fc19097c849de47d07b235cef2d719b64d4798;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca7b8583516e210cfdcc653f407e4e5c3d77f59b75731e93bb5f3106818de9e20d0295be531e96bee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee5c80a3010a8204ffb3ad966160f0c15cc238301bdd50c7241d267cfaef1b2b560169b49662abd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha35b9e6b29a839312fe21457fa920db67e5b45561d99ea84ac5b48a09ee0b8ae588e5e1103a28167e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc19ab66a89f41b4d87f4e2c3fbbad761e7c5af94cb87e4ad2d825f3ec8e1c9af366f88aa0f6accd0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56c423b3b5f72b34b3046854d1166abef87e360214978aea57e63964a5360cb6002847f68d367a250;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43697071200681d546c394a4157b48a0a269a42b05535bbab343debeca74a186226eb59b4ac06a6b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd8971e3d4c00ba4f30224978ef3b413984b43d9ed4c845752aa3da3fae390553d2e3ae2862c95a14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bd86f53b6cd8af114c2ad5fea0284ccf5ccd0e55c1ce06dee4c4a0f83df3b1d68acc43311b00c493;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a1ac97683f39477fc4ff5e66805a011ef4739abc96149ad74c71bfca5b1cd85d1fc93fe4adff4b62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a50d762252391b794c5a6cd51b97c98945e01fda8c157de63c077a8a89aae62c7ee2e25a3cc11a1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7c1e1653e7cd456536b6499176023d27c81689db76b49ccdbc1e96afd91a9d808f65e46400cc6242;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa40857b3dc25bb8e83886590e0121ecfba2dab6baadc4fd0c2d71b3f94e664a84fd7cb48e857b17a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3585c85a4b091046d508691ea28cb58488e2bc6f409bd43e88aa6567d7c3237eb3449c8e8c2e7fdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb597a356c4f1bf4e8516c6de0e67ffb852f2c009ab3bd99cf5b5cb7e6b4a6ede26be6ff753c5e6f80;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14f6e569aef2977ea3493629b59b5638dc61bf9dca176a1fd30c43f879664484635e4f7f328df86d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a88d55ce47e942ff3915bb2f548251a343c496d3e6a7a4dd078698b0a7f5d6f1f299c042727c5bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61b4125a06a96bf8d5d0ba1ae3c93d3d582b57cde183bd2e605cb10a5c143c4166d6978f7e9cb961e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2fd2e0baf9b3d62ad19c98446c2b3a9275a5a6d249cae1bfbc0b4681252deda26841daea55f672c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf065cc491e8c4ea49a44d998d682142f3a2e12d9d4caea575cb78e5cc728d9899a019793079e91dbd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc40cf89410fe90cc7b7b03543b5274ee9cfa59326608b8dcce4b6ea7a01fe0f57142882152641dbff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f50695c5b5f73a07ce7c3bb186f33e619f56bf642dbe8fa712ea9ed0ee8fb63e2fcc91140a9250d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h729297df01e82f683ca8021b14ebd91d18ceeaccc8c98a090c88d0450af38e010fed64248f6e36f57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5032e845c2b403649137138a6f09e51f18d425ebddf3245ab82e78ae634e8894a0a91b019d2b82450;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e95176ad5646b9b501b6d3dc6e83cf1379e537673aa6768fb022284a76b71ff9f571437a4cbbca37;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38a1c9e45cf95755ea5069d1cfb7d09a9f85d96d9d645c6f9cb6a21fb9e8b0733def6c7a1b870e745;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63698cc826667bace6de88e928cdd0a8e9b1a6a0c0b011c1b812360ae2f0bd8f3bb3d5cf1c72046f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e23083c09fce6c52de8e61fe6167d9efcf3fafb9e5638ba0576d2b043bf9f4897750a983076ad8cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24a93d191ee82a40893204e611c60b7e56f993e815db4ff16fb164876cb302469fc8926bb1b78c2cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41c48bc0d2ee42a9e1a731876651455045a6d5c0c45b5117cf31cd8973e2a8f1357b3bdb7feeadc1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h611c33b38a42ebdab760f0223f9b04d9ec15a9d657029afc19e95926870e40c4af44f8700ba970c3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h591c17695967e2dcf871c2f74801b09f81d8b25701c95aacb539e6700e1cbde7f09a03f7bbc895afb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11df5ca568634c4f1ba3c36631b430cd6d5fbe9ac35131ff13cbb23124f11dc08c7d15cf2622e309f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cb7e27f51790fe32d7c61f009900ef75dd1df7bb47ea7b4d17fa955ccf04b4da844dfaa4dfe1981f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bf20869033d4b5d4a1c0079ef18f4c3eed829c0dd8b0bcf803940413b11899cd72a8428a2387453b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha90467a4bff82b89964999f33a83828a947d2fd92a1f627793910fed65b2bbd968910cde8dfe8c74d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c058ec32ae2cf081afee8b3cda15ae81e7128f4ce53138357874a260abfc71b023389c0f3b96116c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77d8a09d9c79871131d7979262900c4b47233b676011d4c7b5c13656253d0d165c05a3a17f294e045;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98c60847c48fdeab8ee3796a69604db860a2f3d2488d02717d1404d13c48fe906daeb82a37119b60e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1edd245f09894baec5af73be75236ef03552e219e76b57d48a72594a3667f434f08e9d1397b06c4b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a67ee38965cee64787f7fe820ecfc9dfad2c657cf35b7d094f3e9e00c85a4cb9a676b09dbfd9e41e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75fd3712b64309e854d6663e47bbb4278c6bf5250052ddb8b2662a270ca1b2470d830d636729cce80;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24ec2d433c93787814b4bb75fd98fd771f7e35119e574bcc6adf37c5ec0418788df979ba65b5176fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcae82a8eb0ee1c652174e8efd7b2c06d7ef3f62d5e51493d60a2346d4fe653de68bbb8ee208f8e8db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c2d59c5d2cb7e5c07933704ad30b97ee5700ff5dbffbda7eee237a76d2da876441fb3f3f269c5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40ae40232e15d4b4c00a42d83754216a54dc40b094795e2aa71591194239fb8975deb5423ea1774c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc51a0dbf5ca1e2119be69220098fc43241e10028adb03a54c496309000ac5076626fe3ff08ab2ad4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc59b4b8b566291bcd9178992097d3dfce617ddf934b1d52c61c2126a8599f22d9458b81657911ad36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74484688502a37216dfaf4b071049b8f9ea70e8bad65dcf64984286acbdda0bdf070a7e757a08bc8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h760ad18bce1db858b3816268dca46e8f168055424be67e84920a8ebe949eddc06e6a513f07b9e73bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab3894222eea2c116a3c686e7234414845efbf5657e7e2968d0f896191f30b198820ebe26239b2903;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f4d4a0b2867d15bbb8221c996460f4e3e111f046acf81112b83c49f163fc0e2c41944469fdd587b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf37a1e245362d89f4683b3fc4a048f1fa254552ab8b7c4f3e80cba166c121c8f3456b0fb9a6b43db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf30c1af9ffc6d2f151537eb3dc7fc1bde62be608ce03691e4990a6587111dddeef525c47fcec1d36f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60f31c7909f298775a5bb946e3c0f3ffaa6338835af93f8fe7ec94d2f18017a073ee683bfbdac9887;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcad64f38c1f4d8c431233353a265f058c4aea100f56ded12e2c822d7bcea2ab7e029f183f852744e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h833df70389f9d23a5fc52999489bbec4a334a4ee6fe843ed78d2db70b19504e77e34e68f990eb820b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16db5668b8b24d87d6f1a8cdfd5258f91e11abb26bee147f996186371ed66976250fccce805dbb5e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4201d7b9a7697123a975383813f396510a74566e0d13a205fdb24424f70a8e56efc395d854bb45f18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cacd40520f6e6b84e10650e1aba09aa73d95c59750116db31dc3805a85fe769c05743f1943136e1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae590ad4a224b173cfb8e89d08d4c45cfd8eb21eab3d5f5c2d1aba2fd071ce2a5949288b682faa4a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5b9b480b6b892a1ea38c0a3969a2bb27ec521df0f3d0c8d2b8315fa19734674587c3e00264e999e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dcb8f3bbe812144144a54748556d29cda95522439f5556bf355e753bda61387075a72689b4667d05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fdcd5971ae3755d2078964638aabe2b91d2933b9d2e22cdd7e72f8d47a533d6f7ca26f3c5c3c867d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9f72e6d1aad220be80151cf9b93b9809a899c95e37a76cccdedd3502e6223d002ef866b8b6a6afb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h846e17fccd187dcb13515e772e120be3d14c01eedc76ecdd5d2f306d61c0dd16c21c4e4481f9f2f24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6b72f728d0c6e8f9ca86879727a2a664141f0af36472c42c9f69e1c96fd6740a19ac06ffc132d9e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f9dfcfcfeda86bc40a5fd18a6386191890b2698e9dcb9da4f87b2509be6c7d3a67d4be85c77d6051;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43908186cd42d03a6e74813e4a2d3347058a07bb15733b6d3ff6f8881c3df0dfcab386f03d3de20dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha144cd64b0506533051f2393585d22ab8bc63aab42fcbe39674ff6eac110c3a20eb81d36c84b18050;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6505b352cb2af91c4b45138560a2d6fe71ddcf659d008a4379523011d32057ca0d169caaa8dfb8cbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcbe17bf4650a479126970ecadd6ba06899180b4da891195c611ddaca53903e6069f0d0a7bd4c0615;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f54b8a2a99548537ff42de197b193063f551f5d31d73efdea16a629602d8a2c9ea0f29da1b70e09b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h135fdb50492f17b780086f9487759323df2780b303e294d7b6a890609b2fa10c5500923a3e25d2e7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedae338ae63622102ebce966f2048a1cd621f5313e26fea5a246361e72487f82a5fc8e634883d1439;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83b4e634e5a0a3cf13bb9d83003653f763d64b4e18b6517448a3db6edb22ef244292c01aa685abb36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44c2fa956030b3482ebeadf54bb2f5cd54b3a7bec0839b1ea3e3b47e7c7cdf2230183e686577f7273;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h439f963c0c5c182b6dd05cb588ecc9a0eb3696f26a00e5f38cf349e8d2cbdd15ed77eed9ce84378b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1df412cd35847ff5e2ae55f56744cff6eb7007528497a2d9007a91d56eba23cdb0f5bdbb8ab6c75c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6088743e3b2ed1a701a7ee58a2f00c44ea24790f8903c8a5ef6687fb6f8c8517c55aa5dab8e1175;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97a7e20b4ef4c1fe19b43af0a2658dc54f6c95cae87959317e08172bcf271389fbcd5c7949a5ecf24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7137f0d3f2ea44beaff47a71418b24e7dc190978cc8b7bb9a6369340f8e88d217ef27356453c72729;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d0789c16cadeea2db4e60c671d902f3b24d8fbaed5591bcab2da66407fbb36deaf247ecc76f1347c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73aed5fd8c9926ee57b08d0596afad49c38cbb9aa6c6c9928a4c60a265ca160fd7bb7e885a433838b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haae664a79d157db37d9aed0d095f50a4457957f98854fbe5885026259d1a7129a06a687d4d6db3b8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b359cc21e1edb8ec6d08665d34acf6d55bba074bdb689f824c7c1e7087bbd8ad26f0f27f713051e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h638d71f24211ad5d50841792f645784b7f7ecacd2a5bbbbc6da9e82af7454f10f20ea7948bbc18051;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cce2d007271303ced3975c02eafa1017fd4f644ddbe28e252b6f230e6af1ae52fc424df2dc3144c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f65840bf6346d350fbfc03e829a2573db4af68710b36c5db7c53c0517b04a5f10170431f1ee3d54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d830e8c4f800df5c670f3c8582ccce578fcaacc62a4fed071cd30aaa5ff85ecbdc34fae39d34ab5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4383c5183de2728d346964b81e998bb43cbe0f07ac0f1ee20663fd729bd421cb9c204be5d91b1198;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eaed48581c9c1e4e5f41d7ee985f4e45590c478ebb829b50baef9162d8eac84289bded800bc458b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82dcac659456bf370602bc0200fdce2d8783d93edbaeb5271a416fd42d7873e38bba858253772f453;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22a30890083e60c60b3e44f39f0d4a61bd1c088df5a4de1e7bcc57e44c96832631c56cf8da9d0c1b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bc7dcd975de697161e78fa49f96e9d9e5899e1b7c06a48096a94d46210b3271d5e368ea762f78a02;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0967dceb3f3361c9d645f58702286e3dc82b50725cc7b905a3f596b79251777c4fa1defb2de51f3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd40afc8734a4c124c1324ef4b974d81207e0c565daabe320d6f9d72ff9c5bf30820245798c3533959;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1137e926f9eeabf5e619802b6efef9997393cfad8e2f60bcecf4467d0c499fed41532e220d2f763a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64bf1f8d309bea052e488bb06bb05d160280e6825bb71783c51bb48a9391b8597fd6196f2263d880;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bb273e80d49d04a0371972adc99e5ca11821f2ac0700587df607ca906a255ec493bd4e3cef77b360;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc70b09dbd9853d5a52adf26dcc84179308390b636f9ec098f7b4664cb650ced1cd3f1fd75f9d56115;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b7e6ecddd03be3a949e3cd60156dc3213c65e60ae00459170b7769266c4173d1899d4756b1300336;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a4af2eba0864f74f1b64544ede06199b6a9e23974e9ea6daf891a77da957d2c5c1fbdfd9df00bfdc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd94f226cab5a27e439a9cc5fb32f8753344a388c484b31b91a4fdef90416d0062dd191948d7d388cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7adf1464f55420e2ce106574c2d32c3c4f3e90edb5d87bcc5721b72f969040de0dc3090c704997c57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ef182041a22cafdabe75eef77f5a9b8b4f0c67ef48974111f87841ea808b982f91daf026c8f731fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ed1b2fcc68696a4ba98aa5cfd02d4e6259969196d6e508dfaaaa1cd1534787eb53e13c79ca2dd154;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c06efad01d172c5eac9ef490e6f6b063d5d7e5e773a77fdcd908d43b9dca6a1ef0a9528bac06d51d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd755cc4dc43c8b43dd776f8df8d0e13bcaa5d3b18c1b3dc5340fbda1079716e4f430e1f4869e77e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b6f883af603aacd5e4adb80f10d5b3f797193ad635ed7cd758a92236150fead4d681f76374af96cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22f69112f7e9a351b48984c8c0b4e4afd8d39670358abba29e538d64301014f695141bdb89f0c1979;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb477e0b20fc76038388668320b6a9d748c03c7f6e423d4ae8396f2351d77535525053a55ac754fea4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9defb43188955ed7de958340ede32e78ae6e4949a6beddd1bb20d46dd09a94f2612672db90611eae8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ef74bf6f391b1709ef780165d6c03fe7f7b1b17d47d01a41fdd7369be779f94bf95e8cdb3dddc5c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h236dc677e2fcc85ac0090cda4cb9525d7d5783b3cdc352611911d6fc953b1be47afe304caa2cd42e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82aa4d9f14e0b41ea587f98b58142dabe157788080ef08be2ce24547c989200823fe32e26e895be7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h390d31c75fd0755380b1cf04b63a9ab70208ce55cb5488cc63016eea244df9bae1c494d0779304db5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46e2f896fd7f04662cdd1295f715711d6bee4547de00e19e570e8440b91f370dce75895a891ee8662;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12d354f688954c31f305a48bee6417a74ae69f173056ec17430efb5c9d82c216057a6735f6c2f8936;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h276a97edf367331713abf1436e1635a7a4871809c9863fe9cd7dabd3ecf829010bc622e8d84aa3fdb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7c224c709c307cafe44fe34dbb692f6b1ffc305b4c71580a042375ae6473528e99229be2e27d479;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78d270b57a035481fce7ded38a8ba35347714a99ebf558a75d08f37646437f66d07f2911aa9c1315c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ce0c32ee029c487e3c5edece4ea0c5dda1b2457493da6deb3e726d1c17278c90fd7c342b4da4c391;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd308d101512f426857523f3d04c153858214695f2573503892a0386d1a532506c9fa22c12acded01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6c8f88ac8fae9e23be739f193e568822308d9d6e9b090d7c1cb0a8e9e4c436a34f8dad8cbda6ca0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8255983e21ddec9b7160c48ea4795cd8425227935d698ecc008cb92290f22b900e2bdc68506f3f13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdeab2795c1abdefba9c88e3bd68a4c39c7388fbbdd2cbc2075b954b1236ef4d6abf9a1b0d5d009fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b6e9dd3aa20d8f6c93af1886ed5d1ce19a8f1a6af12536e17136957d609b462cc38f773ce88bfd4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0f8505edc9f1b55c71854f43f96071975c1b591b0e452cc94538b9adc60f9e435755b7dee4ad0bcf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88ecb62f816078032732c7bc5be86a96fd3a668917b256f0ee31747061fbd02442b2b04771a4b408;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca51f7b703e80d17bb737c051686e10e7b6b2ab84e263a0c985ac0afc018d41eafa85be736b6c386a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc16a5db7d313cb79119c1e5aa8513faf26f509925f962ad28dd4e1d58d3b8f0680dee1bfcba974bde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he45144e83af5701baf8ed7f72d281c1562b707655979a91641c8740b426d12c6f3b8b742e32a5b157;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6f3a8688bf538ec715e2022bd7c471dfc89429cbe18a0a587b3b3dec9814cc71359e589a273bb4cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ca3603a8fa35b313cef823174e146a8219b397fb679e90896240689c5056c83a26f4e0b48915dabd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa0ab3841e03981fef11c06586065dd82c10f2f5c9f4072d6f1f0cd6f30bcdcf76376b80609d3b905;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d1e407a05fdce50487282e9e7468f0b6c5d6457b9f349cdf28448b93657ee3e337d4d4a496927a5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb149307ac35743884da3e18af35772395342d41ed9b715597d21b019458945f7e2cf3b24c4e48a146;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h405a8c960a39727fddf8c5e7a2b05598ca001183ca754c9a64e7adc7923711410822b3459e116ff69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h118b2f1206c52d770254956372f660c8b3d6b678ff9a7442e8a57602a77c0b79d8a527bc8488a75e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h444d2c5a42f503f018c39ebb931d4d22e987e65440221999f401ad6f9d31268222b7c97141a5b97ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78610f393685a8c298a89b40cbd3e0c678bb717f3ed7b2e15b7d76c328b2e585c9fba48daabf63aa7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9abdeaf5e3d9fb685121249154590aaf830454d9004c9355e6d895016e4a2ba535cb0d3e8348e991;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37f6fd7f36d5b13609734404cd5ee6dd3def1cc4c45320d34b88bcb3883953c4a98aebb6b777d4321;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae5c24ad354c970fb2e178e979df91238d9bc7374a8edb366284b949511569a44aa6220eaeef9b406;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eecde05e0d6e376aa697a79c9699b4f6825c807d87c631d6c2980d693931dbdc82075dccbc954cb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a07bf60e5390449a471eff9533cad350222a22e0404e65d677464ec0709e9d53a3feb5b17a19bd9f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2df9e468ac9f65a1d641de1f62ff19de736a3f9340e168b525ff369cf322a247ff3114f44a13a15a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7bc1bd4559868bfbb13f4584d4b9e4b9aa98081c648023e47a0dc96fc2e6c6fc8f7c878f414d6c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb0cf859cf4f370213479031fac4407ca4684781dc2b5ecaed8dd46746bf038062536b5fafb56e006;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96ac466e62fdfe65cb416110babf3a7cded7726de684347f1d1a82b33bc7213806e5e94cf4ecb68a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2740093661f3f1c224451784cfe40189b8602a80db67cba509e7672a4dd24291ed4d8f1805e26eb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38996265104dda7698af9719569de26ec8b7ba4e12678211f531a3e04777049ff90ea8297ccc2fffe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b29a0bd7c8da04f963074490aad90f7efc2ef703df5dcf9585675c8dd4bbe1d09e0efc0b442be95d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0cb6a8a9da158784498501d27a3d1cb270d3341081848b92a87cd22cc1875a96024ef4ad8a93c692;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h540d2a688b609be5720aed3c5dcb18f01c92bc3015bfb7af48cd80d11c3e351fe75c4de1186fed140;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99585990def7ca48fd70efa194890d3c2339a7f231f3262be4fdd989bc90a9ec203bfe122be37337f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5d3508234a10a6d198cc3a0a1b5c761e3663775597c4e12385374629174e76e0813c3e4477a7e591;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cdfda2e3a76734c28873241b1554113ae50bfd0fd056147023942bdf17dc8947fb688d219ae9b071;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ab18aa0a521d5dccf80e6eab12e24f9ab821a193cb90c3e04aa72a802092976d55ec2a8dc6874284;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd07b55c0dff6bb29e1d0d1edb721dc2893e419b4e8c81e8daacdccc4f713f7738155fbd1e5d52695f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h627f000973358f0d0eec97a3b723d7f5cb7b058f8060ed09f578198cd7a319000c4bf971dbc2647ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha724cb730b8c4609e70388d7a3bcc1e910d445fdbbf2878cca22f3fe477aa83441320168af6358f45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1e5557d3abae4b5028dad70ec4f164b7aadc961cdfca689223a669ac84996bda530e576eec8a70e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2adaf4c326db38db4051e9002b44496903a53eb58f70f56a1725133f5512e98d2d0204941a5eb2bc2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1db3043f7bce34dcd72fbb3ae53d60810973f38b1de1429db5e29016db9e6c17afaa5e3d9284f77bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbd0b925849f44a580f50bc7a9bb65d987f750550ed18a3d782f50eb81519d484da020116d51a7061;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e334c693d9dd1c53a67972da4242b330904db78727833c9bd5fa7cb5ff7be64232bc084fd43fc9eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2719109e487bc3126cefa86b6351d00beb886a9a8e16354eb1a491334b52022f1173232889b2806b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdeac63a211dfa1c4fd91df254d573b78bf82e62274a64255f0eb05cfd8a2dcfcc5f25bb918c32c313;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h915d7d24489e05e656f9e79a6cac04e74224239c0689607f0845c6f765cffbe08cdfc00ed6763f44a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff1c899987132bc80f76cd1070c24d2f59787647200d1beee4f87f50911e657050b0b8ee6a678bc48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd672239eb1aea5b8c19ac02d575fe87bcfacda47790f93be1f95b66d3f9094b6ef1c5831f37442207;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h233c808bc83b1e4ef02f2aebde7044954184cce8dd620f014d95e301c6ebfb10b06cfcd6f1435c5ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e064980ecd6d20fe386f052e8f2edc0dab4b03810e12494f786f53fc9719a5bb86b33e2a86b4c6dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3186ba8b9e91a93d51292958e14afa2ea148125ab1de6b8c8e29307386581b02ee033cac8889cfd8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h803bce7dd704f8bb8335e3897fd359a16f85096700aec63e103c3998a910fd555f59289f699669fdb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93cc58663d3fb7e160fbde4fa30c54e513fdc29b18683ee3c1f9d771fb3c35588d1f1f1a7c81bf02c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46b9854b26be023aaa84242f34bf76272d449d5011cd3fba8713cc395390321b570c89226bec47486;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe1436662dd17c57c219ea70fe79462a992b2622cb2d8b785805bd418a40ca788ff58a79d3e125677;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e40ba87e6c91bf6e8df877b975789449311b53511463901fe95de436f3351f2161f0613ad7d45395;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4494f9b8d27b7a28008de59c4614668142e673f1668604c2dcc737165ee92d7a84f44cafada9649fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heee6e5ad56c9088fed08e6dbf5dd7460e9d4eb35d0570f66745e30880a978f8d37d331963e5f41e16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aab57e59638c1de6ebdc427540ca9829c5f8636f9245e12f9419212a534fdae98970b76ff9f8a37b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67276da1983824910fd24a99f50c33cb9c26258ef75c598105d038f89a1fe9087752d9b27d323cc36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84ce142f2658e9883d38a68dfa9cbcd5552558c8410dadea89467e10bf57eba020294fc49e8de4eee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea2693b833d1d13e8ed64556310e5bb8e1a792598df0f8810f576c0de798ff8b85a99dcf4025ed49c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff2aeb76137e54cd9520057ab2af8cf59277f3964784b21b308398781666dfcc29e31bfc18a09b11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd02145930d7861a533f29e604fc420042298310430cc75c4318d80f597f77d0bdfafe3c8f63852e3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf17633442d9377e7280b9773150e267bca5bedad4fcd65efc7ad774f3e472eefb190001ff06708b95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80893cf7b63c07b6e7cc703f38a0562623e3aaf233c894994d5756085c5052826a67a014de88ab061;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ea2576715a08462f20894e051f4a04b349a9e4e361860a1b998f0d3de650970bf5e9b9aabc0b1a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27420e66be53ff0bc71f98489015dbad1df08fe65ee34561dd269267aa56e3d886d2d9706bddaa7f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf908c24be372a180126282c69f26d828e52c47d4ab83f5675e9aa2577c109496e26fbe90a0027e656;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ef26682082183f78537e94569dcdf477f55c8772adca485ed7a76e1e8c8f79bdbdb473e12ab598f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73b9bcdad973afbcaa40281d272542e9336fc7b9424f6e9ce0de1dfd5ef765fe34171d4b7766d6d0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77fbda822e13ec35676aaaed4d1cd23bfc98a6421659b7f4793271310c6accf28708f8b394d9cd780;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5abb357ad2f9e98a551292365b042dcc5186ee048236bbb7a4506042df3fb3a7c86b89747464d7dd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69cb92f890a21300c90db367e6398f6c15f40842d579d47af861425c2579998ed7236749afb9307bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90a65b96c54826fd67098d12f17869ae359ba040b075649fe4208de99ccef670c8d10646cfafbe79d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8fa1cbb984b24e96cf25ecd3057774ad3e24b9cb6b5f9cef5e6194ae5c36bea27e8c75f98eadcc81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb44442357c1daa29ad44253019bd043327fd902adc7bcb9074c0deaa8fc90dfd8a248b60130e79d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2998748019fee2a4a8d097b5f4da7334ea26050d935267431490ffaed414f834f9c71ab8a78ae0fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8c3cf84b4dc4be58e2587aa663252402d794c14b46aa26e917dfc3a3bcd0b5864304f1cf9c86c150;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb92bcd03e161460f98073166861d7df2431a494697fc56afbf6fbd842a96d83186804a99b4d265e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h893beb6d6bfd9ac93e1903174639fa96f72319a425d58d7816800de979dd3706c52095ab12988ba01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dee866fb5796ffd9a8d62d8394c399d13ecf55d798856344fe550519f176463d748cffe58456243a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h122beb7057bd47f840dab20c214f92fecb7c09139bbaaf44adb3b6d48a7bf13b53f9102d7be416a85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h233c810684c33a36021f326a93e46ad432a85f36738c2c24d67831d6119822ce63942117dba31e9f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4977672beed7a6ca2955a5f79edcca550329028c3ba0b40f7034a91c9c04ea9aba9c3c6bb3849e3e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha03cedbca33a894fd361000c4080ddf47e0c95893b2c30050cb3dadc6d152f04ee6baa5e90686f448;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fa9f3ab317017c9cfb38535092cead013d5652bebe74f163ee9e5a0ebf4a6e33d9b56183080af2fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9dd4c4b83917cdeb881868e7429aa48e0dd5d5df11de6cd1e6cd5f7475bebef8faac097e67d4ede3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd193ac23945ae1f06b42d8f7391342a1d581aed8f26430318197bd0b30800ef4a2d34dacfcaccd88d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd59b8e8ee82624d5b40b139ef390d51ca311dedcae85885e4b61ef66e593660d7f9b8c515f3fccfe1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7c38c446af784bc1f4cd2827e13f1597cb4b696547a6e72856d714d33fd97d5f9cf55b79a8f3063c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3be269d5e7984fcc7fcfe70f56d1d5a873f1dc615c3809094b642a9646de24d70348bec51f6ef28ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9106a94209e33fb1561784d4b046c6f1b1e1d27e8364adc2a7470be01c7a4ffcb0256f4696524d03e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc973ebbbba722a4bfdbd841d2c74694458b897da7f5dead71746af791c5d7b5c17389973147cb0a00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0db90faae9f09248aae1eaa334349a819295742c3975e7003e22b16ee4c8ecc427b13495e20c86f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8314856facf28b1b464bc2cff8274919d60596aa3b6c4d1db53714cf48ae71989ac066c139406a76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hada50076806122f23b2bf6e90dfe33b2f1dcaff0f143ab77726f1aee5980c510be6223aafea8d131f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e01403a861ef534a6ba2c9b6fc87d5c27692253f5f5ec4e93cb75c0bade1cba3b1180013d04d766f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb552c9912f424acd2aefecf43d9865b9e95c37b70857336780c2c92d482b3c80f0aca484343f80f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7704a6735083fc5c0744b23045701f509aa333cacaf642d70579536ab74e8c98525a621ca0ad43a2b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c903ebc96741d0181a840a2ee4bbe599ea6bec17ec8e7c73b2ced115d242e6f973fb124be84652d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c8a5ee7ba7135db2d863beb5d1f5de27a3e384cd0d111d7c267d91475fb35d62c7a72095319cae48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h661cbb46d46011ec2adee7f1528c30fc6cc1bd1ad67f0b85f89b565aa09932de56351b5320013e1e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf92e7d17020dfaa70539aa6115c3939b88e0f3db192d9d26d5e5db217877952116207e27161514883;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8601e51fef3cea39bc524a926961a61ac9f11cbadab1e434fdce46699a6faa7732a4d04386bdb05f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a6ffce857f064def34c34d08068b5611a2c52a24bbc23efcfe242d8279bda97b3b4b8b080a5626ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfced0428d38474ee44e67bdc7e715db61a70fc925b34d32b3a9f7b7604795205ff678fb71b9b7b4e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a9c59ce88a703cf65d9d9e8189d69374b5ca8cb76c2d0a7b25238e8ecac4095e647e83d40814d4ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7d4fcfa84e475a47626b937740f0842f150ce6f38c4c06746670f33a20bf042d3ada5872ac682098;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc33e9e1f5d793ea93b013c3d85060e99e6eb4a0a2f8b0632db761f51edf0df9b46f9813295e6fc11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8fb7db72ba017171dc389a5cec9c9439ca8a1db41161addf854fe03e442f0579d44f960aa4c492da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4205ad5e6b4da8eeeae3744ad4f5d8aabf487d152af9e96190fe45b1f74dc0471f8a8cd14976090d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7dc790fb81d8903b86e7d83b893f1d837b1558a3240ce83b8142bbaa1ea0f97cfcd18334e08cc02c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7333203bf7a5619ae2e30a74ba9d592f99f9b80b5466e48c0e1ca270419071fc20cf93b85e06da7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haca5142dffdeda5de9db730faa8495e9688a9b8c2d2ed96c544a15a08b1492bd5b592c5d8aecee449;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5b227dd60c1207cf4e9b78943fed5b68787c005b8e3dfc4ef2e7baa29a1dec2f3ac71d7267f5c0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c3d5f84d0f4389ac90de13eef420ff0bf5298ba5908ebd9703e2095b4911fc4b3a2e27d5f6f135b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0c74d13414dbe1c4d6feed76e0b1a728b66b2595d044467b8a55fcc686c28d663297d0a8b878720a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h942e89031946353d32d99bdf8cd02c51f8a935c086f20c858c0de84c5238f386986fb83f3b149008a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6648f7f718caa87b1b3840d0a3baffe82ca32960f35f2adcf49652e5f9166e7986893ffefdcfab69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4c42d182cd3c0c2dbfb06d3fb8215ec0688e34b79da3898a14a1f299b4a4c1432f433dcaa2421ad8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7859b79b1aaaa182ba6a27e5bab9e8ee838a6fdd67fc906aaa89dc12bc2b8ff93c0241dc7b6391526;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b3460c9f4fa281ee922e3848b58b1f01c5f92ed78a6c894d7142e4287b09ee7d5bda68ad091d1f3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14730e8b84fe8d858c2895b52e7036a7f75d5181614fde55f8d45826341eb5ec31a782c83db7b0801;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4961c397b7fbed8b5416a7cb2764377bde3a4854a29cfbc146cae2a622bc35237a5b007dd18cf970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7235e4ad378c81b0ef2332ccc8d21913cd4b80a0eddb348f91512b4954948f038ca926ddd39e22bb6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha19d0e9fbc6a25baecdb14237bcce7dd05293902e4ee431aa3801df44d6f9267754e0dd59198d72b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f5c5888d07c95345a9e20762680a5bc4d900a2051f7ba71dce67e56c3c3d28bd2293bcfddda73b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86f416a54414694d4207805f744f8afac3cf7fe2a6510b5d7a8c76030950b09166de3b27547d7070f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20f622f600e1339fb9b0e32a04e91a5fc479b6010224464907404f42030fee9daec220ab85c852d87;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8ffdda09000d3a87db3c6117b655bbfba36b40465089ec163ff8ca6534c1109b7f80669321003851;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6044ce15dd8c25135d605d77b4c38bfcd766ea194446500538bceaa02ae355f0362b277ae765fed13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6c7301783f6da80811a5b385e6872954e8b88a82d08b51f2d3a6f6642bf8bd90350b34b482f3bdab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8929917b17ed0edae94a5352aaea1932b8c2cb3f16cdec0666063ca4e1c6a921eb2e3441e96fce95f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb66f5a5780492755c3ede99141d3d4fb5f1087982f57bbaae220b7b801b12c7e3914fbf8b8279bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h226bd701485ae622555debbf1799d63d28f548e7df4e19ee9f25d95c8251757e159040f9817517284;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc4ec777607b1fcc76960ea1eb8324329a399d8a6cbb6b16f441045d983f15c39c1aa098197846ac6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb17a15d29be687a125050945ef790a5587fba7c1e5f9316fa2f8587173d2dd3f60fa5f458eecc2f55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab92aab3a867b5c332ea57a4e426f453bd1874704664719c2fcad6648e4b8d9bc966a0314e5aef37b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1572664bee8c2a7223317207a3f9b112627f3ce973f6bc0833b5b888f1ffc0713242da2e160b49287;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1697a2b6c161f601894f5f8557aeb9201fc7d892afebf9ec673663be95e7138b056522e7a47009e2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc497985be2a2233e40402080986b5750a68e92b6cbae33f870728e99881c6f1a16aff617e04eba1a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2146854f2f2ee5c041fd65f5b90485fb1ada59a0557f499105a1fd54711cf88a95d8609a630f55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa216871684c2294ad4ae3c5d39cf485199cd432e8529f73d297bb041f66c87072c0060a7afb30da6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h495d124b87bebe84a9dd8916b290400c4793120d0e7536af07703bd9d2f7df45ae74e7cddab7c7b6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebc2c27822278049f0f187f9f50e23936a6141a863cc71d92348c31a4b6b59e4dfc9f7d0466e80b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfec17720eb745bb70e6144a963e5d154ce3a9555d98eba9563ab236fa75a0af3c1c636dd05dd02a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h328d75cb9b504a6235c34b8d482b4a69e0a6f33f410b6bc6c23deb18e6a6e64697ef0dfc77fc16c4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf3c28f10a5e630f80fe2d5576809eafc34010e8439f2612ff8c4fbde5d95276d4f61d1d296b549de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ac506e6f5b65f9e81cad4023c99ea5d756e7c8f986ab7db14b9ef018933c26d78de82a5d89997bc0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5d75ed607873d9e0385ef622b780cf7791553de2f149da00e44fe80c8d943c30616c5fb207036e63;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h380169f76b5039b712b47784c85e4d3a820dbadaf4df2c6ed187de14819196c3ea7252936e09d025c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26dec39720be59746b1664dcc9bfcd0989f81dbd60a07260ff31aa220d627f4c1e79894114ca30ce6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2e257745c34b3150f7e4bbe5d21f6bd2a83d54c56f3c9faea9d98d613fb1e887af9f50c215b0735b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ac67f26de64802df062698312645859a293e50922f5771feb2795e1c839b36c2f9f33c51f9cb2640;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a64c3b7cae549522b2f3c313bc93891e587c41bc62accd99e719d75a328a1d5c03595ff6babe9e3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c718b1851089d69933dc5f0feb8fc294678d2e94924e595a2c102d95d57b60b9adf4a1034ab0c19d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c9c6bd40185905b48e24d6a8de2bee2ef4a7508beeb310665f951c568c53cb09b4c258c1896c414c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94c62aa8ea3335feda167531b7658e5366ac6d3775aaae4015b10860295bcf49903e2a812e4c02383;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h262a0009cf26e0e7ca1f10b191990a717b1a02a124c9cad49179317c417363155e96513782a3bbcb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50b0e2dc39a4dbb91f80eed8425ccb59d28ed1f13fdad586840960fa8d1e419c2a8e223bd16f620e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdb91f7be9689c6f433da6ac676a29568e6b7c1acca0fb20c1762e7d1715517c678f0ef6a0c3152d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha497bdb71b034d00b4a12a582bd6ed118b91c154d3ccf565318881fbee95d1a11de9546c540d1fe94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7b042191823d5d49eb6187d4a278bcd04ebaada8f2bfeafeb22ddb6f9a07e77a2e295163a97cd3e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h781fdbbc585c5992c97badd83145ba9972d14da43fcf17c5f1bd7aa11ceaac3190298e5a8b7b22dd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f44683c1f0d860962750775cd81fe0ee4edf19e58ddc87c5ada7b4e6fa02c021745cf34de20872e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdf4a16a246ea55c81116c87a3a586958e27da0295343b697c3612e6eb64db022c4cd02bd88ebb9ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8efae3add12c978de075331c30c915aaaa4781d556bc4935ea003974ec8e955a7c446275153221dae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2736400e379dc81e8314513068d9f9842170ac2d946109f9db66c0835ef4a3c605e4a97534c3db6a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc34a88ca5517566f854b55b1a8ab34ab7eb75f27e6d49a626af92a0420038273f7ccf1edbf0863b04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92bf6485e7ccf1837b255c67bc61fdc0ce0bc69d03bc944a6be1e0299cc3aafb9ad4a4cb2245ee20d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29ef092ad971162dc522cf48769563f0a618ed0e24fca6e2df707523122b02d620bc68dd1d28714f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0669590e38c755072f0310887e8aa2788b7e7dfabfbd11a154fe01c11e43928f15fba9a0fa992b9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc5492619d83d301b6df8379dd20369c55baa8ac4dd41762a6d2e6395bb8f7d360bc57e56cad7102e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e6158ef6c151d2e8dac2b6089f8c18e5f9c68b67084ab7ac8cea48d31cc929ecfd5460247c56a524;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3013a1cf3cc43dff8c4a40acc3b8775edc34b9d8db755587be410bc7cdf7c726b9b51e57dfd6ce983;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadac850176803c096f914fedaeba517059b72b2ba7428f500af8fcaab660e0447fd5f4658aef94ed6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47fd787488df5a8e92f4c55749239219dad37b46d44810100cbe7fbaf93c9e2ad1a7939474874208f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h617c99f32f45ab198a12734ff02645912b394b3a7530c4cbeaafa249a52b3077495266f9a501a8bb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3b7e1ed6a75c6bddc7893df2118d0bf1887a818fd8783bfec4b18e0e7d69fb408db796f156c946ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1632684f2f5aa2793fd6ce6534a76c189da1cf6f336c52549398e3701fdb0da9b3e1b5875f96174c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h988e54a0defe5ec3be984ab4000ca8d2d08aafb9cce00455c2ee5c689c186b4210435b9ee79250947;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70c6300acc453e68bbb64de11cb01bb4955bbe06f71fe8ccd5d88721766929bdf9c36af411b465414;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ba8d732f505ae5a80a53e38b7a1758adc99b22dfda019405b3ee990b8c76c7b94982e9d3b35f3fac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h492379c5dbbf27bc29227d08de275146eb31898506b41477fd962c031243b35cdf849a11d9d306897;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb6ea8aee5d9bc4b7ed808a261b611ea00981c178dc7ce4f1cb19f6d74420b57dca36b11e02f3d238;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ad8f46bd73cdc73179276b0fc455c8247484e3cfeb5b480f837d392c543ffbcf1afc8a2610f35b0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fdd2e116bdf4a2ce5cb7eb843b3cbefd6d28850e18c4f58776594d9db0c2b7981073489123094c41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he74d4a27f5bcb6951c86c78d03e176793a570e69605550a5560a1f833b510114fdfc815436fe969f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4347b896bccce849669dc15be5aa490c6ca3cb10b5be760c0e4b3c87410de835cefbce7fe78eb35c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71dbcfe3723a496ca7482a4b1ac45f8c116df7694466eccc7ce1d28982e557dd3dbc4908044392517;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc08c39ecf7406687888f4f15975d6afebd47c38c241ab914fe85a41a673e2d6023254e8164a95e219;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda459116b678cc17d6e43c888f8c6993338d5cb5b8d5f15ec03563e393d444f940c3203cb64ab8eed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94446277c2ce0e59e1d83fe27ce8934b82ff6fd280a981a07261f072032080f73dc83455cd26c4866;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4bba5ab4027cac978765621e11014b5a002225668e57a2a9d94cb78e45c3b915187a266776d75385;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc32226b0c4eda15447b1e282695316f6d3d9d2fa2bcb253d8a253e01964762d6bf3e8e8f1bdf250b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83e30a5d00c41278c73d3deecfaba7d509326f836a655ae29c2d5e33e1740013069de56373df29f86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2d2d4c0e67f59a7c6e8eb63332ce8f7ee5a92d6f3d09ed558804407fa3dde24cf4b0f7bb635f554;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1093e67fa06e1d39d56d5239575cdc327c1ab1758d4841b0534a52d465dd83b4c930c8a3052cab4a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68f3e9fa0d1a3833cf5bbea6d0b302fd4a647e96d0eb296ce4f68c853b84db6e049d78c3365a1c3a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h753edbfdc92555ab1d09084fce0522d9aaea76ff4d54d07ab357698469793a9b4546f298ce7681624;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec2debf30f1525be0708dd797a7477f0320eba19709cea6aab2d0e52e8e3d791c92373ad7c838733e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd950d1eb585d4ab3d66d24c71df142e0e43c814c6460306c0e185c04abcd477dcae309f8fac4bb38;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdec6ebe0aff10aa5fb38297c3d5ef371c61178648cc408425af8bf9de49ce74a6abe779b12d9c590c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he04e3428ce78e4340abccf95aed78c0832ea4b5d5496c81b58c837d3c92fb5fd11cace9cca74d338e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f3e107fe6fb2ce3d7574d05eac8c0ce519fadaa68d285820c1fcb8ba76c49e62c78cc19241744cd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe09ab08cdb3e16ba14ce8db71159fa312d2537bbcc9e61706b653a4fb9fb54886570253e9bed5649;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a3d62463f1e486f050556467d88be4183765265c33999ea61256d5fb624ca8d909a46facba3ec0d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fe1b93910d846a2791701b056c21f8b0eaa79174db885212faf62b2c48ed69e65381db67571e79f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94c7589c3f7637d1d870711a018406f5dee834f2aa48eaff4da8ebd6e74aca11fd71922adee3a29d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc052dc250bf1fca8f7fd863595fb4c7c10814a466b79df8baa6ba9d9ebdd36737585a2e72508b9fe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h276f6df6ebfa37d51e7ccee7e6e4974bfd2b360ab15180044a71105c53a6ca93a9b014cbecb6940af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14554a147f80e4a726fc833fd74ae335e17cba24636e144dd58c7c7fe1532ba93485974829ee0695b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e2a0a55bda476ac7e7d79b5d58e899376f1ad0091cb0ca0627dd9475ca302cf920619bc196f72650;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c0fb31bba1116715175cb8f8fbe76ddc75f65195ca691d06bfc70f6615d416365beaf9a0d148e8ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24baa84a27765e9973a60fe72bf1db97757c045de5462253477ffe48a4810a9b988b8139650a8ba2e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc28becc04b64e34700dfe215cffb73ccedf75c57d45ac8ee96adc82c9051d57b9a43f3c693b67adb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa3eac34de45b12348232df7cf9236ae2d5bb0956f9e1a832893b02bfb3855c2f948b514e73313e46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3caab80b516b4a8b1febc6a448a25c4af277475b46018addd9652d210f930664856317f81eddb34c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f1e3f3a2b47573036dca8a78300a6baafc2e34a7213737e80b3d1eb288802455f81f06c329352456;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h654c23b8fdef5294c4db2a34a780982f531e912ff12cd588d1141fe056673676ca022f14168cb7901;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b9150da2b30684f2bf3db69f3eb8a9fa5dd596b17b3c7e05fbd0ea05915fc14e7bf54c2811da4b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafcd0d962e55602ceb1775c4fb57ce139f7a5f7f856dd21db85726a2279f1d95ffe17a038345f045;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h193b74356f8d60fa5bbd505ea9e90c1484ca99d4bfa28dc56a852982e2e292f3f1256142bb7719875;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbd1d9bc737722f2adc42040674b82cc01de8726d85c545c4dd3a3fff4f0f3e248ef9db3cbbb283ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdc3dba7204ac7bbf672696c9853eeb1dc5800d35c587c0152f3d0f61a1005f198f2b20cdbd7c565e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4eb5d21c2776ac4287c566631bb93b43a2a8e753ce8f728de938a3c36cdcb029c2235e5ebb48590e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h121c9a889c491bad8df4652fe15bd772d0bdc84f94c806388b9739043e275e6e8f811f3ce57973903;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4856daf9a4205d6ee42ec03a874e50339f37e0cb7599123af705e70df14a31e5a03ffe2ac681504;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf62b8a23e0efbd47f649e1af1db4d41d9cb1e618bfb5390798934302b9398aef327a65dbff69b0cfa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha104ccbbd382d284d4638904ce43a8affcc2b87bab1144b94964e30e33ec4d40c319ea4449daf2aed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h979c6e0911110aa9405ae0215b42787257e9a983482f7c4ffd898f1a337d75c00221ae5cddb3fb56d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94d7c919d16ecf96db51b362c8d366d67853585ad33493b99d4a8dd0cb7a1355ebca1202482ef664e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73ebf0a3d789b4bb3cfbebcd0a32ee9e204611d666efb5652b95e616096221ac2f849d28c49cd01ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a9b7daa102e8f3678a4a262277aca286ea16189c46d62680ccfa7990961e7ae01ca42dd75f6a4ac7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43804cb4a5a7714be7caf44d1a48da57a1b2c351d9b28d406c0081a73d8c0f3fce443163015577795;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf503801052a30cb354c9d5a111c1b91689d74bc73436956d944da39083d7d909a5d236a63066d3166;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf02ed30a46b80b11a5d75b3b9d837e35e7fd0ff249f3fc8366bbfaa2443f417137589d5dbfd16bad3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3985a04aabf20b5504972ca780daa37b978275361f95754178be922bde16ffde60b66162e3c962939;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b5ad79d056766dcea167cd4a034afa2e9282820f25417298ebd1711cdeffe0c229465b633f824ece;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffbe8ac62dac4997e658bd8ce68208f114236a00041070dafca0d361877d465c19517da10390002c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd407dd1726a205ad602cde2a0fba9915809f5825d37c4a849f9a4a32527738c0005459d7dc4243d7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4da1c4e9e6b6e6b6828ba662cfaddb345aa65e6287efbf899d38cedf3f94fcfd762dadfc12384407a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7501c537ea090570a387dd0b5abb2e6a072b533c071d24002e58ab5c46a60c1419ad5c6e25a9b0d18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ee8e3644d46a9f2de03d71b13fecc907f84de3791b77916b76ce6c3a65103686ec20569dcd5452cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8b4df5b5a815e1a9b9054f86cef27f518471b74bd547389cd4c90df876873eca5b64f9163f52730a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1de55d6b9edcfb09db858557152ed98637552637ebf94dbcdebecd48e4860dd7217771e384e27a93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f38878bacc5f289decd3e3dce8b136cbbc4d613c2964f50ec4e538faa8168e7a4d527ca48a46a0cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f3fc79a35ed5e71fa4fbe9108a545058fcc591b21a4df9588652bca17aa3f7e38d6212d849b3d2d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9287742aef1183d4c444c37eeadc21b554ece6ac856b1138aa11dc368224493ebeabbf279c0c83c93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13a264724119effdf1e17125016ede3483b1b13f11c2757bd57a5efbbca5cffd3ffaadc4528983a33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8851eb240bdab7d5de2cc87f74a9f65437bd7acd72575ca26b9f0ab0982563091e7c586746a7ed9b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9c3adfc2e530d4aad8f308606dd7598c44ffdb46aa2e2209b207782827ae05fdda210300988f01a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99d2993b248fa649b34c49ec8cfd9508d5031a89dcfacf8c816f49491ea38b4fc434058c4700b8ff1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea8c07ad0abf59b9f2021fa1a9918354e7d4beffeb2aa09e47db32d2866b14859e48fd6d7c19b54c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac0c168a1a2afe472ff7421901d0d93d567f1efc139ab2e53f44e00ee1f72e6cb6d5a968dcb92e7d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h884ba63750e87ab173b01c0f3d149da2dc511189fbc8cde510fb19b3769f6d0448116054aa28a273e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a07a83c39bf651eab0dbad9ba81bfacac539602305068ae0b3af7327352e879ff0d3acbdb0d31ab5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9fd8dd24ad363dc58235b85e3fb7efddb4da6ed0408374609ee7cf580ea876c65a45aabd3e06bdde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h136508495836c2ef09173294af6edf71fb8a1fdb7cb28bc2ad5b117c49ffc09179cb71873b3cf109e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26f56ab227e2c868f65e8371f1b70a3a119be3a7b1faf99a855de747b753541cc65d3cf51696f3b86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e229d5502f97949bd0b4e37b18b4d61527958a4cec81f4c7bcc8ddf2a910c9943a9aada2b40d707c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf47ab90e9cf5dc4a81ea887bfe06ccac5bddcbdc44ac96ba93dc4ff8cd07cd754ff0501e7a3991ffa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haefbd81b0c956fdc1b7fd58b9b31df35857e814c4263d38d08ad6c1cee5b847d54ed153965b61e24b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68cd6c77360f3b04b33ae52a7bb41609aedf78bf1b0abc57eeda70ad3d9759fefdc3068149febd5cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6ee77b8ae435acf71ab87439437245353a9d26d502d6d0da92c6509bd138298d71c92fcc797897ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc930a023bd3e33197e1121b6e0748383d5ab4d902e910bfcb392d65bb5c83017ccd632f6cf3d7623b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbf85d6d7ea937d226d86ef16e01924d6f471c73e3054fed225bbfb3236e956e623a036c019200133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he300f88b613a47a63647df35e71a45edc45cde33f6c005f9c364d89559f937cbfe165aa6c0d32608b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8069e2876fd037664c999cb5a5366602194e3b5fff0eb7842b46720cb3ae334b24edd2d959e8863d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65b43424bd745c68b5f0e482875e0ee586ad435f0a8441c1db82c207ab0d91efb86ed0e070d8b144d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d650c4aeabfd8ad363e1b0ce3d352cadd956d021b5f3e3ce3e822c2dd680006ba858e9676dd49eb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf54fc175093b84ae13a1663804eb44a955021e19e9d43197e25ac3df5b51b924e66b1701dbf157a71;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17baecb2de45ff223cb61130849553443dc724e27b8fe66982b0e7684aeb5cf963366182be055cc17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c2eae262dfd5f8f5d17e8ce4b59534777c256d9ce318c6d6ffe7cf775abd97ea0bfd7d1fecb87d45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33ec489cfd35887abfe69cc4ef631d68711eff969f7f35830b306123848734b536d9b0c1b037708b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7166ecac37a3240fe1839261e3331590a62e74a5db338ae6089063e10b87cf7901c9ff07d3cd94989;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71d95050c7a54e5f3091a6f8235bbebada26184239148d003fc63cd44221c09fd5bdc1440f969aa92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdef79fddf6e64368dbcc498ad5a2aaf51d66f7c7e4ebca25f114773cd9f883ef2e5043c6e42d28e15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bcc0947dfda659883da1cacb0b79e0ca330a13650a465a1b768675f16740b81c3a1dad94a199f2ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h192553fe1241d6d4a26aced4552ebd05b4c9ff6808d0de54c28f057822bb519fd747466819a6512b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7939e79f5399018c117eb070901be2550f065fdedab730d9b1d138267e67c87559e71b06baaf1b5fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefa4b9c54eedf0ebfd25c62cf4a11438ca1f41d313cfdf05bc9554992f778c4649fcc7846528067e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd1d62c00a85a6ce3bc1b6f29239436d008c78235bcef932b1c3d54e06bdd982843a335c736cc9298;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73e0ebfdc27eb4e417780a8831550982a10cbb73beda790020d3204d3b851db207352c5e17b09a236;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9010ebf0c041155f8df15ee97130a31745993d91cc30900f83e066196a85026a1a75794c66dc3dfa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb72815426962c321a2183d9d7082a336e0dc9b67e37a30a1fdcaf528c70d6c5e491ce5edd19c8da72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7410d91503524751ee8a21e1c9d7b57fb0d7f494d7af81d303bf769851b98e9cd72c54227f35f4a35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h639b13c725bda8103b3f4b37f6a51865c9c4576eff30c0ac5d4b5e4b2478820b3107c68b51a61de3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8879af20814ad8d406fa7e394247d66d7a6120e45296667ee705c4a2f9a0cf2b82fc3e5fed657166;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfb4fadba82224da2a3004730e09ad99448740655763582b7b9ed938077249c1f7c0901fbc8c4f739;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e63c14a4d54d0be353a49e50ddb6f52486cc57f5184e8ae2620115e7607870d4b958e4cfae1334fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99cc14acee3222ca0aaabe7708c90ee6f9554038348d17cf56d01bbcfe9e1fb9ecf8b41bd5fc7fff9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb320555dec80e808ee207fd3774b3e2565937c2858751329c5974cb7aa090b5f2a0a8e0e1224b95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h760baf7a7675864afe4179d796d5a97b8e8bb55d39afbfdd724b949b933bfe0653e6dd7c616694c14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdc05ae1883472001114d31c04a83a547204727a1a1dce6ebe83c6320c5b5e4e539b3a72f29572fe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h274c2611a55cc683231e771f0a66a497c6ca0359981267118d3e5fcf6a0278ed82e1aa8e56e5061f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbc6358ef86d424b130776083661ca90967f9397c3bcd5ec1999b318b4d4f98b3b60de7856e853126;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3018c07e30f2f8ed1674d2480f210c2dfd800b0ac82b49fa6e2070dde895a50f037a13df07f2f35af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47bddf0dc206f3930bf309e031b152f4e2892920143a0ddd8ec8a6d5a46147fd5b7173638a112e4fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78ec4bce445df198afc3d600cfdf0da5883ea2ce37b1e91d54fb5d074e8861bcb06eeaed63fb6c026;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6a1c265e017b6b956ef11bdc243da4cf0f4f8f7f71cbd8295015f4c5acd9c4d1c5ce25fb1eec3a2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb198ccfabee4c6a7bc4f74407dfd5c3e2b93790179ecee28651a289ac639d8e3f24adb129745819ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3fe231406626e5e49d2ce53b81e01e84e151de5cffb30f7aa39a69d60fe25bf6b75db1080689ac85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h381e2f25866bc5435108e8d9af7202160837efc5120f7f1a96b2f5aef4684c5d38d4490c77f6dff8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb29eab9060f7db5ebc979111c4660de6e589c63901f93eb4f9bc1dc3386ebb657c38556262a4b806;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h859bb37fa39bf62cc8dea1ae169bd015f22068d046ca74d58c967e5c1157c44faf85983fd29708281;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75bef3330421d6763fb2bf032981ddf0e7d22b3a61a34f3a78790181355296b2d14eeb5033e808a6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80b12768470c1662817f3b77922834029ef7670e9e8dcf6cbe17882f854301dea047d4da894c83b07;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2901f0f72adea29d6574183daef75560a5f6dc56fc11b46399a87d743f3e954e4a8d5e2885e7f24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba8624d6872de2ada85ee443d3692eb4b6218c7eb8aa5518bd3374d3fa120349cc8aacb334cf97b95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6b92eb4c0d1a296fb00488dacedde6ef6984b3e4c33e0cfcd0e68f123992bdf9b9cda5dd07574bfb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc449c227e1fa641355eb5de0f0ff82692ed09ae3aa42ea43b43d142f4683d8095ea2269678748e6db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h662b5b2541a65f711522800b22bb3a3b0040c16b6efc66d62d37effbf08952987e0f3ad317f449c57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff893b3f2d5a3be9aeb7af4713439e057b4f5ded0c26d2a078a6c72d62ec3e8ddf416aa01f4a546c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac0a5ab0ec19f205fde177137843fbee6e6de6923f76a589275363bccc3264fa2e46f1d1772aa2a9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7883ba37c3564cefae651b69d82ed235426c6037aa1d5c69ba30ef30256a80115e025409b0b3a2e19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1fb469cbe1a65504c7877dd6eccc71fb57bb67d60e22e7fea925d837c2aa4e30f2f7f12f1bf24ad0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41a24bd8f8e7e09840e03533aeffa19fea230d32a562ce8db5866c2719d4af430fec11e999a706083;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h448c6f69cb22b133619350f4ec4735924465c5d452eaf60ca456b16faa3a599dd591828aa5178d529;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2eede4eb8b390076caec091e16f51fe11341162dcb7d60746cf9f3844509400d17ab677063a32b082;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca85e854b5a1b180b61ae9980da320824dbe1a7295b78c448460a482cb8bb9eec3f6e6c46133a8c93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee1ed112a3f10529de21d89b7300f5c335caeec7a0f44e49d20672a50cc04249e3a6b6e7a73d034d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c969402054f9eaa80e0e40df59f90d0c2b2d954050439657ef5b520ebb4bf67688ac11071e884cf1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf254b5f36b3ac6dc3b098f89764f58fee715b71cb368dab3b2224ccfacbe29e53c87f095bcee2af15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd69dbb57c7483dd8e555aacb4b97228734680ba8dbf78c183765dc6a6370c1de49c92f3c5c335855;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb07acc0e3ad1f438ca96bb01cacd1b77987b9e31754de673f33952ed16e5b1445f7b6cae1a7e69ffd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bcbe42b1b20701196346a15b13747840d58160d40b281ad31fef95f917f776dd2542df1667bec50b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h308ad8b21badc0f4cd822bf6bddc7c7f169bbf217b32599e47c502b18cf7d57b90b33bf2772e5af17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb15cc1af34be57b17ff5eb617441e3cb5d8d0adae653455484b539654cdf2c43caa80f8dd6fed5fdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b71957d336263fa207d7e1bd5a2f06f389a9858b40d4c86c588ccd397cb98e7075bd632882e8caac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cd967f1d184de8b1a6a8c71a8409f8cef18de7c15042460e5176010529e1ad7d3955d3bb3d5ccfd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9daf59b6d0efe600e5f1fc46aa76f33236ecbbc304be0bcdb9873c570842282bbd77a9ad1ae4934a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc22686d4393af9f9086843fd660c3ea42a16e852d2c37d354deebe458c521a424f5f9db8e0c94df11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603bd6f469e98e7fa3a563d55555f98a53862a06b29fa6dac094ec9c0e1d01cc750e211080cb7fbf9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha07194747324a58840a3eab1d9f374474a67281ad506e5696105400dcc4e5a3a8bddeb335c1396c22;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ecc3ed096a92ba6045bc8bd5dea41c83a255e1c49350b3545c8d3858440f294954da22181a57c10b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97c91d597bac157568a0191b7ce65b01e893dfa770b7d6d7e42784026efece2a39a58d0e607787886;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7116b671af4e4d58b8ee78b8af69323029deb5411957d2be29135d900450399d03da7eafcab93b9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e6be238b83b405ef2c580578982003393923ceac1dd8172b1c66513b42b76a62428ea1b4bcd6067d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77d797f188af74f7875087ab45e17fbb6ecaf58bc5ecf2670d9bda30f0cec00552237a2ba328ca225;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23b2ab18acf1f8250597969231dfe3307026e1a2098aad66c6e9a5519f438a24986734bd2a84528a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec5d179386a97f3cf63bc4a6effeeae42d4c5cfa7dd4395e399a206384a740a2ac487056d2f18af6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb48441dd2cf0d68f91275e1d81919db7c1e39ca3847e87ab8849f8a8a444c4a502618ca01982851ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h575897ea402c343cf3d27e10637badc67b7388e26c5ea4375bc0f28ab77b7edd3619adc238f172529;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d3660f6274c71357613d60984a594fda9f695bd460f3326cae23038e1f64ee38f59ae2c89e8d31ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27606a74af6a8ab6442ad8493849638807125033a8eec67fbfbcef5dd494efd309a0efb8130e76458;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8818ddb6afcffcdf872aa0407a897853bba3286fe1a2d4ce3d9c1752ea94c3202030af2c218461b03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42ddb2d45882100d1313a90c7133f47af7d40fbe0499648308711d4055c148a5f5a5f98350686d3b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59ef9b2cda7ecb6881b9b1fd731a4946d2d3275c4df98486fd187ae693daf7298e73f65da0ff473cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ec92bc373ce413783af3f87aaa664e5c52e24c34d91fe3db97681e6211dc6b81e86ee869e0fa5308;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dcb848b404d76d58a17c08c89c77a86f4d6491104b37ef53b74d547ab20d71411477fd73e540fbe5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2fcf85372e5e9caede348136b2086bf3bff4737129b8a398f69b31ef899cc453e843e535c4627216;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc527a9d838ad83fa549d4de0f7934d609ac2a1980435ecadcbec4fd8f86d9287f51437fc48ade3627;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb063cc4ab3c2a7bf9b5b43de144d67103a5c565946c03946a4479ad2111fb46443db0ee1a6fe16c84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb526b220df41220a05f988824482da7e43c094769207aabe940cb15377e3a25144b27dd17f0fd478;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39c775551b4937ec578ec06d1d919b1d2b3afe7a52b30458e13509e8e1318cf20682bf0a08707851c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6714a90ee959a49b64f9ee789f8e9c85f4fd280330a0f8c061665458ddc79584848cbfd2cf35c5475;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fe3d204f40eb9682c798438c4d6981ce14f70aa87f601a2d573029467237ae28bb94e87df7d5d064;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d28bffc27549e3a5cac950b44cd100fdad06c1550f77597372807ec5d14c8940d8f7dac041355235;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h417c7a1d74a0c5b20a2268ad5516d3656d71e07d7a0e154c6b70694fd3e19d6a01ece0019faeb4924;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedf8b67c73e78e354b138be91871ef05e6a7b375a8f314e37a3f5ae0fd5278fa40becf366e9a166d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25f12c02611d730fa01054cc589ce3a92b5bc3e3cff16cd93618eef94ca4360923d598cdee123460d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f932ca3bf5d441b4f6d6b07430541b4756c4eaae835395f9cbfcd4ddda4090385fa7cebcc5dc59c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a88f04f1af5b88466d59242b137be8290793bf2f75c82c4b79e5f38d4598fd0cbcfaeed1770b074e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h481f4bbbbce0b38730846227e05159d4937f3cca79766fa8de18d293c0837b8f0b9452f3bdcd5bfcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49f370b744e3d920e5d460ff03aedd74e5ac38af1590edce022dae9524abc7632455d7018cbd10d7b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h695245c5cd9a50b2edf9ecd606f2bbb5604cd2dba49e483a967210e90891561f8f269882965fb1778;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91dbf2d863ac2bfde72a217621df756c811db2f54be4a21f53e393307b954cb438b983ee5d088a16c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29e1e1b2f7e80de1ed6899beae4fafe141accb2377d12cd7c8e96802381e54ddeb57b9066636e568a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h400b16c5dd6a6f29cdd78f78585751c8aec54d76265227685aa447ad9fcc27c9dcae55a1062f2a1ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd8d633c105cb7944d78d0d795936d5769254ede8bf39c2106843b09c67fe0b1dd3a015e0873a400e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea30763d4fe8d616a8ff01d3b109838a354c40524c4d390fb7aebc55ac923fe0f59e4e08a541c46ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc89ec7cf7b8fd62067533a369648f1c483e5f5e3b452059830980aa4e60cffc806f4c8d5b4745b902;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb57061c3386f8dafc21aa57299a4d82aa8771e2b0ad3d78eed939f34ee2381cae0ab0656072a5039;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb83e53afafba3e9c63f91b53c8ff4db3b72a8427bdae0d297282410c93fa0c8683e5875e2b15b3744;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a8907ce0875973aa1900d9656c4226c62b61b30b85bac9486d48a50eb58fee9a1bc48ae9eaba64d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfb9f7f39af48085295fbb57fff76d5f1a604b33fc4a25d2d3bbcabacc9f0facdd8a213ac2d272191;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc8e7d0e6a2f3f4011255fed5da7085cb89cd6c846fadb085ed04c1197b95ea539f2d920a3f445145;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f627a96080d3dde941dd66eb923fd637096721b59176982f1e5a5c9be74f09bbe66f8ccdec14cb54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47ed20ddaacb52cb0c2608c56fc8012b72c60b4d0ac4401a09fbd13c7cd8928cc3b31f5c35727eaba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h626fd4b84a9f184f5b6fcb9327f26b192c5c13cc4baf23daa860bc7bb580554a7a5ff861245f32086;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c21715d346e27cde16eb3dbf01c23b8aa052c218c696ec18a22268ee09d8de55471eaecc4d1e8e04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0f5e228959545c6deda8a22317324eead146a4adffc4234319a15e0fa6070067a47c38ec2fc48f7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdaffeab4d5d0f82b028567a35a0f5b36617dff9bd485fef7b4eb22105368f886e906c4a9f3602d1e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1496f0379a79612d978b2b0395a2736d37d35061d2c212d56c6263e57c7f71c549f5cec90e08bf1cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h182e6fac14dec1a0cbc05466f91f9bb6c79c2acff298e4ce664ee82560dc0d3a28c06d21dd0f7ed6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f95ed6b96bb633163f052aa2ff53d646b9296f5bccffa771d1e85a345b734150592f15625c836887;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a9094f220256776ef246bcb0e1205f219e8dfc1f50c5696cebdc487bf35e7fd5452b198fc3bc3445;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f70fa14c9ac785439ac794e92eae9affd969478123577b1bb49bdcbf801886237f3c5336477fee81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c888b525ca099b02eeb801f3360a93de819c1328438c60c757588d13566f2d5a8dfa885fc74e0a03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2676944fd9a9a49cf1234357eff876df493271d6d0ec2cd8c0ad59ac0dd32c96675aec58bf9b8dff0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9022231cbf8726cb79427736eacd0ead9c2cc3b355b42abaaff8d260b3ac3216e20c8c9bef2efe05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2d979f45c153b0ca99de14d46f47e1350fd0d44f3cd3dceca961e242e5a8aeb4af1564b509785331;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfd5f58939c89753dd8ce6bfb4b516fda3eb06f814001c0bb55545374513d7acc6593286e3e147168;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf4e1d3d14b38a8acc46d65140f8f4f9546649a7c51954c3e9ed1898bc5d1c0b2f9fa41dfa0e36063;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceace939a1fd0d5adf67770f31f8b05cb510ae23dbaf4a0184c4b8a4bdafca7b29c024abc1e34c9f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2be0dd77e10b60f061572a87a8394e6cb6794ac41d78c43ee16d36cdd1927da22bf62f737ad8fc686;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8be432af89565c9cc2fd7784c6c9b0f425525f925703fa4d072030650e40fa843b74df48e9ca3ea3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3eeec726d796adf27f47444a70f15830c6626ced678a620f898677fbf0cab17676814cacfbfed3f37;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h715555c50d45ed4bd3ebfb2ce3d9d5fc09d45334df601ab52eceb0b6325cebed15dfb750ee0b06d03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90b8f7a29b360fde18e18b3c482ff76fa60b65d4260e9e18b0522fc812c2ee5f024c44ccbe6d65814;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a02ae4b1caeddc9c39f16839fb963c0934a7bc70adb0ebd7232dbb6e753cfa572ac22c1ea89bc2b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a40c5290bd992f2a004a7bd8b8523dcfb910118460d65b25ec84d7e7acd9c5770647b26a8f6cd8e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57a07136322fbd1c556bcb2c6e2556d4186c0cb54f35552f289e23f3f7f987a4acc6c6672534a8547;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca299c15f952d27d68a93d768ebaec29eb540f91d581c1daa7ba489e1bd792b3ead3e96c50209cb6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h837650276e5a69737578e37735ee94b369935f53fae65c8c3b4ba0ad1f48235a94557b39aecc188a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f1ec3e8b7ed67d22d7eb4b85a8a92db21db6b4297ca4894e58df323b7ea0261ff248abf02bec1b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbc24ba1b9b1967330083bcfc04dd4ca2d7bd076001399ad9257ce46678e14e3a2b20e1655abfc182;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8b04506cdac0720a2daf0190fb21ae36fccb00e45014701d790bdb6fdf1445df3b0ecf616dc79bab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf635082a6d006c4f9b85385ed9af82912cf92501db8f5740f3e3b103ba06659c7f697746b30be0d16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h291232d0a42475d819698bfc3b120c1bc57499ad55bf006b2848d5fdf26de2b2e20256ad7416ba6ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98e57b05fb6909a2a2c45da74ecbe2f1bbec70abe6a294dced350a837d88edaceec3302f6bf3ab6a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e07f0870ff9ebb3700df09e85b2e9bfccf8398f7ba3687b25ef1ddeeea0da9e542550b9ba8029caa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf27d8e3778f9904bf1268ad20a1f4fb83983470cbb2157e43710ab0e7057c62e65a7a25dc287742f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fd8d7452ede0571e80af2f86ad146483adf4be21dc597319d0f1ac6d1cad17ff10cfff56f35c5c1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5991a64c2a9ff7468d38173f1ff6f98931596c43e12ce3c45e2fb5576d9cb11083dee05df9341ba5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d53842ee757ae0d422c3100a2d6086bc460d12cadc6d87f2e008a59e96a94362df016353efe62ef3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16f510560de42d3fafc67c5691c1b69fcae7d559e13052d3204be8811e926d8fc47b0801882f379dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h328161ae329b58f49cff7293fbb7a9c7596b25780ae3c9918135d684e961899775fbeb41cef7b9e7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h137cd8fd6ef01888e13953c279a990ec8ed6e2350af6172f29ff4327148bd84385c0239d23207618;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee2866514b578b842bb52358b29bc36b344f142212e58fa90c4246599bdc361f09b1629e63677a665;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31cdc7a59852073f6f42f3da3c3d70e2b0fa05610430cc0dc66f2d63d9498920e15f12d8bdb5ea3b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae93437282b13855112f7b390d2470474a820d7a05a15fd906f14224e03e26a6a75d18e28a930dad4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h300696dd7787a1a0a56f52e0e304513fe2e440e771427dc500c3ce73a7bfe2f90b476232a35abd815;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha542152f98d5bf2d3005d26692d37f68432675e015ab20a3b20b83e71dd9eb306c5aceacc0569847f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc646bc088e72bbc87fcde4f70e66bb5bc108e8b307113e85578afc2d7e3090a8f360cd12a6c3fa39a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6363b0cd347329ac9520895965b0949461ab1e4fc6adc17eb42f53c14ff25dfa225aa952998be8d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebd3d0c5bc491861ed91c560b7278eef31f978116a72abfcc9df0b5bb258d2d6afc79086b29456cb5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb437966b2b15ebdac08982e058a5296881be39bfeccaf7acd1e773157a32babd55c9a1f7a45600679;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34402a282ef85b19d6faf86cca8cc9bf45f76905df17d3be2caa1b3d2c1f2575ec4143b3642a8c2b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had189c0bf3484b35b4be69955c3975753bf0edb2ca515c0f075820c7b234dcce0fdd864fcb744d7d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h889802895bcb947d25b81bf0dda302d385ed94149acb46bad34b9c2173e872b5c92e2e856402d44e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbd5429b6aae61e5968291ebe140092fda911abc4d18fbf2add9bd8ea9eb18d2b9c25549f13775f50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab64fbbdb1ed48c66efa18fd00fa39a66e83de8166ff014724e0caa5269a0e8b82a3c76cc07abb42e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea145e5a091810c944bc8ae500efacdf92cecf02589656860a0dbcd1266d7c3699dd1b0f37daa1a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49f225afc5949f4befbb7ef8738bd9c33e44328c1f3259276e5e42b03b46c08d21f601ce3ac1c1577;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35f8e88a8feaf8b8187f7528f1a680e7929a6ae0e39900f27648937ca031bcd9a0507d53416a96864;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4f62d053e49742b91fcc9514afa3a97e68932f57d5c405c4510c2b9c12e2fc73c7cc30f44916bce4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he59159a7480ee591be67590f9eb973487841ffa971dcc5023b7619015f45ade49351c7b881cc80518;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf099b1c474f2d45f98b437f1abee645e38c0f3fc8048bf423b360c1fa27bac0742f5901d7dbbc0ceb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19f1fc276642e50a41b5b8fa3dfdb0b76011fc433560c8ddb24c4dea8d6551aeb5a2dd79b2f3b235d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haafa12d43ef189d791b6059cb7ff6c09c1b8204b1649152386def1f4c2e5c0396fbb61a5d34ecec9b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6821124f2d5383f629965231933c7f3c757ec0b86286f946cf0e7a41dc55ff504107cdcc72db68c9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h952fb216d03d131e52fac401f652e9fbce4dc626b339703c0f99fc38fa0052cc994ea1b66d3b3e15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a5757fda7177641b4c5c090377ca51a1ccf95deda020f327f08eaf6f8ac94d0ee70017c92bad09e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2567050f197031bce97f00614f455fda22d9628fcdeb10b0bd984d28582803387c546d7ac3d755a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f5f0a60d2af370406905e8c370875d7efec29290540b841787a003b375f1ed5a30ea88a19c7770ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b855e0980583bc574cfcce0f1f3142f9694db6f6e7b437f0caac3762303981cf7e11338f38a3a00e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h687b745b3039408d9d63fdcdd8dbfb30449c9eaaf0ed13c253b5cbfb5d3cab13ccb4000b08e09aec6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h981bd55c0464aaa220c760a5f85ef2483ff3b963442d1de71c9848039b3b4b50b865d28174ff1f63d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h763896595b57c831eab017ee6ac7708bed2d9bbb8de088305104b34b96d8e2c3c1d92a9ccaf89b5aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7619343420029a08a27dc493191a8827367c5efdf320afa044ba357d9c3230e282622822d7ce41e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcedcff36c6ec5cec93e74c5caac3e72230ee90a2a4de1ddec0bb513a4eae3696f9183dee90b734b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4a71b7b860073f4b7019d9c3cdd300c4f52844137389ed9e6ea2f66d29e38162e3982c6373b4c73b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h935b1698e86ac1416e41ad35b4df8297a89d927d4122cc2c1a48dd33fd0b013b0b0bb91cb084bb297;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c769e092faeba8af055e8daa77052a523c63cd5fda5ab15e5d38864cbae51bc856577dda28c9879e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceb98230335adbe63ee7f155fcc535325f34ea56b8363e42b62b6b8465245cb084a49560e93051ba2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73611cb60c980325c3176ae97212f8c78b1d4d103dbbfbaf579dc4c8aa354807642a457071c611188;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ecef374a64cc1ffea0bf774a07d9cd96ae724732272c521f851b2828f43bd4bd83c98ca52dad72a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf479575350561a1ea3c0a0dc3a947b6fab5bbaf9f136e038af0059fa496befb6e0a02d459bb1e8c23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72caeefdaa0f6b972dbec4add136b9db4143247363a1fde557e609f6ee0ff3b3e1a1a8240133d0331;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1053acfdcc02cacf54607f187921bd8e9d0ed36bc1cf7c9bf6b0c8a31bf74a38e84308e2cb7d91726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecccd8213eee3505756016db06aebbb1e21246395f0cc3909ecaf84fdbcde0a392f270719b4f469a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a5493c83a32b4c97f1ade5d1ce103d75af8dba642787708274a51475fe7e4d528b3f1f9ea0351e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15807cd27d266af5ea9ee655021a993fa1a3b2bbd7621f2b2213f22ad5df8b03660fa4943b7255e82;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443ae3de65d48177e56ec6522abd656e71347540d8f1cdadaba714015ba50f4d0793c5ef9a7e03e24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20654919d815a74bdb09e8e4102253d6cefe08301d9fa98fb700fd3c161e43c1aa7a6b2fa169c59dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha690b3e4170261d112208dc8cf3744df8dead1b1723657c753467226120b9c6e5515d60e980da06cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h480403de7ddbd900293c7feb81cfa6a4ff08b2ffa8bf3ed46e1d8c43deb912802e9a3c3bdbe2ae0d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0bc2dca6355d4912b21fc89afc0edf873416c0693c69a30c638d277ededa724418f1c24630ec4718;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74fa00fcd6bdb94be99ec60c2d8e0e03ab9f70c25e6b8fc6afa252ce2e10c71be09a6c52045b4aeb5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc187417f7429cff37be2c85612af1841f154ab45f5e4d90354347186df7aadcd5c2f9244df3ba6869;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9435246bc76de6390bf34c6ecd272b7dcedc02a2245c9d141624755ac3bd55017cdc6ddaeed7fe3f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h178c0b7c518a67f3875409e7060ecc9bef597d361f3f5b04ce975dc6774fb9eceaff80415dfe992de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h929f20ac5448819f5998458eb8373b317839ee7f3e282e8fb85f1c043b1bd464af5449c167b08252f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h627f249dce433d1a0e1718a1564390041f9054af8f8133fd871c3b29eba3c134c2b23aca12fddddf1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5bfbb9d3bc34680e66614ce8f0c383d00727db7ce7b5f87239481a2b5e7819a19b3c2d1af1a8bf8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda909a129650c80d4f880f6e2f6c2ead2f48817fa5a0077f1363167a35b6b113f44b64a650ecc6211;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed641515004cf9a3275446e185742f8055ce003aba4acd0a3f2e5fce39171d636722f73b8f4b49c8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aa499f6a359c3d62c6d459814437bab70f343aa381a737806912f3190af58cb29250003178bf063a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h543e1c0fc18634ee9da3992ecad0a447e6a4c8a1e619e9f07a40a7ebd3053194878849ba17498148e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94d38c92badf4a46854848f1356d44ca56d8758fcd4a0ecfeff4639062717c3c5196bce53f1d68a14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5a90c06508288995bdf97c7043c6128b6540e773b3da7733531e2b7af640a166147464496195bc98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4b6c911f230716b2151192f1ef8db703166faf954d3911115dc8389c821cb0ef646eb397a186b0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h525dc682552872dd6e1d94138d0bdd9ad9d8aa720327e9dccd69e390429d605e665302bcd8578daf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe297d130a6e88aa1c13161d93d30e13b5447d59faa2900bf78abd021e1a46c6a0b31a2d58613cb85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h467e89fc14379488e07e196a23657dc67794c27ec195873a6c021cf0f8bce78c2b48dd95d25787c0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h902e36addc498cfcce97642b5eeda08ab3b20a7a2e1174882fe971162b3a5fead624e53c462f99cd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21241d649319f1472739fe529534258f6e1d360da875115c6941aeebf730079473fe923856b42953a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6aeffe3a8060ba3e3f9fa35f121d8acc64147b7e0b7c437007456ae893c091e5b1927e633553a27e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42a62998af5a10a80f8ce31d78e7766e34c7ff3c1034b80a986a73d49930de18f3d23e7a614e0cbd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdc266f3ec7dacc1ae40db10fcca6bb30a030bdd199e982bc90b0e51f34e6dbd799f1f61f512b087e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf3f74b435946b4826d83edef3101a289d90efa75f96b52ed0c10283abbe2f4a3c3ecffe3efbac54e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h855e2a37f275141c93395bae55c0379e4437cbd7ce8c6697b5f5164a3cfe95063f889e0d1a801ea18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h648709ea79eca656293ee39c902df02b1710557cdedea5719a05f33aa4868029b90b69a3254ac18ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65e04c440382eb7dbd53d564921dbd48cc26541ed55b1c9031f11b42ff078368fc5874394e39ccce5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45ad5a8765b178449274a8d602da5fc652f440baf964891fdd6f97f3ff311f25352267a45b8d6b5a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haed5c3b64f75bfd8b17a3c904b8cd2e8e088904168cbb19d4b5832008bd462e0445afafbde8a6ba50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd60b516d96401ba676e871d54485d963913ec67313e3919cbd11494cbe3006bdeb59c295386ccf22a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h640520c3d1928c958b0bf9166dedf6d312d48442d27f801264aa3884b38e8b85ca799f06c4d7a480c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8197b036a9b4d5fcf4f9beaaf7eb13d8a083c92f0b4327ff4a1122a11a6a2cd492da53d8cc7fb1894;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1aa9f7b9ef1e2a5d62b5842fc16fe2849a24e19b5559d76aa3ab28180c90b110328a7c099c7a3afa6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf24a3dae820c1b2721813d661a9ec5e93e159a995967d44d6883bc851da075ca1293d4f19d9e39616;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd720f2726a4775942cc9bd6ac6608194a817ef07c025a45a4b39a465411d59c93d85324ab98c493f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd767fc69fd05b73adc659f220e461a20578c574b8314cb91137d25e12f1d1aeb0d16cf48b1f56e00e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8760e312c93977968a7ca9d20cf3fc797e290e827d5df6290cde38286d7cd32f29de865bd9a38b13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4a7ec5c3f6863fca468ab27f646dd15df60402f417619ad55e0435801514b08fd1ef00467d5f8f90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b2be255a4934aee0f2155d5e9d211fc78900e2351a173ffa8b76e584c71585b801e8834feb89a4af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h366cdaeb1bf10fd6d89314e9ddef42abd172800816fb075c1fde3e382d98a731cf230e92492825e06;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6bcfb8b6939c9b6eefd372a9e12dcc2d4e13f6795e2c1046e522d60238d6cf88fa0b5c4ad040ae59;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee48497a638886dba439fd32fac183dc012a63e20779c7cbeac13f42eba118363ba0511720426b19f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e23608e4d2706ad1ca69d7c98ad3602d13bdc92e885b31321ed737c81af00adbde61d07edd6fb684;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58e827a6f551d8545bc9593cab9f7f4a1704778dcabdd975ac4ca0d73a039e459f137fd386bfeeb66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd158b9a51710cf38d9919b6d5c17992c31591d48d9bc3b5a46ea1496138c8f78189a0f0c5baea9365;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4403b275b12d9c0fd4be9af3bfdc6d44f577eea38ce1dcd918318d8e0c237daa6e67ccb93d7a7eab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dea08028183398aaa194d9d30f97db5c601f9891129cf1a2f88308b6f9aec1b06ceb45bf69ffbb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbc5b9e817f65795f8d0a2e54bb0c07039182555997f1904bf6513e0b9e6ec7c8eda3f22501ba8fa1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha97d46075fa7abb6f5749132bd325d821b1a0f3c258cc3a7e4f0d889faf34012f89ef5cdcfd55bdb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3805c65a3ce7e7c1168539c2a84c64e0f92cde972502892a4dfdb802773568fa75adc0ded0b9cc0a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3316955df76490eb7977e910ff05605db2a9cbc79fee0c0a993de8e07ae239ce8575ba76a2dc8ae92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cfa1fda6f84838d5d1b5db203f9b1b7f5be118baef42e1998a4af0adeaca9024276444cf093b093d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4db2feec64e05c699425609360677d4df91c08a501e33a8aa936ba5f81b57b377af98b44f73bd33cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha45502bf074be8058590b658b78708c74a2efcb0e7bfbf3c6d6731749372fc9c98fd1065cc247e217;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10cca639f15c924c3790d0b0548f77bbd0a7f5d2d5d516a5b237c5082fca3a66a01b85cc4f7bbf957;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68ed5c21943eaaf3fb77ba78d4681d35098eee9a6d98ff6c938e15c02debe3d72dbef09137740d3ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee6e4ed43397e0e4a961fa1a653e7fb14aeeb94f5ea1a356d7a1b53ddbc49f886a503d8a3c4b4bcd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59df84831a1059af7307cd7a349b78a91270fa9c1d9d8a0ee18fc27bc2c139cf6c5f3c41f1b0e53d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75aeb1f3e77dc619cb003f1de1850a6c03e4bf320b522a9d501c83d4129b30483f999efdfe626e46c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h366325b37a424a08538da902c511f8cdc44a1fd40b70f966178fd6230c1a827732e9174a6aae8736a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e856ea7af4df9f859b82115a29f128f9f4ce6ed753077710fc9ed4a7a7fa5e7ea2240b6fd0083019;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dc0bc48bd27e5f684ee87c412abf7f1a6c52fdb86eda30e5aa81b31a9f5b2ae0b8a1a3d77ab34fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e95259bf9e0734fe0e7afc739aa922909d5a31cdd40835b506591e31d5e18cf95039f8ec4be8c5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c1de0c17fa6b4f5a85af01896761dfa07bba492d995c3c48b9426a632042683477a896b49625f848;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd1e5dc6edbed9c601a3cc73dd052815a28f7f548a6989008fc8d864d76a84777f261580768f6f0a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecd53ec850ae0b9e181c8bff4501e8da86d693a5d7b9dcd45494dbe8e14cfd34fb95c2979740395ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7520bccf77508851fffc12b098d95bc17cc614802d35c1ae3753ff49753f8d43015c36b50f7f902b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccf4eaee93f55a6406ce55f44b2c0294f83db13ac72fbb44f71c8bf14053dc696e7eefcffa14fbee9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74796bcc120d2e21c5e3ad023908c44be674a3c80ad7b42c3deda866581bb72ae2d9d3b6a9f3c51c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h488ff2dd37a49010c6c48a825ad8fae7d13d445c69158e4a71b7b5c8f763d646c577f34ee3c604633;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd98bb469a37885a6da6f852ace0517dfc51325ce47dfad4262e26dc1338974fcadff781f5ecdd471;
        #1
        $finish();
    end
endmodule
