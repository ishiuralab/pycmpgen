module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    compressor_CLA32_16 compressor_CLA32_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA32_16(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [14:0] stage1_0;
   wire [9:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [14:0] stage1_4;
   wire [16:0] stage1_5;
   wire [18:0] stage1_6;
   wire [11:0] stage1_7;
   wire [13:0] stage1_8;
   wire [14:0] stage1_9;
   wire [12:0] stage1_10;
   wire [10:0] stage1_11;
   wire [15:0] stage1_12;
   wire [17:0] stage1_13;
   wire [16:0] stage1_14;
   wire [10:0] stage1_15;
   wire [8:0] stage1_16;
   wire [4:0] stage1_17;
   wire [4:0] stage2_0;
   wire [11:0] stage2_1;
   wire [1:0] stage2_2;
   wire [9:0] stage2_3;
   wire [6:0] stage2_4;
   wire [8:0] stage2_5;
   wire [5:0] stage2_6;
   wire [6:0] stage2_7;
   wire [6:0] stage2_8;
   wire [7:0] stage2_9;
   wire [5:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [15:0] stage2_14;
   wire [3:0] stage2_15;
   wire [11:0] stage2_16;
   wire [6:0] stage2_17;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [4:0] stage3_5;
   wire [1:0] stage3_6;
   wire [4:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [1:0] stage3_10;
   wire [2:0] stage3_11;
   wire [4:0] stage3_12;
   wire [1:0] stage3_13;
   wire [6:0] stage3_14;
   wire [4:0] stage3_15;
   wire [2:0] stage3_16;
   wire [7:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[4],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_3[25]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[5],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[6],stage1_4[10],stage1_3[10]}
   );
   gpc606_5 gpc11 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[7],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[8],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[9],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[10]}
   );
   gpc606_5 gpc15 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[11]}
   );
   gpc606_5 gpc16 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[12]}
   );
   gpc615_5 gpc17 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28]},
      {stage0_6[18]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[13]}
   );
   gpc615_5 gpc18 (
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_7[24]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[7],stage1_7[8],stage1_6[10]}
   );
   gpc615_5 gpc19 (
      {stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage0_8[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[8],stage1_7[9]}
   );
   gpc1406_5 gpc20 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[9]}
   );
   gpc606_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[10]}
   );
   gpc606_5 gpc22 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[11]}
   );
   gpc606_5 gpc23 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[3],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[12]}
   );
   gpc606_5 gpc24 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[4],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc615_5 gpc25 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16]},
      {stage0_10[22]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[5],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc615_5 gpc26 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_10[23]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[6],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc27 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_10[24]},
      {stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage1_13[3],stage1_12[7],stage1_11[8],stage1_10[9],stage1_9[13]}
   );
   gpc615_5 gpc28 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_10[25]},
      {stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30]},
      {stage1_13[4],stage1_12[8],stage1_11[9],stage1_10[10],stage1_9[14]}
   );
   gpc615_5 gpc29 (
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_11[31]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[9],stage1_11[10],stage1_10[11]}
   );
   gpc606_5 gpc30 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[1],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc31 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[2],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[3],stage1_13[8],stage1_12[12]}
   );
   gpc606_5 gpc33 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[4],stage1_13[9],stage1_12[13]}
   );
   gpc606_5 gpc34 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[4],stage1_14[5],stage1_13[10]}
   );
   gpc606_5 gpc35 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[5],stage1_14[6],stage1_13[11]}
   );
   gpc606_5 gpc36 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[6],stage1_14[7],stage1_13[12]}
   );
   gpc606_5 gpc37 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[7],stage1_14[8],stage1_13[13]}
   );
   gpc615_5 gpc38 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_14[24]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[8],stage1_15[8],stage1_14[9],stage1_13[14]}
   );
   gpc1_1 gpc39 (
      {stage0_0[21]},
      {stage1_0[4]}
   );
   gpc1_1 gpc40 (
      {stage0_0[22]},
      {stage1_0[5]}
   );
   gpc1_1 gpc41 (
      {stage0_0[23]},
      {stage1_0[6]}
   );
   gpc1_1 gpc42 (
      {stage0_0[24]},
      {stage1_0[7]}
   );
   gpc1_1 gpc43 (
      {stage0_0[25]},
      {stage1_0[8]}
   );
   gpc1_1 gpc44 (
      {stage0_0[26]},
      {stage1_0[9]}
   );
   gpc1_1 gpc45 (
      {stage0_0[27]},
      {stage1_0[10]}
   );
   gpc1_1 gpc46 (
      {stage0_0[28]},
      {stage1_0[11]}
   );
   gpc1_1 gpc47 (
      {stage0_0[29]},
      {stage1_0[12]}
   );
   gpc1_1 gpc48 (
      {stage0_0[30]},
      {stage1_0[13]}
   );
   gpc1_1 gpc49 (
      {stage0_0[31]},
      {stage1_0[14]}
   );
   gpc1_1 gpc50 (
      {stage0_1[30]},
      {stage1_1[8]}
   );
   gpc1_1 gpc51 (
      {stage0_1[31]},
      {stage1_1[9]}
   );
   gpc1_1 gpc52 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc53 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc54 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc55 (
      {stage0_4[31]},
      {stage1_4[14]}
   );
   gpc1_1 gpc56 (
      {stage0_5[29]},
      {stage1_5[14]}
   );
   gpc1_1 gpc57 (
      {stage0_5[30]},
      {stage1_5[15]}
   );
   gpc1_1 gpc58 (
      {stage0_5[31]},
      {stage1_5[16]}
   );
   gpc1_1 gpc59 (
      {stage0_6[24]},
      {stage1_6[11]}
   );
   gpc1_1 gpc60 (
      {stage0_6[25]},
      {stage1_6[12]}
   );
   gpc1_1 gpc61 (
      {stage0_6[26]},
      {stage1_6[13]}
   );
   gpc1_1 gpc62 (
      {stage0_6[27]},
      {stage1_6[14]}
   );
   gpc1_1 gpc63 (
      {stage0_6[28]},
      {stage1_6[15]}
   );
   gpc1_1 gpc64 (
      {stage0_6[29]},
      {stage1_6[16]}
   );
   gpc1_1 gpc65 (
      {stage0_6[30]},
      {stage1_6[17]}
   );
   gpc1_1 gpc66 (
      {stage0_6[31]},
      {stage1_6[18]}
   );
   gpc1_1 gpc67 (
      {stage0_7[30]},
      {stage1_7[10]}
   );
   gpc1_1 gpc68 (
      {stage0_7[31]},
      {stage1_7[11]}
   );
   gpc1_1 gpc69 (
      {stage0_8[31]},
      {stage1_8[13]}
   );
   gpc1_1 gpc70 (
      {stage0_10[31]},
      {stage1_10[12]}
   );
   gpc1_1 gpc71 (
      {stage0_12[30]},
      {stage1_12[14]}
   );
   gpc1_1 gpc72 (
      {stage0_12[31]},
      {stage1_12[15]}
   );
   gpc1_1 gpc73 (
      {stage0_13[29]},
      {stage1_13[15]}
   );
   gpc1_1 gpc74 (
      {stage0_13[30]},
      {stage1_13[16]}
   );
   gpc1_1 gpc75 (
      {stage0_13[31]},
      {stage1_13[17]}
   );
   gpc1_1 gpc76 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc77 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc78 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc79 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc80 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc81 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc82 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc83 (
      {stage0_15[30]},
      {stage1_15[9]}
   );
   gpc1_1 gpc84 (
      {stage0_15[31]},
      {stage1_15[10]}
   );
   gpc606_5 gpc85 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc86 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc87 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc606_5 gpc88 (
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc89 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc90 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[3],stage2_6[3],stage2_5[3]}
   );
   gpc606_5 gpc91 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[3],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc92 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[6]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[1],stage2_9[2],stage2_8[4],stage2_7[5]}
   );
   gpc606_5 gpc93 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[2],stage2_9[3],stage2_8[5]}
   );
   gpc606_5 gpc94 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[2],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc95 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[3],stage2_10[4]}
   );
   gpc615_5 gpc96 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[4]}
   );
   gpc606_5 gpc97 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4]}
   );
   gpc606_5 gpc98 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[4]}
   );
   gpc606_5 gpc99 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], 1'b0},
      {stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[5]}
   );
   gpc1_1 gpc100 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc104 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc105 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc106 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc107 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc108 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc109 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc110 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc111 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc112 (
      {stage1_1[9]},
      {stage2_1[11]}
   );
   gpc1_1 gpc113 (
      {stage1_3[5]},
      {stage2_3[3]}
   );
   gpc1_1 gpc114 (
      {stage1_3[6]},
      {stage2_3[4]}
   );
   gpc1_1 gpc115 (
      {stage1_3[7]},
      {stage2_3[5]}
   );
   gpc1_1 gpc116 (
      {stage1_3[8]},
      {stage2_3[6]}
   );
   gpc1_1 gpc117 (
      {stage1_3[9]},
      {stage2_3[7]}
   );
   gpc1_1 gpc118 (
      {stage1_3[10]},
      {stage2_3[8]}
   );
   gpc1_1 gpc119 (
      {stage1_3[11]},
      {stage2_3[9]}
   );
   gpc1_1 gpc120 (
      {stage1_4[13]},
      {stage2_4[5]}
   );
   gpc1_1 gpc121 (
      {stage1_4[14]},
      {stage2_4[6]}
   );
   gpc1_1 gpc122 (
      {stage1_5[12]},
      {stage2_5[4]}
   );
   gpc1_1 gpc123 (
      {stage1_5[13]},
      {stage2_5[5]}
   );
   gpc1_1 gpc124 (
      {stage1_5[14]},
      {stage2_5[6]}
   );
   gpc1_1 gpc125 (
      {stage1_5[15]},
      {stage2_5[7]}
   );
   gpc1_1 gpc126 (
      {stage1_5[16]},
      {stage2_5[8]}
   );
   gpc1_1 gpc127 (
      {stage1_6[18]},
      {stage2_6[5]}
   );
   gpc1_1 gpc128 (
      {stage1_7[11]},
      {stage2_7[6]}
   );
   gpc1_1 gpc129 (
      {stage1_8[13]},
      {stage2_8[6]}
   );
   gpc1_1 gpc130 (
      {stage1_9[12]},
      {stage2_9[5]}
   );
   gpc1_1 gpc131 (
      {stage1_9[13]},
      {stage2_9[6]}
   );
   gpc1_1 gpc132 (
      {stage1_9[14]},
      {stage2_9[7]}
   );
   gpc1_1 gpc133 (
      {stage1_10[12]},
      {stage2_10[5]}
   );
   gpc1_1 gpc134 (
      {stage1_12[13]},
      {stage2_12[5]}
   );
   gpc1_1 gpc135 (
      {stage1_12[14]},
      {stage2_12[6]}
   );
   gpc1_1 gpc136 (
      {stage1_12[15]},
      {stage2_12[7]}
   );
   gpc1_1 gpc137 (
      {stage1_14[6]},
      {stage2_14[5]}
   );
   gpc1_1 gpc138 (
      {stage1_14[7]},
      {stage2_14[6]}
   );
   gpc1_1 gpc139 (
      {stage1_14[8]},
      {stage2_14[7]}
   );
   gpc1_1 gpc140 (
      {stage1_14[9]},
      {stage2_14[8]}
   );
   gpc1_1 gpc141 (
      {stage1_14[10]},
      {stage2_14[9]}
   );
   gpc1_1 gpc142 (
      {stage1_14[11]},
      {stage2_14[10]}
   );
   gpc1_1 gpc143 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc144 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc145 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc146 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc147 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc148 (
      {stage1_16[0]},
      {stage2_16[3]}
   );
   gpc1_1 gpc149 (
      {stage1_16[1]},
      {stage2_16[4]}
   );
   gpc1_1 gpc150 (
      {stage1_16[2]},
      {stage2_16[5]}
   );
   gpc1_1 gpc151 (
      {stage1_16[3]},
      {stage2_16[6]}
   );
   gpc1_1 gpc152 (
      {stage1_16[4]},
      {stage2_16[7]}
   );
   gpc1_1 gpc153 (
      {stage1_16[5]},
      {stage2_16[8]}
   );
   gpc1_1 gpc154 (
      {stage1_16[6]},
      {stage2_16[9]}
   );
   gpc1_1 gpc155 (
      {stage1_16[7]},
      {stage2_16[10]}
   );
   gpc1_1 gpc156 (
      {stage1_16[8]},
      {stage2_16[11]}
   );
   gpc1_1 gpc157 (
      {stage1_17[0]},
      {stage2_17[2]}
   );
   gpc1_1 gpc158 (
      {stage1_17[1]},
      {stage2_17[3]}
   );
   gpc1_1 gpc159 (
      {stage1_17[2]},
      {stage2_17[4]}
   );
   gpc1_1 gpc160 (
      {stage1_17[3]},
      {stage2_17[5]}
   );
   gpc1_1 gpc161 (
      {stage1_17[4]},
      {stage2_17[6]}
   );
   gpc1163_5 gpc162 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc163 (
      {stage2_0[3], stage2_0[4], 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc164 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2]}
   );
   gpc606_5 gpc165 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc615_5 gpc166 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[2]}
   );
   gpc615_5 gpc167 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc168 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], 1'b0},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[2]}
   );
   gpc606_5 gpc169 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[2]}
   );
   gpc606_5 gpc170 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[2],stage3_14[2]}
   );
   gpc1163_5 gpc171 (
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage2_17[0]},
      {1'b0},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[3]}
   );
   gpc1_1 gpc172 (
      {stage2_3[7]},
      {stage3_3[3]}
   );
   gpc1_1 gpc173 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc174 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc175 (
      {stage2_5[6]},
      {stage3_5[2]}
   );
   gpc1_1 gpc176 (
      {stage2_5[7]},
      {stage3_5[3]}
   );
   gpc1_1 gpc177 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc178 (
      {stage2_7[5]},
      {stage3_7[3]}
   );
   gpc1_1 gpc179 (
      {stage2_7[6]},
      {stage3_7[4]}
   );
   gpc1_1 gpc180 (
      {stage2_8[6]},
      {stage3_8[3]}
   );
   gpc1_1 gpc181 (
      {stage2_9[7]},
      {stage3_9[2]}
   );
   gpc1_1 gpc182 (
      {stage2_12[6]},
      {stage3_12[3]}
   );
   gpc1_1 gpc183 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc184 (
      {stage2_14[12]},
      {stage3_14[3]}
   );
   gpc1_1 gpc185 (
      {stage2_14[13]},
      {stage3_14[4]}
   );
   gpc1_1 gpc186 (
      {stage2_14[14]},
      {stage3_14[5]}
   );
   gpc1_1 gpc187 (
      {stage2_14[15]},
      {stage3_14[6]}
   );
   gpc1_1 gpc188 (
      {stage2_15[3]},
      {stage3_15[4]}
   );
   gpc1_1 gpc189 (
      {stage2_17[1]},
      {stage3_17[2]}
   );
   gpc1_1 gpc190 (
      {stage2_17[2]},
      {stage3_17[3]}
   );
   gpc1_1 gpc191 (
      {stage2_17[3]},
      {stage3_17[4]}
   );
   gpc1_1 gpc192 (
      {stage2_17[4]},
      {stage3_17[5]}
   );
   gpc1_1 gpc193 (
      {stage2_17[5]},
      {stage3_17[6]}
   );
   gpc1_1 gpc194 (
      {stage2_17[6]},
      {stage3_17[7]}
   );
   gpc2135_5 gpc195 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc606_5 gpc196 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], 1'b0, 1'b0},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], 1'b0},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc2135_5 gpc197 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], 1'b0},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc615_5 gpc198 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc2135_5 gpc199 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc117_4 gpc200 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc201 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc202 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc203 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc204 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc205 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc206 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc207 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc208 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc209 (
      {stage3_10[1]},
      {stage4_10[1]}
   );
   gpc1_1 gpc210 (
      {stage3_11[2]},
      {stage4_11[1]}
   );
   gpc1_1 gpc211 (
      {stage3_13[1]},
      {stage4_13[1]}
   );
   gpc1_1 gpc212 (
      {stage3_14[6]},
      {stage4_14[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor_CLA32_16 compressor_CLA32_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8f213b1e749ad8503a67b856442bdb04c3766f8415f1e738a5d4b9d01a96fe73fd2f87d38ae8c8b04b06c92aece2517ec1bfd36ab3fb45c90c2cc4e97728416;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h78117f8e139e65be82ddcf2aa88f5d6393b81e24e6faaaacc33be45ca03fef8f0357b87a9e1224ae583c346eb1919df1984cb7608c19e7d83887d075049e1e38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h34a6780a1a88536fe5a2b06d1d8ab2b03d0c5ccaabc32dc1dfe83bf597570f279e82135d7f899f20ce145406e42d8cc2f2cf6cd0511f99c96714746925b964c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha4c820414feaa5b679eb77fbd51fcf6ef8da3f0e4f6072071a72902d2572c4a6ab4efc900f7383d440cb11823e62354df9b087ef8e656d61cf98651cd32171c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h87285b5160de7c0e0d6c9375d3c380226559ffa51a88bdc186a7db621f51681e607e778cbeb1fb08d60924df363c0d4fd35bee7828ea83a19f806699d7cc257e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6953b0f2a7e903e1459a708ca2c8f8e9a4a72c93f3cdfe2d4a97131e4ace7c4811399e3ccd0cd68a479fbc72d3f59fee633ab436e26a722382a521744cbd4fcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h364c25cb7933831a5b1216fa93838022b4045b6112cbb94fd545c37baecbcfa7e11982f28fbf4519ff77d3e0007079c1d35e7b999044f5e94a4cf7753c641b26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfd3616bce56df7e4a6a03863cf1e973da46eda5c983e620162e72a1c04accac9c86f2a6d711eb82aa39e000a889c3709744d1efa567222ee11bfa75ce0db2f1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h52a9610f4719706be36bde88bb3a16b899dc30d8a2b11f72a143718be197b8766e1bafe5758a8afaa12ecedd626a163a21a01beaa8440bbfb13862d5a65a3d2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7a7a40a798ba16280507402547da091ea8d12a89602f27eab7bb1a5703603ca86412120cd946bc8c3eb0c85bebf190484716c5f23ee565c9f65cf6972c436274;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he60e5ff322ee0ccdb8ae459d59fa6acb4d35fb7c7167e3240f94baf55735fe379bc7bfa37b2ae9bdc1ec3ac8c0e042a2412c522169edfb58c55ed76257dbb183;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7d5cdcdb792d48de2f18a1ecf5e68e142db7b3765f4ac7e104669d65217fd998e2aba1a79292ccb28b23187f51faf6f19eff5f4a41629f126d8e3394483a1b3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf703b92ac0008cffe6daf248f2bc2c41cf07b3ada918066cec04e9494e803245a4c19df796385abf3e7c2468c305414791fdf9bd509970d945d71e773d50cfef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hde240e12e4b83749747dc13c6e57b7331348c38f3356d03c253ee99bd946780436db13e11d06b949e8e0c7d161d08625ea26c7c5e5d2a2b28d9f6ffc37ac7ea3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h705674bff4a8cb8ee0ba978f794cc3b12bea7a7518c37a61cc6f701c1a90af67bee61967d4cf9d7ac135158448db2867cec6bcb619170e179bcd725be7fafc88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h560701a6ffbed4e370c0bfb382705220cd03ab3554af3ba86a6999330a6afaf387e50727f59b810625fb88e03a1b186ccfbae4250d144dbda1f08d9254c68fbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1d87536e998fa6be5848043157ec43f294ee841a4e725f5fb4b539ce9b97c0c25a2bd2ef7a955229ca0a71359a295417f79b0f709c16e50f40afd57740c04d98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hec882c0377980054b93c97a69460177d77c4b4b10747edc4758f2210bd1e0e4270e030fe47f0798ec893b8a60eed0dbbf2b81b19d12af1e71ba6e7ae8aaa6c90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he2d77abe73841803e209bf1037b49325ef85113727e2bf5518e7fe9cfa895b5940f55fbff2b0298cbb141b5809301ff1cc07c7147159f04b2be1552b456fd873;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6047255067960a039f31861b7fc9bb947a18985258707b1a73237d1ede56687dbc7020dcf9fc389b25b84036e6e541b429aafe6fe35b6dae5ac03bc0bdcc10eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4bb53f1519827caa4586cebe72f42f2f0a0076b0537ce0d924a1a09fba1126d169196780b1725d850dddba16bcee9be2e38f2cf11672b4172d154fcff646f2ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd2788240e7c17007fc5f1048f8fa20e0a5ccb212859e0628387eaa3191d50e3337336c284357d9c6d250c07a8b50923ee966d77d6db2e244f124343c43232952;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hae91a642ea35f6f853ff641be1f5f749b7913df75eb91030ce27f4afe25be1e2409f7de085e51dfef31e12a950fb2ac3db73ded97e8cabe33cf76af7f94a14e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h32a392efe9384c988177437fe6342ad770b481cfdb7f330ae635a31786e23d48c99e6464720f9d23117f345972f93e5cc460c5411e8bc5c3880ba82e10521053;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h39090f51ed425a6fd3e2adfd3cd8f5e0005a98de94836d461b375b8ee41dee11805b46ee8f40a2ac2e26367e088df04e06ae971832e1441eeffbfed743032f5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hba29f26a3009ce0552ee5cb86df01779c14e387edce01369004bd4e907f2cb61aa1dbc79d9f91e5b6de4a25b4cde1d570e53de757c6a72315f2cb868dd89c68a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5ae1bbbf493fdc44c0511dfe7edce1a1c918e70d27b6dbc8a382dcc98cba3834f6841d4e9a422ea06dd57e4d02e20fd9330ea9b36e9df91dde06cd54737a0953;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6aeeb0b128000080a7bed28a8c633f8b4a78295262d30f519e0ed5a7bab678d92771b764075d67fddec11ac5e7833178cce4e565f19b501bd4a06189d143cb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc42f36390d6e9ea915579ffb95d1973a2cf82a04f7bdf766300d1dfe437d57b692eb0d89f858c8ee21e0c5f5d1733a235fc728606f9ad9484e0cb1aa4ca9d925;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4ae46a76620ad24ba1f554766748cad84e7b16e2cfbc55921df3a42900e816cc5214e84b8eeb3e302dbb91a156bb8ab14c4408f84149628ec9e16d8194bd6512;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4a0b39b6ea87207c120b8e3c9ab1f3b757cf0d4817265c0d12187613d629f5136a71c377c1a794169b2de1c419e2dce674ac38c3168e0aeb73daa26a189d3f07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc870671cffff895436b6df3606ad2d7ff090013602b434b6d2592846f43bca6514e74d466040aac970b4479499fb33b6b40685e2e263b702660d7e612ce5e2a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd27ab93aafd1328d2c7e7af86378bfc8e7b70ce4616a4e526b8590b036553011de7bb421aeeddc958c5113a2c63bfdee996b68cd1d62b92941b3a62be52d473;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h39a512ab77a9c0ad3ea5eb9e67abc104651cc69f3c3a2266d438becfa04b99c69f0a1b5d011f582a0057d0de763a16178e45b5a35d154a804bec279f0bebbb9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h821c758da62b1436b32ff07701e28de818d8ef4433cd0890b3171e9ec9e7ea310b8361d4632990e24931fe3af5968d5675f31c1a74a32a46aa0308251b45a1a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h73248e1d8c232120df8fc660200b50f6d01d8fb603fdfa7c29781baf1a7d548dc79f41acf3da85c24845659d00949daeb27d7f3d7a707afbcdaeae31ea6a3cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd1db01f445d90d839c00ddc9a26dce38aabe1cf429ef407c668fb4d34bfb027b58ea983e4a9472ea267c349abfccc3c572b3b433147a656adf6ddc762402e265;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1765caff53a9c14b47ca436bc604bba2d94f109e2249077e51be4b0dfc1ddeff4dfcc34d264fd61d8238ede6e531f0c678edab44d24e27f6936cb9b82aa6ccd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5e22e181d5b9d891891568868ec8263905698875d094f4ad39562de7f2264904afb34afb275adc3cb2548febea281cc08fddafeb877c6a25d0fcd0ebee8a85f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haaa826b37e5f45a45dbac6bfbb8cc12c22070fcecbc33c4c3daab66139d3600b30ea28ecf13e0e5a7e673f2f113b40bea3ae0934f0c5c7a9a726ed6c66c5a98f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h49cb4daedc9a350b4b973baf82a7ef0a5194a247dc1da13f202cf0d6578ab11c7e831de207fe573809401ca78f426f0b575318010af0f6886d23ebbf7d2332e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hab6240fbdb83d1418d31efcb5c27c09f76ecd71f43aa6595dde8896f9996ca71105da7c00f880e0dde4b33f27d2ef7e1a3a61975be70d742cca7ddfc5a40d034;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h16ce1c69ba79242c24339f8758843f07b3244c0897e6d713e0df9576f61e8242d8528716713447153e571c6257de46fb27576934d316650d71c905f505b941e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf6151538d9c79569ac773a9bc3e8d669fb86aa8585b4c7073b6efc5fca9fefd45e59b90a6afac4d71f931e1379d6b46a7b072530641da9fcfe7dd465c63b2a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h46fe65f9afa57beb9bd71d1b32ec15e873544fb29eefdb0a81741f998c1e678dd9cf984d8e6271b5ef130c12e1229b42324daa6fbc7308520a56c276b18a300;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha7ddcd08aa55c5a3967e842b8f3db20002e9d33edcc63b34a541c746f001b03fe839e5e65b9bd23ccf0cf11535e994fc7477341d4450d280eacad8e13ba45163;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd423c355d8f269c75f147b3bca503778ac37a3167096cac1e67dd759603b04a656c9e08945dbbca679e99c1473bc011cdc2da322d54879e6fffde1dfaba3c870;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h34764e239e585b22796099b701a0987f8a191d01cbf250541d378c0e512fac9ccc5f3ee96a757f5af1f71c18bb14fcdc418a55ea9ce6a0c1a31a9f6c21293a0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5a2c399e032485ead5c49aae812d189c496ebcef223191cfb6691f18c4d6e64a13ac19a32cbd5b913145bcbb8fa17a0c4e7e7e592263bf41d1f9440de6708464;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he575f0a5cb85a8b22c0d0b63cd21d45e98e1c65eaaded080fbcb7a9f34a7282a4dce794b1884e9155fc7640bd49d798b7b3a3991f45dadcd3704f4b7e31ea981;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h41e923129ce908df9d5ef7ee27d61a64bcfb2e31bceab7628d7a2bbd08a2ff23a9f4c1159430a17953e9db0569c18e5ce7c402c22cb47d01ce199765ee0fbadb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8024671ddccf9758d02b085a2d59496e65aa53795edef430daac28e28c3940e9311349d4819e54712397e15e437ea78487059975f276dbd288ae6793a454b40a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha39e047c7e70d997518bf048b39c5e3971bc3c8e1e5ea3f3a7d290feaefb42f800e32024dd05e831de3fb1ba7ce15ae8bde0c929bc175cf76e90a3f53713851d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h18115f4a9bec9874fb062e07d3e11331f9925129d116debc82a96463ff412f5688a5905fcfd33a3e04f819f1fc76b4c7caf9ff475d418ccbf22c77b712f9bb5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdb3c8498d06f13fdb6ec9540b4cc8fe46878d064ffafb1d57e39e9fb2ac7e0d19c88b7092c9311dbaa1a2cd27464d6580406375511e949ec732bca89fb987420;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h568f47e3b3f43fbf3b7aeecc8224365393ea3413065f31ae610138387585ec20da5e78f244f32d9619007438be4f925c334e2e5bd4907a910072c39ce74d6556;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb05c2d100830577504fe582b766c65dc34bd22f1c9272471dbded930330c27898e58e82ad25ffed32a0c7b8e4752ccb411c8bba3e1b2a923998742c1804e86f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8852874d0309d673aacf362dbfbaa167a03b7e6b199ff0f6190313d096abbe758977ac60dcc22275a205a58c1ada742b24a35564684d11414f80cd3943e0bd12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h41aa8681af5e767ccc0fb4282b6fd84dc69669bd95b838e4d7b7af70eedf491d3df08ce81323302c76e67d29a7d2da5399acb794462a98f144a18e24b1b30845;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd22598071b9860dc5e0183acdd31ab6b5e98f44d28080dadaac9c2dd5757ee6ab67164a391da329f503dbd07c49127646f6d69bf3a8fa55859180528c88864cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h21b4e300ddab58b4fdec356a6498b05eeac51186ef30c901e787a25613cfda0fc841a94002c36d0c89a1e73ad9253e98787e7acbafcbeba04c03c16d7bd3a772;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h22b78fd726bdf49fc7664d43376cb141a6e9a7456d6f599372460ad3628c15f8b92a6800bff9c4ff845f4fae39d3607cbdcf396923ce522f4fad16d73de90730;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h361b86893ab01589bf4594828ddf713cb8f5bd0979960e2712e785f8d56f47654f93376fea8704d53e2ce297c4a9005f9b70488c2aa630e1325e7221a6c14a63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf98af5ac94b5aa5457997eaca9ff923712637c6d9abedfe7d9051129387d42856b0d62785a249a531ed4195efd621ab16853354d76e4cbbe2bb0211ecb59ae0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3afbe07b4733bd4f0493379a7854f4500a8c1f55dc9bbb001eea871c892d606c39e990947ce17d3de7b4a050dbe32197c6855b9bd9d7a626037d5b4e74948823;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2fe67a6edbe73e46d6dbae6b43216ae44e377329b40967182359c28ef76527b85a080a6309d2c34cad964c4fafc8756e7db92cc5669dda9c45eeecc49878fc57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hddf84714eead5799909e52e48510d1b140a1300051199faae471e149ceac69e63e791e5aa06ba7bc0b344db94cc9c185f95efba3254345cde3580cc0b5d2324d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb7599306c7c90c7ad0297d7ae3ac44398c6698e5a3b372d0ad73fea1e6974cf68f265ff8487ad2423dc8858d96acd658c63b5a79dcd85705b090a8e10ea0bc47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6abb3804258a15e4ceee2d2e16fc471c86b130a0ba3611f4aeae7ded6a8f8a5f59099f448bfefd3c998c2af5318a5f22778ec22ab59ee82f5df791ab0122d29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb677eed1271fffe165ebe8ccaeba1aa334aa9471deb8eb7e5ee5ff2408bc97ed5a85c7c66a655fe38e002aee007d6c296128fe6076c28658cc261c3bedd93c5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he1fe8d0c1e1439aa2ae2626b449940ac18eee1c237a694f0ce4971c65d6ad98e5b98a1dd86d3a25fc977e0e9aa085d39ded10ae92a48c81b6ac06643e7e76020;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4ad42894cf6e2a39e608b5fed760a34d60142f4ca9430ec8e9c5b078eb53139c9bd69bf7bdc464daa2da56326d8c76265bfda9eefdfe99497dcea9ed06a173d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h903afdac9d3d93119d2e68668585f70f16fa7a59fb2f76c827f6a2c8b95f14c2be637686fa0c0d974454d2d9db483439587f0bb6cb3e22f20a36960fb1529aa4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb9f3ce6676a32f5c1cfccd4b9674318a5b6ae25bdf15d68573763adbc22ba4852cda054ce185b71624121b6baf6ba4ea3452942a8a7eeb8acb772055532da0f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha97557bfec4460b912bc573905177af2573216a132743505f4ecefec84fdcd645b4633d4ad597e1d68d2b8423445500e5481d668e7f331b04e37a93ae3d5aa29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8ea066c92bbb1f7f3a3a409e47007325c02ea0faa6d1b6e8aeb575489f1e92cd13cb8c51f1c10f26f4afe8b6662a51198f8ba34464758d2cad7bc9d478c54ec1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hbd9f83256d3418799a8d9b7c7fb601625dca85f5400a90d08c07a7beeed27c55913f09a835f8d4f9f7dbb7c7fd5a955d181110558761599a563c002b3ee026ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1e54947f37ac937e5a92086efb586ba1526b096b8ba85aafc6dc099687135ffee08f52d13dc6a19867ac4df0ac2802425bbd9abbf5dfc49ee17ab4a0e3bd4cae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h751efdadca7b2dd112dbf2d99ff0b59087ccfc72fb422b2e1e3db210d297c958344e5c3d2fa3c00b53996091e244f4090c70fcacabb494343c0f7beb30382d98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h12b9705eeb20869158212a2a476136df3e0f9a2df9a8dbef400773c1254613a7ae2e911fe2e44b4f988458f68493de40f18c1af2be96f769c1797dc2a53c08cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc1028a6a490ba8684ad5594a31b0f566d8fc433eb2cfcd498c4c21d75644cc8db88b7f3b9ca2bb02f5d5c8057c2d57cdc1494ae4853e1c0f82c0c57b1cbb3840;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h71486f5cc0293cbb82d4693543993b4f523ef0c94da8b5cfeb651c5ea3e27d70b4e3f9d4e1d451281154d8869fe8acf8d410b3d9ee3b30191f2fdc34711213ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8c32c1688e53ece7f700c0a8160e975a37599fc090c01a6a592f00d99cbe602916f4c5a0650a7ac8eb6e504695c0f328cc31e159a73422c6ff2e0b2ead832443;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2b8911a052fa65fa292c6d6f955e95a9e6f79dabecff11528e027db7fd9b93f36470231dd6d20353cddc811e75ef294a62f6cf3f24570543bb2a9eb1c2b179b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd2f4feeb8390320a5198827d8e4e64f27a8f41bb03daf7170dbb9b5d52b356b9c2738c0e62e0a0ddd13b38017fed4a54e3b6f06dad4ac10979d9652d2f86eb8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6d20b212dc2cc88fa54805823f588186503810c0c0b664ed96a0befde4d7fd949fcc4c79c80f99aa688ff8de81dbb45817e9eb990bec94ad534145c5d8061255;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd06979b736d28a2fb60d37b9c86f3ca5c521b05687a99ca026bfdac26d01ac5c88ce440e61a95cd4a1556895b29e4925d2d28338b5dbda5f761b37b8e933a155;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2fe507d17456b7836dc74e598707cf09bee3bc67e80df389363e4c39f2b19301ec031ddc875de481206d212a3d208cbbd5e50761c21abfc45d1e0f404d1cdf8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h976a84a063f0bce6fbc2fe701e729e45f2eda90c3e5958620aeb7bb9671d26b048d657345742730b3e1e5f9d198c6a113224796d5ade1039c7dc07c21498b81a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h664e3e6e2c31ef629ca36ae89cebe832b859081833fec2352acfa12d153817fd413e8636468ba24383f1ae0a0bb8f5c83973285dbf0bd047482e469b5c5d953a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h57e4e1f82822ebaf5b33830133c85d887e1e30d83ef6258e0fbdb66a5725c57c9ba0167a1fb8579390c25f18bcd3e0491eb0df7136c55d6eaca5c07b4febc69c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'heec408ac07535ba2d3e5c27657bae7c5905b445ab54287fdfd7e9f802ae185967cda6c170cbc445e9b677681718c4260b982bef38484b38b936028c1ea4130c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h327f6ac106fa8bea38f90aebed91072b1c197d5f5c45d75a848422e163083b2d955ee44f96c6dc0726be4cd0946cba2e3d72f5161be3483f59d29edc97e64241;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcfef1178425cc214cabcddb5ce342afd3e6776614134db4c6ded7b6c4e0eec385327578d99072da6b1666b42745a30e3a77687f122b43338a2a5854143b0eeba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc063d5b45077c31dc91ce8fb2690b113f0a7909d4be8aed2b5916b8122dfe85a2823b9bcb88392e5ef970a029dce5f6190e2d7be7284a87125456df715bf5998;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h71cbf35c33537066bed8276940fe8ae39b7ed23c54ecab23aeab86c5e534218573e9f2fa2fd54710f2a193a20bdb43dc269789ef6ab592a17fe2eb3c450e9e21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4dbf9e0cd05a3797d360a7cdfb651b4ba4e8453f90d62b3df90bef7db783586755ef431b5da187d7b1967a02e891d8be12367700183d17377069b96fe8b12948;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h17d0002fdc2c39c21ed5c9c5cce77828c606631d9c5605aa3addaa026cf65a48917b88ed6197fb09139f4057e585f2bd3552036e770189c9d972b0537ae14db1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hccfb6497af4a29e78459ba8ba45b3d3732b2892997937f3d100e0a79f836096310f5db5fc92c8d5cbbdcfeb17e7cc34b0c6c1ffe4ad0df2a4382f61d8488b06d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd225fea79a77882ff70ccf9ce45e5505fe183527893bad1b313eba62fc97d5154b098c81c6f6c4d288671f6536943d01fe8431fd59f48a6dfcdd00ec61800a65;
        #1
        $finish();
    end
endmodule
