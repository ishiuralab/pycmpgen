module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [26:0] src28;
    reg [25:0] src29;
    reg [24:0] src30;
    reg [23:0] src31;
    reg [22:0] src32;
    reg [21:0] src33;
    reg [20:0] src34;
    reg [19:0] src35;
    reg [18:0] src36;
    reg [17:0] src37;
    reg [16:0] src38;
    reg [15:0] src39;
    reg [14:0] src40;
    reg [13:0] src41;
    reg [12:0] src42;
    reg [11:0] src43;
    reg [10:0] src44;
    reg [9:0] src45;
    reg [8:0] src46;
    reg [7:0] src47;
    reg [6:0] src48;
    reg [5:0] src49;
    reg [4:0] src50;
    reg [3:0] src51;
    reg [2:0] src52;
    reg [1:0] src53;
    reg [0:0] src54;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [55:0] srcsum;
    wire [55:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3])<<51) + ((src52[0] + src52[1] + src52[2])<<52) + ((src53[0] + src53[1])<<53) + ((src54[0])<<54);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40f952dfce6ef31aa4cd7b82afac84b0b8782e2198b02cdea99b8d1e41b9fdc691fa3da388e1a97c035d69d07357f8634f6678095548cf85c2bc1546f1d2ae92a7f41ea1f6b37c4e3467eb916066ca55157105850cb91204ea77d9eb0add92e33e5c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfadf61f68d7571f275b3529b11cf1931c4b5231ac3faa275a5553a10d29bdff576b19fb5ae146b0e782d5216a74e007144cfe0a9337797fa5a19ae5fdef8d9c9d759a222f74ac70664448c632e8eea0cb6d52f358d3f14b2b87d8d448d6174b2664;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf071250ab56720fb60576849fa4315e4ac4114fbd036f0ba082d8156c6bda088ac1b6c84aac261441e8becbfba280869aa8119a3fc09b27a43a82aba150e9b4dda7e36a0deb3f1fdd90bce7380bffa677d1a9072db74e090682dc61eadbe039638b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c1bf21824077478ffebc2f489603faf59d7c6050c3438d4b772ae6341be616a8a425dd9a4bafe6beef82add2d480c67adfdaac947e5d025b4da2509b5aaad762fc37184e713949e80129a458237ef465aa9f1b6ea2a04e3d5fdb0e2c955898bdbbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f4e5805ad3a2ff4dcf894ca48aa56e7bc43b6736f99931cee02cfb62c127b774c686d82603b11a20ab582f5831af55960e2108ebff127a47ff4ebb8bc2855a7883ec3b4e7e16419f5eb2170403dd68fffe5d59fbfc193970a4dade34848a8ee2c4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48dcb3d01c21b022bbc5d763968f5e14a13f8ce2458c55674c43c7e03f7a2359de81f3fbee0424e67924c51970f08f948c913fa0f5fd72626eb5fb7205ac935e04a344a3c1c41ef8fecc34d0d263e095ae96c426ac2de5d16ab6f869a443bdac9e5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h699f9af3a8192a233c55b231a13faac25147bf994b1e6b089a86c52d992ad2e7089427f261225c92e300fa5544dfc45d4c6af2393c5963b8163db34a104931433b26ea036dfdca3fd5b5683974992067f69c6ea5cd6e4f9372b51c575b098fa6495a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98beb8237fb55f4fdf8b275732a8a55c4972dd87bda9442825afc4d227408ed9d8451d5d2b872675c8c53c9cdcbd97ca2ff31b0975418759b5e63fd8c9b96083ac337975df6f49b6fb372ab84d97cd86fa893f4cf111ab9bdd69635e24f54cdc2bbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a0e4229f5326e55f6f2cddaa2951e1cc89c0e323a46b56260d18b2c3c809f1ad6f8938ee197f93dabdc87f78a6bb27a8bf106a9ca59d3506ba1c9f3a446d200d0ecde40f3b36af23e539c0b7455b3fc3c37a6af466649a3faca7b852c66474c36a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fe1df056723966a720e826e8bdb9a1d2fd2c2c62344819b307058f34940374c0174bfe8b26ed2b8da58a8035806f16d2c28f85b3da3ee6759b452ecaba9fbd2541c382e54ccb6e7623f64b3e7714bf48f4d93a2c859676999da462afbc923b0cc82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6def80bf2a508c845c6d6ca0165020d0f6db469214e5e0f77cb23d9824b144693f1cc6ed9353ce206680ba9b3bfa7f52badfda59cf77b8178d4f0f6cfcf54e92aba4c1f11e81bd58db27da2fb0d3e73195e7e49631a24962c41d50fd92cb696c8a62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98fda15a029c6843f901cef111c7871c5899fe664d7b75e34aaa636b13e4ed084fd840ebd2ae398aa6db337693fef96ab573b8f99d6b3b88ad8e1ca5ce1d6c78d86f654a14ae0b475f1de14b043af956aa7a71015d97c2c03d4df334f8f37efbd3fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63e867efd46a24c2eb86f13cddded7f9fca4458d61d05a0748f792695aee880e1e5ac289b6ce6d2f76c68f6cfc674913bf9f568fd177522be60d748f9b73a5d60f1fbb48e4959e8c619853e95c4441096500ee17efd20da62565cac77385b8758ca9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d8dd43479e2e0f4dd21e9db52a519cca952c09373692b49b1f140ffe5eed075578fe6d89af29aff269cdf6536e31214c722692648a9d2d5181e67e159430b1f1e9799617bf49d9e5e2cc50ce1fc7bd17a923e13de9e1e28c4f96aa28bd288cb6fe4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a6eadfb5504351513efdcdffcd556beace50bc0a9b028d609cb6d8f56bf5185d91bcc31f964de04fe0f0a076a349f5965d5aab587d6b35640f4ad7e9b2f7aa5e7ff5c1d2d6499f9e09a6b8603f47756fcd5a8ad0afc9796ffc71fb64e06fb2fa5f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b8f0254d1703c6254c36361d2f1525bb1bedcde949efae92b17e8283ffc647377b1870aa600907cd5258a8f82b5d8e57cc32a7e9f873c7faa6b827ac904782a6c151eb573a338fe155a1f131bdaa8ac3dd2caffbb5ddffcf7bf88ccb27d1edc985;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96a13351ff4a0336ba9e49ec8930948192b2a66ce14f6ee5210ebb42b9054a70c03199f0eb513b2e4cb7dd219e51bd0f05b2335402cbdcbe8e8a9d6a5438b78fcaec05ac4ea109930bd5ca3c0b119f7d9e5588dd00cf144286727a3930f941b9a62a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70c3e4a7b16931c76724c937ef3f8b9fab769ed11dc9c63593a6d31170096c5e29b7b859701f1edb3c011b603b9715ad6e9e175fc47cf62e8e2db39360f4e41a40a05755eec246d29cc3d61b28318b691935b1bcc51cdea1fc5d68294d573f45e90e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf032d88ce3027fa76caa775fd31631712b325390c453d4d5db6d55fd2bfe4ef1b870889c3b7dae252387d933f57184e6993ad924c960a1495bd980bd38a156309cb40d2e8ca73eecb2d6f24890c22432357a3f322805a85e78e32e952f3d8b4a3a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77172b082853958dbdc14a67c1eb49919eb883666fcf37e3698f13954d716f6468e220c9191608691bdf35e80747cc3d5eefe24445636ef46cc9da52ab4708f54e8f9390bdc5a6cf73f9576182ff1929eae6000710ffd3d2ac2473bcd52f82018e1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h516b018d848a32832b81a33f34e7ab120db0ec4bf81d20d16ee5ba0fd9ca72aa829b3a0c0cf293f9064e492e23bc853fb40a06572ea9be348e1b349adbcda1aa033c72ba1fe2fa71c4919cb4d4044214579c7f708d1a5f4d142f255331a87f8d4d17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26c91dccb47a8793d810a17df7bce0246a0e89b25316b3f9070c0f08a8af26ee211e1d13f978e397f2296350ae5eb1b7fe2e7506895546f29813f2a93ebcafcdb5d5469e5ef70d43133f16e5959af31b0257f4e6f0f1b20cd6a82ad8dabb842917b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e0a29dca52c8ace606791be6af156931d7be3e51a699a8707507d6ab2aab0e12e3c755f0281aa3e7010dfe86fb2c1c629408fb8b36439a7288d5247801f4fde4392e6a6b9b8d87276ed8ebb6303d28a1b73bcb678460d72aeb6f61ac7500bb4567c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0c5802ef152c25f51058ceed4d2f825e1917754dbb42f5f1e5b518fa2ee527c7b9424dc9668f542c633452a85cc7efc024fac9a695b8ea45d5e49a62ff81e24dce6bfac8edb8b5d473260d882f64952ccfcd2072a6dbfe37fb155b37681c9701b18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19c43610edf690f2a99aed78d4b98e5cda8416e5e28ef0741eeeba9c829c50f75effa6a7688fc2795b2abe7c2e0bfd8a0305fc67d7d8fbe3e2845ca98ebda4180ec8ea36193b23db6447391624d6fe6350d0c4d07386877a4921c8b160296b5832b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11f920f9c86f49898307a1630866321ff978b1aa325db384f057fef8ff3eaf5b814563295d43ba2f30c09df12df43ce638a142bf76dc6f879d81c303b54d0acc1a29ff6d63b74fb7c384d259544c967fb3b95543313d1fdd21b5b8ccdb568fd7b51a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78e5dfb8468788a617970a2049007e4a12a36dbb1f5d1d2e298e2c45d79b21ca5da4c33de1ae9512ff4dac86d40f744a582854c0fe0f105b3958ec6e092ab628d04be7788c499444e46d0448c1a2dbbf596aa4df9150aaefb9a0b6dd86699d21378a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2434c03e289fc1c21f2376494535fa4b7925e80fafcf38e4749445424b68d64680830b735a0fd66260bf67f8aa3146962a4554a5a84f35bf8bf92d38fa039c942f31e14d3f77091bae92a8c9379bc807947e609bf0f3167f71a7d7666e72d2b59f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb25a3d5570684ba112da8e38fe2f55aa1d4bb296a5f80142eea49833f9fbba81d69ab90f1900f4f90b4bee8fab07f44458b23c0c355a75b32c9073724f40f3c00d2cb6c4372b581cffa073ddbf7ffac42f0ec49f3afd721c552c8cbe0e29510b29bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h170ee4543a44be326e54f1c6bd5c517792791558e09e40cbcb5a859d3b1196a8034a00888b84aeed5dfe0d0dbbb473ee3f586164e0848232f128d28a1ecef1c4b799f737ec1161304bff90ead6a01d8f70fb67468acda3389996d25742e8fc623cc9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77f46d98118761920caec70348b4dc490246efcaf6dc3fdd44e476c0e66e0921257c65add071a2a08234749debcce29875758219176deee3dbd5c2e01ca268c8783f3cf9e0d9df749291b1a11d8fa006317dac92a066d0398527c8586aaa2e4d7ed6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had5573064a0e8f1cb67cc47dc630aee60dbbb7ad4e5a5a90f7b1eb2f9aff739c8279a62c155b3bf083c4226b90e757c9846cb4682c267d5a0a84cee7c2adffbd98526712cca954da4e29e87d6b8c4482781b3726030ff8eced23a3661952572b124b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95a352545d30c3025639320877faf519765c1d874376587436df1709c0c7fb64c5f671c7d606773c94f72c2339563ce9ef7858073f5ad2a64f1620db290fc9909e0e6fec851061da3030296c1f8c8c8a560c92d80ffc332b4da5e7f0a0642e73493c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e8eaeb49e2bb8cb7e9629dd0f2d9ddd1c1188bf99d5aa142a9220d5ac6382efd62e4c3f5f0789d5561f7271adaef2d9d1e3ad12a35be05ef8256298d06dee1d1fe17488aad3c2510a42198df3064ae66f9052a8a926faf6ea48264cca2bd8219baa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he745df8f44ea1acf8ff9f438e67bcdec3a4bcfe7d52c8ab7240e3fec017a866e5db2e85806de6cabc0cab11bc61a028ad68b9a59e412f1d3f27c96ae6be913bfa5bef196ea32f1dfe8992e3819b5775df8ff55ed34e3dde1a1e9f10c539970042976;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23906597876b8a7d6d44dcf8c7fe5c5f28ae71cd6675a877ff9327e4e054b5d9d4c862e86187ea104c7a7996f2632b2d06cda4f6fe4677f858e60ae444550fc0e3b0500dfcb0370c25cbcbbc8523f98d329e499ec649fcfde3b8b94c1e6da3bdfaf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h407ccff9d6613018e837793d876e6f5944a48053dcc268e07a85235067faebe4ee9da3bd7f0144228feed655b775b3d26354beb69807e4eaf49f94e3a06ae664e1aabf606668036e5eabf8bdd1c4a35e01e3d0188b39fc85a0880a1b677d2c0bfd1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bfa110164d97f29a233a342674c0eaf5c614c6a43a2d6c782019052361119b6852e0fbc923505f5c358ca291e03c50d74d2027601adb6b8d664266d9352e0f2be4ffa473ffae004e788b41ea800af2a0e0f893cb87f12baf10975e1b2db2b74e0ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d5f05db63825f8d91146429990595a2f9a93873169167e4c36230dfec484525276f31cf775e723ffd08685b5ff137137a96a3172bdf05d4fc983b7869a8ca2cce4d407714db245f4086664d248ad7d430b4dffffeee1a14a3ec40a20945b189a56c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88026d33301ea12a1f47fa69bca44a5a937b8a3131eb9f2b0cd5fb3216f9cdc87b2855c688b5290dfa0487bb8ea6181612511c60b41693b10c22cba6ca1247eb263b249478cb8f6b986037e61694e58e5c61b84e0d7ac09dd3c401615937506f5216;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93dce65f5032d60938cb7fe7e720eba3ac19471de858405731855ce6b8041b1b3659b2fb5f979866c4a9cec834f1fa48cc47a9ac4f70dd74b20efdfbc07755269783f6e93b009bb1e3a5612c58896255b17dbc45aa46a04c109f26986be4edd2c83f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c2ba8fde7dcbcb1b9571e1afdbb0b42deaa99c35376cc56943566237d5d906ab79c9d80476d3c6bafb73782483522c81ab423fe8e9e21f7f76e35a19524cbeccd529563258cbfc2a75f964f6efb6f5cfc13ea597be2d014b41accd8997455ea6dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16afcc80adffb849d7504b2f82a43dd595d264bf5832f833276841aad9dfc3eb76ec8465d924b9d4217d5a344834446ed12daae8ca221b72f91c11c9a9e27420b0469f31946578b48037e2612eb572d6390476e1bc83f3a02d53fd1f52639a3d3777;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d6cbac2de7a017753d6e21de8dd2fe211975604a992f923736852acb002356199bb1de1b722f0d113926574d1c2e93bd2a374a7445079c3cc0c6d7fdc858e206965fb5a7b22bb3d4c0ea526ae64a3a0fde61c1fb8b9287ed1c7d17a8b8c50cc591;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h130c46d487cc79501460b1e28c71fb5a233e36a814d9501c9b95562f98416412add65d86d5dea530dabf7e701449c3a1952cc27d143ebb7d0c462da2888c945ab6f3908389b31802a5418b899d4a775d7a98aaba0bae49175cf1adf8e3d615cf3dc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c9562cfc3a0eefc5be4ffea465c4775a8b71cc4a76751c11c73af033cc9feb3097a848889767857d3e2c0576e20ed22a5eab1db535f6aa23d25e06fa8c9843c01ce8ccc6ad53a9c99fa5e6999f1049cc7a868f2be5eeabc7e903990cfec9b8b011c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf11c8cfd413944d8cd4b9264157fd1f1fa40366f9655bdad0517e5e565479d51d1e43b70d4b992d508fa5093047bd233c19145e50dc5f38b19488485e4ae2f6107e75e1a45c999309fe297620ebcc540df338e2980fb6cc16c8ca851bca6f9bd9903;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h141fecdc4b14759ecd24a2f790f1f00a0edb31bb3f5deabb9cfb9ba4d423c0395e31ed5a940ef81248ae4a53e5067ea27f52d742e035d40aaceea70430e4ece2b387af014b374d2eb4798abab1163d457f083f3bc461e4d12fb63076723fe8e66f41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1d031bfd20d0344ac1bd9ba948518abc5066a40a0db817cecf7b7a1ee6a3b3db9d5631f7d41abf273b576467ff22e6042eb5f74aa482577112950dd3c1ea4fa9aec8b8238367bac87cce8a6e773bb56e95c3755bb5791024c52170127521e520f8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3fe8be155cf39a3e0c727f4b0366556a4d5d31fdde9dffbe283405f866fc7c5db89dfcf61988ee6be74f85834cc79b954b5bf14a2e87a3e58824bcbc36262ff7f43ebd3cb6af87da8fceb81dea3484fa60cb86fcf5df3624b97097739966c9932fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20c47b9e6226051c4e815593dc2886a3040f3a6533a17e2bef06ee9737cb2ad7bc453ecbcada66e9df874508d9591768552e954d35da833dfd0bc3b043cc95f5965594610eb2b80345e13fa810d90e269bab3dd8e6ce89f61cd3aacfdac25233f9fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0f908146572093695b27926b3fccb2f425e38de94b29dd88559b25d8924a61c9ffb7c255786a68eac7df12c552ae77d2b0ee16e881a28403a5c84e4e83b026562172c9e8902d541a58ff2479f4f8792c3109ad19094a05493a14906e17589fe4d6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64340e791f058c47a74b3e87efa9094de0f029b43ac068022e0f85853a13f2c7d7cf9121df046a1727098cf5460845edd8fb3b2a7c482669f0f1e0fd9085d53399c206289f4c643851ae09daeefd06a7b868ddeb3757df072035dd027b73cc88705e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0df6bc337143eff8631594b657bd1a9356e9149590a8d95ebdf2fb7e6921f043a8ab809b2efe1ac1e2bf30c5f6e957ff293fd88dc5ab5c2860579a96ca0f2452b96ea8728e22c040df37f2128fe5ca96bfd92c04c6078839b2cbddad266dc2917c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a8c5429d7db069bb0d68a483b39e8c81b5fcec5c96299db009e4c40f01daeb0c15228c919d4ee250c997a5164b2c0716ecbeeb0e52ae206ad7c1aee5b9ed73c71e0d44794f6d3dc49deed055ce139c082984898088ba8a675b5c122da686199d6f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94a57c70d96480c5abf32bdac4be7cd63a8beebb2bceb7b127643004ab779c90efd7c41fdd5d4a90f7f01da8ec8a928571fef031da8620be8438ddf96df0208f3f90a87353a5dee90027261e25abaf07182513a045746330ed95a87ee72d5c07af9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c76627872203a56685dc4a25d85db38062cfb0ca5ab601f774cf6b15602a93a664ac6736a24d0d6861702dee656a6956bf5fccec09ab278e7c1ced8afed28c01016b2393cec1399bd079979ae4996ebd9e950d372bb889f03dc62d7dcf568a9a7e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae1db5ec3dbcadc3e5889eacedb47c0dedbf9ab8050a4937b387e3fbe01edd5c9444ca957b007dfb0d5a91d4277dcdfa4367cc99d8ace50f22b4f1f2234f5c62706b15e1b90c98baf775d177cb7ef74b30d537e7de9a769f0d136da5511f0734cb88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h117210ba6203b233e2b83277d4b663bc8dabf55597ed935c66bf750cb609850e8d4e3b5e20f9b38bed380e49db1e27e215a826055d5593ddede853f2ae91dbe8dae926e60704c96193d9d0a6166fb303560f321009c0763d25d2e5780c5687bf0319;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc9d9ea633e639c09c989c7ce32939de4b856ee65430866e925e51d61ca047bcd63b164254a08e0c470e81917faf1446b61851fd028cd23212abb2dbb9522616853f4e33550dec5fe768e79056eda12be282eee494f3815468af28fa98b2d9b3c8c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1914134ae934b38d5f8f231b8c10b98d04d58066c3a693cce6ebaa35c987debdca81bfb7eef82c0f4345b0da8cfd482e0492ca81260b3bd5853af779755971b26ee30e8fd6ef8d72ed1b97ebec72e3c59a64f8f57fd2f1c83700297cf7f0f1c7ad69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24ed6764f2d9d33cf0493c2000ab5add6d284b0515eadb1a1b9c3ddd5672fbbbaee925a9702050700c5d27698f62aa78a19b280c0607148449daeac6e296adee8b5fb5ae0ef1762a57956b60c650e697d82d48977e3c0312233444f6274de4300bf0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8ab2c80f9b385ed3c6ed4ac958eb399b3d38648549ce7c053974c3d7d4efea7fcf9b06fcb8b55768ac39c4d726f67c45c85d3796dba66071efc843bb16b76a30983f85d6eaea46aede22397742302404818518b4988bfe2d44696ccba0f272d8c78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf386b0a1d60bd5445f1a9479537ce7f9f007545bf79324c9d2bfffe0c97f54872383a773644b97379a97c18c9a09a4b3edca8efa84221c12f6cffc2c632e4881cf64623ea9794fbaf2484c7d4c1a1273bc8c9fdc1c24f7c74df2478749061a45de1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec50fe36bfbdf03a715f6bbcdfeb2036b82c5225ec58e4ddd23b9eb1678acf43b9d3578a4e5988da390015c16a6cdc82eec1dda47d57cc7dee2ce5d9b37fe39eb5a4222f4a16576128d774a3cc81b66a693036cde9ba12f5a3ff8d2be4ddd9f440df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11027aaf1146bcfccd1e624fc9c3112ac357cb9bc4f531017e2f47a5071f5b84316befc5fad85d6684631687ed24a9fc12cbca08d6d153330cb487179950612e0fde5d8fd67d1b43d0fd4c2dfa3f507cd7d333c4576e65a18ed6aef9dee1e4f3f012;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb481c0ec208aaa2f26a45b88969e876cc76bd2a16a26b3a628a124e117f716af03b670787b7a8aacebfc2a36feaf6908a593137145a42a8591f97f4ee73d658aeff0e6c6d2b67b828f26a94294fa443011edc4c816b8c9a6dccc39b2043f248ad295;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a4b898723729911dfba0227db5aceb5102ead4fb3fe709f23d95afad1b2112513d844d3b485243a9ba6cd1096f5425f71c42706885494b9a9c1ecc9dcdb4768ce4155dd1f4e2d00895e93dc585090413afb873ca7fc96362a49cc61876806ae5807;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3abb38e12157addd52e5f51028bf33a7f315736fad9650062991ccd52c3c1a5c76920e0ec27d46e3b1ec623cc3fa758a70a16b642348e209ad092a7e2ab5088b884a4d96f3f7c7d4475f0c7916a5fa8cca8a24cc348198929789e9a9a6dd4a8a3324;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa6d75f32e2acb0ffa1ae69b035fc5f14d261994505c1718235b603774bf73bafaf8c267d925fe2e327637e6d17185d86c55016a2c028c5f28ce1581513babb4f9b2bd9570411e898b176a138221688744bb543fa248561aeea24433893dea53cab7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd527e2b72273bb43fcb389e7eaf55b4d11f6c99ee29cf9d1d965ceff9f0ed65c325464c37018e8a4c804ee14ca7e8b0b31bf611ca5d23257ba8e8f899704bbddb7591be8b18e5b1c40712f4d8ea23282682ddff10b1e9bfddc39b75a1e253c6e12a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf31e4e1ee082109fb6f7cbcf8f3dd645d9cc670f1e2aad29137d0ad583e52af8e64f97d266b137b9e4e0a6e61c95a7a5a6f6263f29f95b28b15895f5155604a0355a163be0baa041751b769a3c4bc3f66b23adbcdec436b695ff4de8a8af7fe2f63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h456baaaace6691db15fff19657123bd1d3d23f12326fdcedffe5887f0ab771a60c78cf5e59a71b380953398d67715442e0714f4ca6153e388aea3db66d6ab37dce5264b6a9158da4efc71b3a80daed5709522a41c7aa8ef203799b114ae8600ecf95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5426dc205f8f9e5ac85a768d952541eb0088afb89c3715965fc312a68c7544b6a7b5baf5f6c2ac57178a97aa45fb12d688d270549dac2bdd699ed7116f0144b0c7f0a0cfd05f233e511b4b724447e40e80d3c8553ac9785b3ac08f5d465c2d2f32dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ef6b6a62f7f53458d01041506b53fe5e053d05590bd49cca604e11cbb160337aad2ab268ddd6793e9e9a6a93feb5d20664c27cb0a2cdcf74db05fbc71306b499849d9bec92511025c730bee5182f85d6b512819a42a1b3dfec4f7215a100e00f6ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h776056d768567a8d0e7a800fe07e79c1acf554e9a09cc1e82cb9e0497e9e85e12a906318efad02cb1da06bfdf520c41e894c7b5b0fe0ba7182b4d29bf92ffafed232b3ab67425cc04eea7ba744587e509b6302f7f7c7f20e0064819c486aa21b7b0e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb397883968c40d6a95dc81711608cfbba2602c7b4a577209df14cae052482866503a3bbd044ffb676db4de8e0ab118f8530e40f95272952b23d4ef49184a542c9cd03aa184ff6e656714307b642bc2fad22dbdaf2f94b639eafe2b05c61c1bfba2d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fef2c3d67bd5ff1d1c6a0edcd7f5f8eb5eace5fe8bfa8cec99225c4d2b3ad9a7a774979d7db5cde945494e71dc8b15f93fe89646ccdb004af70e475aa78bbeea5f4db57e37addb77f5f31d58c806623762db4c8bf2cd12ef4ea9df03019f67f654f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11d6e27428ccd68800d80b1b8fcbb475825572c349ea2241b6f3f9f8213c69c031f2ae481207469830a65d0694b3478242a6ee55cbba3af40f841dc9a7c969d775ebe3f724e4b0c0e49c27d371c712a54cc1706bb19af34a9f327437c3b8e22249d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e39fe3df939701470bb8e4be6964eff92f8c304974f97d56f7e36d239365416342043d67e1816514c10baf2d732b57a0715dd17442f9033780873858e4d7685246a6befb2a34c20dc20dd0924f569f86a892d6f26006c26c479c68db02666f94fb9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2484c50e6df4a139d9b4a321f66c4f7911d11947c8671f3745efdcac41df674bc3ff3de718405b7522563e29a763b3792b3546c688e82b0994374efc2b94782f906b351030d45f6b90052d0f022ca58bbd77c83d7ec95f251844e12ace8dca753b7f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb40f0ca85a4aa5834ed3268754af02a06ff70dade75475c8d0e1d3373f8fe4add88ec40bf6079395c59ddaaea51fd6341f530772bee1521ad2dbe3d9db476b1bd3ca24b30dee8a09cf48be002c2b92870de87be28facf26f77d58dd23e6798267db2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8d33309e588f9334149f54a44a99c520a1c2d268452b3f56c35cac467c6adc0814cb93b361e3e313b5b1ca298e7165fd4dbc2989e687f517d85e6a25331683d96562de22e055f7fb5f840aaf7b812e170d9cd7568d004a2736d9ae0543eb13cd640;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b8f977d88a23ec9e5d29ca3358a0638531f726af0df1f738956d3b8962bec7b80e37bbb62b6bcdf12db2e102aaa32c92c495dca935e17de636ed12e02adbdba4a4995b98eeb894860450a5220dc5eeea5c406cc413fb2371e4614b03f0fcdc64566;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb43b2581ae4d0d00774da803742b63e8885ec2f01030c3aac1fafde3694ffd48376db6e7415835612413672341981ed1a231644320eac29773226e361849511330a63d315dc7a1b2635b5332874be1bc2b9edfbc41d9e75cb4532d796aa280455a07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce97b071347321977bb0dd4bd09b71d9df66381f447a64ec0839a23410e1d05a19d369e0cf1d95594597fdc438819378509183a2ca237ebb3cd2f762dc20f6042fadf8ccfe5864cad76e120816f4f836f11ea523bcae8a65295cf3bc30ad3f9db62c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75b31608e88a868bf9f2b31629a6904f698491da541ca06f68ec5a82edda2deb02f23a24696a4d45f2599b3011106f004edf3f86b6da86ee5b1bd565584cea12fc561de0c1a08b7faee3cd2ea734b721e53ec14dc9e0b8bc71a53249c060af4d8154;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e36a88e18a4e486d403be2073a1a1e2b73a04c15add99b8c53d0d8d73c81c6c8320b5bb91b9d0a5a72fa088d849daf827f159bbc4d82752c122d8565dffde8c3c933fc78256cca1c754037af812e9ff048466a82b7e1643170c2cd7cb79795d932d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bde783104404a2febbe7adb4f5955811fbd7d3f51e808dc9e910eac31c00bc9c7b6685d2726687dc2cbb5f2e981be2f1c7caa4f0365c4fcd3bf269728fb41d7a462c54416388e89f5dd817a7594a4d0d82c2d55c30c2583405924519f0ac3c4aa23;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had4837ee681c399763ead099db0f0c48fb4c243dcfbab0d517e32e3e57544227447a032b9e6f4a6fb86eb2c705261244f9f356f2fd13cd82a853e1bb574cd4d73a6694f4ede03e678e701f0cbbd97fa38e99c571c184e94616203108f06bed2a0139;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h539a836060ca265aa3c1dfe9610f921d28b280bdbd292d232c563a5597042720a47bf2c0bf0d522dfbbe1ef6f1223a778bac223bc46802061257a1ddae51a2115d51c29d676e2e28c8c485c0955108801418ddf37258452062bda2dee23368e48476;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd49e8fabfe04b18688b35fe59479143def7f30c379757dfd4c22aefb554c15a015f80062d5e9ed1ca8146db5b817150348d01af70d527bccfe5f62ce4335ec1d391f08b258258476a7d6299ef6624a2b83dd2ab56e2e8de54c54bf07940efc703869;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0bd0afc11ff40e6cb7a1203d5139e52987ac08df117dafc7d58dc085a7786f7e2bc64fe2e8bf04fd09e51b5fadd7f10c9d8f738a148d67fd3a29a7907d141481f49fc49c3bc8e889b9b75738347dff2ee13de21b26f87946f86c4f77c7fe7645244;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9ebbeef46e10b630f3c4e99f5b71908325d5c172752066698c3a8ce4830123c164614fa92416c618281b6eefec81d4670d2f7de37b24f589e4c392222bea2bcc5497a08a8a6a6cf8175739c59dce49ba0d802df18e9c06eebd0ebfefc5915e394e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ebcf20ee94bbf6fcf628303894f82ffb3772941b53210e740859c24558d28f63d37e8198be88be132a66d0ade632da615abd556363f166ef020affcb71a4afa0a065671ad051de3635b4cd760ea5341132f967370a587c534ea6f345dd612a8bd81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f6700951440a70b82827bca064fda61799bdc77c843874c8f8401af606463d8d2ae284f0342c67d2fb9fb1f5a262a38bf34d3efad71acd632717e894b5bcbd0a5a4f22c0264152294ec85b1b4b9f2697711d69f99c128370963af5b85462031ada3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0c4ef4742977d64dbe8100acbd0bcf139fdfd16a8ec8f194fb3e434510ca9e4435d069124a4364f2190734fa604eeb00c9c6eb29471aac9b4c16e8bf10b6d8a063b89cc3c04c6863030e16bd0a9f448330d5090e3d12383d3037f00611e8050745f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b6aa4519a67473a2f7943e3be5339e28b909ccbcd92b1128e1708b704dfef2eebceed895309697430d73ef93d08060ad6930ae14e9658be5fff9209ed180e325bb6454e2ae31f14a192c3c91c90a6822f981ba743a8ee9605804d0b8b96963ce043;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8c86c0647dd3ff4528f8c2457822d7280f2c52a066a0b639d1a21bf65497b5d8e0c15b254ba3a023e591a7cf76245d23c7dc457252be77a2ae592c45ce5271957ec97f1a4458f26d5b355533ea5a5781cc6ad1be484c1418d8f0595c68b08a69b04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8802cebfc6c6989ee24ba309c7f4ab182e888211f75744c795463f48d01555f70981e353c1bedef1e17a922a00dd13ba98dc405c6a5a7791d57ac67182d69bde83b3189858300d00c7d764deea967d0e2564eba03130894b24e95f56afd180943141;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbffd222fc4b5d2fb712d14e9d9394d96111c04ed447da569e3ce5425b6e70c7aece1497fda82e8a295b662798484a1aa11f3564140f1b2eb6f46ac7a5dd6dee0796132c302e3283aa1b8960431aa6b2dea7f396bd346f21a122b9f43c89638055401;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2468a0128f13932a01dfc51f9f4372627a96ce9156ff4440690cb18395a875ec701a75050a1d59bd73f66a5d440704395f17ffdcc6d8b9ed2158b2f7c81a9473589ae4b1fb9144ddf21e06d0c7ded24b6b1df45826fcbe2acc9d150724713a3e498;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbd45fbdb71edb063c0aab076a65f14f0b84f5a2436fb3480c5f1db335e40a0a08aaea26486eb7c948c1c06ea9a7d4fc1581d4c70b46f6f15a30fa00bca168e787f85bcd7c580f0cbce8397308c03d278f1e9332c38af1e3453e7046ba43ff60689b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40ffd69647812ea9bd02a157bcd1e89ae48846298033fbb4ed6abbd091b4eeb42c147c6817d7b91e83105c85ee2322c607b7fdf3ece56fbaf0e9ebde6eff15ca26710a9df4c146bd291af8e9e4f132410daa8b9b7de32e8365b7ceaf0c687fa7cc26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec5ac9cc9cf285693d214c2d998c09f17b8cf8fa6199f204f8cba6ac5663ba79fae530a9b3ca2b4998178cdebe510b48d35491cfcdf49eb4bf59670a829142b23c3fdda11c0384936a584312457d56418afc1818d5d0d7e649a23d56589025c01d99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49d2606f425ad7eaff256faa0ec10c8a56e0eed04f818c938f67a4493e8ba46aa7cca56a9e0c0458cf67705f5746407563748997afda0d83c72b81910a05b6b2e2aa6f90ba87dfe6872ddd04e9495b4a5c5551c2a9cfdbc5d6455b33deef9e87938e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2eea6dcdb4221f84f2759336dcc6ec283527de0e38ea5d0efa700afbd7dc284235ff92014d768ed500aa581beadb0bec8bb3b350a8e16ce04a63d0350c8ed3130dc445724c44d132a72de9069e5d3163341ca45a13cc013442bb06576bd1c17c0e83;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8706c371e50d3ad177707fed5943c1c1c3f70f347b82b292208a835ae49574270b21c1eae0188d6b4417d61fbd62e0f1652ad1d521c5e8509707e198510933f767c0517ad707a884e223e9d68652e1413d16fa159e22e86ccc460f6aad5e892307e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ed5893a73dff9bdc0ea9344ad8c6dc81ce902725b56608f62e0b55583fcdf897184c8b999fb5538efa7e51d1ae8f5108932b12e5ae063c87de903cc0de15ee51d7c5814277db48c5334e6d8dc5394859222257b1e4e04daa3e838530aea9d71fc80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c42c7853a9d69730b5ca2d06df12a5c337191dce95e81587cb1194ab68b4bdc0e10f0788ccca096edc0e3006d8b516e3c67fab98406c491147d53d65e5e8afa1cccc325e287e33460a93a59bf0b72f10e5aa5621b7a453f9cf0bdb3634bf6f96ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h738e3c2ffd9b19ef09b940603866f0e65228ceefe1fa0c76dd975f2a95eaa5f01887f508d18204a23b14bcadca309c393600d3edd2c1353351c11b36c10b16e5c96dd3aaab8b81e61d739db782be5f5129c7915b87b529e1f54fda1d640d88e854e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacbec0fbce2f8d8c942d3b416845588d1238516a1e0797b00dba39aab5e9df91115e5154ab78c8bd74b9643085bf9e752de8a95df7e27a037584cdcb924ba5ae95422938628da7109279cd4203bf49c6af558ab99ba1f933f66953d4227374878c20;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha22b8e8dd976089eae8970f958affb992cbc544da335aef0bf4d032406f2324b8a941896e7be4dedf2d72c585d4f85084d374142c112a831f09d2c32425040527fecbf23c128fca812ed8b3b98c15a1400d5064edb60aa082a3ccc34020fef7268e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71b051af65f75b072a232af9e49ae2a1dde83797d159a08c332de19d198ee5a7f36b3b97ba9ac35911dbab702772c7c58314fbda09c0af2762796bf2ac3b5284923151635235c52f632552f8dee10ec76a523f1dd8a045f303388c928c2b7a56da63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c9ffc1fa4fc3edf048d92b78ccde5fe011bbd0dbd6ad11076b1eb3fa2fc8713d83795018ead9d64642d9e8519676cb1a1436adda5790fc08d622d52518d78c2348d6e077a655e28a49f7562454c61f7396ba0671923514a3892ff31becc9bd390a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h195d7e07f8283a3a5c3877e8e5f71bf57d57b644e22e210f5f3a63e4005af11c3d1c53d7a8dbb12fb2094a222d69ba1ce165e3c9a13bade9f1b8a3fc98899f004345814c283b97ed40be33e0212b851cf9d962c55f8b015651899b2ba142db30dd05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc52db3205b3e929bc2d2dbca8c6909762ff6033902c46910abca338654190db389a64e535f49771d0127e23c1a688d739a7774015f6b76e7709cece43c932bc224ff963d227af81b58c788787d9698eeb02f7dcc8545660d05f229a7f2525af2d63f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h782e9d0465110a5056914a3470a6e8c4b2e87cead36bd4d2fc37a159215311913dfcaf268db61beb946a0bde3094ad544da908d1f0f614ba601e4a8dc37f838140a9dfa138fe562e3a276105bcefe82e7d3066dcf487947193118e358e3bae45251c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd386de3634e7a1c2a485750ff367a9c0bb81c5ffa6f6e0946a7853177802b67e1cba2bd303d38309684745f92c71ec2d8f2f0ae9e5667bcec8bef1d64a01c64931f4e189402d711f85a345d0fc95d9a4aaf6bfcf13b711fbede95da6e5a889759042;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda33a7aabec0c75a5de8466f2d14c0a7521a94b8697652d84b662904dee9bccba5dc755f52a2a33e5e288aa475fbb4f3d4ea7413d390f681215ef0b58de44cfe1a336b679a15da21ea96b42d65177a6ef367c768aed9265404e5e230ca4d8891f8dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c51c050a3f3e93fff1da2ead9e638b2d0eab299e4b67951326251813bb3a2e620f2debbf390a7f342c35368efe751d114017a4ffdfc27adf12d77b34745a630ae18cac94a0dff6c9e7106843351f7e073aca22d6ae3dc2a49943ec1d052d6a2e45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he956adcf8887414d8db02015d3f019d0a0ae61a9b7ee62bed97c18dea822b3779cf79465a63f5aee6c05298a15a3883dd4ed64537d1ef094c18ca3460e682893ec13cc3392b4f28fc20d754b3e99e6a1fe4a94936112bdf97f3e1ea73503bd979eb5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96eef0a4fba9cdaa7f402f767ae68f4403d63bd3a91d0e4b14d1be87678e40dde5a171f5b1bb45a8ff769284de386c7e9e372d9da5c25d7d15295ba97b4e75b0fd336634f576d47646541b7b56add5fcaa656b5e14d1a897eff4a000ae24bf101ac5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff3dd46fd96e214ac0291ad511f02d1f7aaf708cfe6b550aac9836a0915746ced2d72ace1c3214d01f1af486ae00ac0949bb97721b2cbaae8f584d2539ea9e1badebce7dfbaca93a45dd07b7c108c62bcf0c251952740a3413615892fc0a9ee267ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h856fb4fa0104eb8b4e33a28d4aa8ab7c4c0383c667cc9df16e97dd62ebae81d8ea03b973d30fa7e73aef1316d1e2d43730ecdcc70517317dfcf30e759abd77181a93ea2917abbbb1c00246eb057d76ba938418fa32ef7c6a45d03521ac1dded6890f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bf13002fd81ef6dfc618ffedcf4a171a4badb09c00970390d83244bbaafe53791058e3e92056f5962f62472564ada47f333a7786c79ab0246ce299e2304ca65b07bb543432966ffa67bea67724024fb950218913c24c3ea29ddded7a3b253c58bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b7bced3b7cab257583eb3d2cfc34d0d42c1a358d3fd019685016582380b4936084c733c35908de66648454b33d0816b940b9b9b3432f8eec14e3a3c5bb04741444e5426df3ba5f7da363c9c676ffbf76d46b4054437bdc5a8e49b0257bbd5c1cb6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26e6c8303750b8f99890ecb469ee1d62f3603eb6e22b4b4823993ff9fb5d6df9ff4c99d0aedec166b66f5f9b0cfcbb6670d02557a6791d56593968da65a0c14cceeb0056100cdc8750e38ff02d6f44f2056cbd690d625b58bf9d26d576cdd7b38dfe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d360a80c64a8db64f7e9e0f5a3599c2b00a8f2f19679efbfdfff8bba25cdf8dcded35a2c937625a3a406f46bb6881372cd797ad01413010f9d01d2da91fd90aa2bd0383cb4b4963cd962936359cdc220129fe03b252e6661c2ce0524804e324e3a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65cfbd7fd862d5d56c3df919ef10304ecfe4289dabf551d2ce6c86454f627b59fd44dca6bcb422fd1f34d19534c0ce63c26e47607ff83650dd9811bfa2d47a673a639f8b5f5cf079e72a4769021137b79336cd832094c93723aeddb14a25ec5bc370;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac6bdf405e410c2d5359f778317073920af926d33a523a28c583db68005fa4a5763421e6cc54cadd13af08cf86436c316b5b9fd4244a1054b847ea6b4ff4af22ca9f5c75acff51024bb52a91450ab81511b4a17bec70d3c95a6c562733c5e5ad04ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e267afa5f4f6eb5538efe67c69bf6732d319ceae5e84c7b1be30d990095544090ce10439d2ff1fae9ebbb19e633d5c7bf9c1b1ae501b00390d565f2bd59b41ccb98c4890f067c4a60c454374a2e759ac5c060f61da8980aefcf997fcdf2630f2e0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9da5f09d038d6922c057a68b8bbcd8f8e86079211478c94de9a38fd45467df36bbdb96a475c121c5cdf287360b0300c68f0fde0c48b27e7e9913a45765c9d4b99c033d7d94647e0d00c2548af1f3bfd11d934ef04c7756c3756c4abb76e2262a9399;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fe3187d70a945108ebb0996cce87ad93d532ebd5ac9bb723ff4966574507bfc2e6c39dc12f3f46d6c6d583f8451d6ae9f61d25e3c8dff6e5c934b1f8909c07ce459e77a499d385235830061c6f1fb3c271608dfda2c24388d264c202acd0e607027;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69e7ba592dc7a31cad375ef53347ab80e882771ba97e236ec46a383e105037656fe71b726312d2832f7891a0ea234654a691f2729fd1e1d70b49ecb15555ac423751677bce5ad1126550401d86d040634e20892f180cdfad20f9c9aeb655e699168f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf659692f5ac2f6737237b2031a2ba3dcaa726a4a7072bbba024b92c4d04d486a0a5d9b3abcc63e9caf6c602811ba15acf0f2d784d1008234fdcd88ddcf8279c12472e838877b894ec6cc5bdfd8f2b81513fcfb7be97273ffbb997cb504c5ab2fb030;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae860e142bb4c1673385a292bda6d8c29faad8a132cc06811b49b981fbcf0282cbd3ed7c770e67b6a662d6148c1a95c8bcffb87355dfae69c3e22ce200030333ba56d84b237ed46142bae9446a96d94a93a77287929f674517a4cca12b44373b0936;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc840b6562df74334a9098eeac15da909cfcc21ac62ef69f3d1e9615182b0cf447e9900c9c649f2b339bc2620be52a619717f5dbfe3423f3ec60528db54d89135bc7d2c2578c2dfea2db65c13ce86061b2cee5cccfbe7c84798cce88f2e80356ddcc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa7fbbd9d1d54ce8f8ecffc741231005d066e1b9f6b15f7b3f3cc032f0e1293f2b5a181bf0f0ef44ee505df1e2aff566af9757cdd351d465f0cf092443efc5633302b239dc26f51c0dbee1727f4a0523ece5381d15085fc5e4ca0556ca4c2ee218b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae73c29151a010f4ec7fe1150e40cb9bf2457f960ebb25adfe03f35d879dcc514bfcb49d02b792c1fcf35da0fe4476c4be42703bb5994fa8e38c0d42a8e07cc11b34cffffb64e969a6cd9d39e1df901dd8ca9ceeea341823d3a21f47fbcaed332c46;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e729b01175075ec3890d53ada01ea98b08a3dea1ab6a4c2a2495861dbdc6601f93789421a6f6c565d8a7aee596d8c34f27b6d1f26ed3edc8a1ce3178122ae5e8485e9b6f9546a3441ea7fc5fa31fc93b61193c4fd64ca9e79ab16665846ae230349;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa61e9a4cd127977605d72b8459ef144b0bf3d812b62e340eae1c2f80fbcba0dc811cf6f364a4e35bcd8a4d9fe96d5632fdd2ca4919e07fd8bce663364be836870ce720f4c8495b7092756c57741a8ea14668a87f79ea406adaf8f6277dd7567957c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36b04046f8eb9de2bdac1b0b04db88bb17ffde7b667fa724008de8d7944c1931167b14aa290ba40355ff8b4fe62224f45a27f66d7588db5a75a9e96e264bf9ebc6c9b4fbedf165d58bc2746935caf62621aaadeca9412de8c6e82eff1a5c5ecad74;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f044e86fd47f8e42d0209fcdc8ddb441327192833f18d65bf915d5c2c344902f1ede4bd38886092d7a9128869048cab67bad03e9bdb1aa12dfb2d34d40fb97df9720dab0db6ac4832e1b67270889fcdef79432e77f6ced0fe0f896ceacd6448ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haed12d9a72350ce0de65eea4a2d80c5ed922fd18c60ad6a5b7e96b83fb557fb0a208e2c2eabbf37185c2e7e846c49bac78efbab8734ce1cde0245b3178f2322c0a44d067fc0d061c6a3facaa1c69aaf1cfaf41c8d8e2ee80e3c1a56578356e2c8aa1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2297cead50ff63826fc34b445f4ff4b5a5154071410deca2f4106def1a3203a18f007781f0883117b8d6971fbaac0dd915601ccb4d836c62516dc1a78d7fc33cecbd06a0e45e68a6d9c3d71bb15e38fcc901cded2561b28c830f1dac8285fe2a6cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca41beded19e32c700a6ed7c5e1bb98019b01d313016a0ca33823adad6fac768728121e480e4ab693162ff45492d1d2983244643a306b69cda173cae5544f2702d52d3bee751a77870c92733a061f737d132a54dbadbf29012b4d88aa1fa0bbdd523;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7db2687db661465e699f80dfadc442584e769339a7cdfe0a8d4f19de560f66af2fc09c712d85941608efa8edc49a73026c32ca3f63cee608b5a0dd5b4772e6a60b80ba853703beb1677f5d578131975b3e5a91bbb73a4c61deee99088b8934207dd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50b8c4d36c3c2feba8afe425efa991f3356f0bf5ae09524261dc6eedc1ab6a5feee9939cd983936f185d299a2a7d8037c0ae294d24abbe355b85250ded158f0a241d92a528930ef851a0e8147e36e5d22bd965501074c6d5eab45cbffae2bcc8c4d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0367309d341637a99e5ec4b548530f5490b544447ebdc6a9705cec5108921d724b6ac7579ced7a1a22c1cfaa0d7cc31cb2979c3ace10ea96080e88ef2baa1acf73e74fe961b392145b132bdccdedf4eb7b984d25e251603194f3959a7f2d77af824;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4d39cf946534750fd071858198b5c63cdc47b724d6a53180978e02ee497dc7ff54dc5826c81700b89bf0a25daa7e5b40b3b27cdc7d4d679aa6a597d871d5a49fcca73c17e0cfea4657c2d1d88c2d3997d771069ea39d41f592fc38cdba761dd78e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76cd907eaa36d0699a62a628889f1301f326c237530ccc42b6a5d960f0b77df08e6ef61e9b0f03ac4920f264107fbbc046f29f3000c558f1d977b8b87e416335a71a07000e13802d49f90dfdf5e43dcd634f6409fe574a51b454c61a95f66242945c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc06d3ca3a8304e248462dbbb23ae4e2d26e75699bba95a4b1babb584edd659d7775ceb381de43a94b6b4dbe395ef9af98016386be96471a5df25728223435ebd107a42c2fb05333057ae7708e20b508463a79d466263178916f99d770c40091efcd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b991fb116d6e578d22b254dee9adb219f82004a1cfd7356bedb8c63af9cb9fd8f891e9c1e516a557d0d444225a2dd9ed064b462e88b55dda859900759cbf4c5a2acfedfd5ed86bf136bafd811758c9a064b04dc5a303dd04a06473d3115a911efa5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bef28ca311f40cda66d053b589d757fa0133226db93a8b77691a3483c9b39a69d80b388ccdbebbbe2bd1bb935e9fe2c3b7ab5482817bda63ce07541f6a12940c7a273d7ce3f44da6f7c2a5a714f999f3819a078b32a67a9895d8384c132e9f3035f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae63f17c21fa95939e2e1536e0368a179c8b56d4af96ba9d2ee036b3ac39f53cfb8ff22977a3d7a4df6656fa7b3d6bc49369f94e44d0dad0c5f57c61aeb7d04c851009fec9242a20998fbd9f856c08d150a5adeb0ca1695fc7762941ed0ad2790d96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf91b4d2624c7d0866f520c9c1f9d853817e95674de33f23f45f52b1c60ff4348413c5b0635e80106a2ff129d10d3572e6ff2a50d8e3c28c395aeea41f2ea4e5bb967b906960386f0ae2c0fee598c9418a3b7b2d25ce069eb79a9e05a39e758c8510d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbfea0a92bf07bb8560e0d485786e38513328d8df6b9a8f3ee905c3337fff02522d011807150577ab1341f0ab274c23fde51b74c99fd5cf947419ea6b4c07c6432be9128b4e6083e91346b8d3e3a84feefe26799c22f866bc45df25fb810ee330b3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h304c4f64b1e84b8ae679d32dabb838779c067a2c3a3a85b9279483a8383c0dc10a03c2e5be2430e72f3a83c16c70fc71b59aeaeaa3540e1a353f45e195c340cc62db250a1d4d1ae80a638ef459838b89eb894f964c1ed2ef9bd192b91d22b1db693c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h651dc249f1d64f56891a81352a7f8e521c5735670d2c3cd83bb90f6d2cb0f665eb3c4ffe037077c3270a316548526b20a2f69191b5afe563ede5c6d97ba513902992cc1bca67d83212a43865d9a423379b99d7a011312dd4df5b2e8eaffd7413c56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cdb45ccefffcf3781ad03a6b0dc89e2b1c2801b1b89099e40470d3d18dc0e3a14799a64509c36cb6e9b1dbe91976a6f3751e1b7d116b3bd6bcac04b0882dea41cde4b31143c3c5c3f07f7d7df3e7c0673768677a64c28c862b8772777daade6604b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he62b8158c9fa67513a26a17474bbb8d9e1d872b8defb41994259c8476d249affa062aee07443a77e3ae970ca3e1c31ec6807d1681e53df39eeaefe16dbfc150b00e078efcd9974d278e5d2ea4bfa7062a7dbaf4e3e9e6e99af9aae86d4a89abcfb48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf34992620a22ada85500da656060c7f81b59487af8c3ca7101bdb6a3b6c8472f4707e6387ddbec70373b1b33f7c225445043d48b6f64bff788472ff017b2e0e4cdf5c5b2fe17e570eadd014a533b1cde84a8ea540a283c0bc7b4703c5d045b4ebbe1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58f7403fade857e0a2f9930c5af580e80f14f2efe8c594c45f0404e4c84ba1f03ecd969760f1cbbbd5d72c3f9b364dead2a4cab7942ea680e2fbf005805b6d3829b5d3a8b824f32eaed29089b22ca62bdff703c16febc6223d036ae14aafa035dd71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d64d2445ed6f577fef549a522efab0b614dfb31c3bd982fe3c26120c6660245cfc21fbf862a860842e28630ea5d33ccb29bd370404fcc5bb588121fe9a9817715759b7f94c9087ef5e8b7d78a7db5293a8aecf9e20e761c56675ee44b66cccc42c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83ae9d601825c7ab9e449a0658561bb807bd5ad26161ce938e04ab2869bed6f22810c66f36b29aabb5db65f3047ef298177d5bf5bd216b7fd4342754ba17542fa8dce148c9afb3bf2646c153520597cb51e169a73e788c1c4a84ebc458f565413816;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h443b142a0caf7ad0c63b2c258ece53251e9a4caf972a6a8897b1a767d6ba4ff66461d11e83e33ee5edec1876e1c0032778670a99d15e7960ee7fdcb2d90ffb9252d5bb0c15dd213c8bcdf8c8ef5be36771ef7fbb1522747fb8b987e3be03a9568740;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63eb028de54102cd64638bc349210c4d6b72940133dcded32ea73c0514c45a72b95bf6aee31213f40e9eed2f456b6a1878f9e33625263390ece9c89129b57874f207e3ff00ecc14963218fe0bd35b768737595411bdcff107d1d44458c8611a60606;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ffcdc2507606d7f2909487b61556df3ec57bae14feb0552e333dbfb0e4604987e631726e63d9c6ad571a616052aa61b1658cbebe88c81f10de71c1ee9aa6233977083ccc63f6a0367cd9154b4babfaa9b52ab1e5606e25dc8c44c049eea51cdb590;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdddf0704e46f4557b5baddc4650e0aa29618f218c0751eb0da6cb959768d30565a01f2371b096901f55f2af4d2b32e9224ac925c5e83f76e19af151bcc66025f88660a895d97958afb9a880f62dba8e597582b4393bd14cc3bde4f101b187aa1932f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf5024936d5dbb3fdf852f61dddf447b847c87ff502f474711942edbd3ea5608ed00d7f09429586d57d97902fc77c0ff3595b3775b37552d383dd27eab6adc031a8fe19dc4cdc9dfa4535a6fd5eab1da5d5e07df3a4f01bb72c6f68ae8a4f7f22094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3af4fdd297f81361977da880bae3af3a01ba2d66861133736941f2098112b0292a97d88e312728740df7086f09529c77cb5c091c15676804d96b9a79b2342c7b6707aed189baadb13da42767700cf5c22ba95215c6022e163056db8f34f0780b9cdf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32487b3b5c3ae8551d1d4e2d98e09f041716bd3a4af362dd8c34ccd05916697ec4da6e5af9b0aaa66228fb357652fd23a2e91e20fa7cb05e968fe13c0aa2e11755f8e67f06a512053e8283e26826e240dda757c7af0bc0a05af8199d79e29cffb351;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7128e43e93154ea56e47a44762ba6b37fc11326be6eb2df006c67338ae4aa9037c8a8763785d58a7a4d5b92cf9df1f3dc3c1c5d1176f91d36c6a99508d19b5de992cb8776bfd7c315957397ff36e972b3b224b9b36f12644b4d6337593d005f5b135;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d1c6e183d53ba4fb07a160505c3e0d364f1840bbfb9a62c79a01ae1739611bcbad787c080d6ed4e35c876c1b385ea204ff1a53c3c059c230a386a8de43362cfeb546961d668d596e2f8058eb5e4f6e3c2f25feed27d35c079bf1f50e5b671ac84fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h355fb32cb6a89865f1cb5875e310c64621597887f9d044765e7ace57306aca8987b1b912f96fba23f4b56e8fe11cfbe1be2eb65c8f125c3baa8d0f12cd08f57ad026d10c43cad4e44054ff36826eb1ea9d680c727c45f89d2a1e20f651f2802614e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a407ca31836fef839999d3f802a45a923d37bd024a09e6ecbd33f6b14115d1040776f17e5c6a46d665ca5caa480eb4ed5f32e574d43c16cb5b0b316d5ff92856fedb85322a8e51baa8dc7732afb0bb01e88ff4a9ba43a437625a6cceea2b894c84d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb3259e0b3a8d2339de9c0a109631a683129759747a340a39380849726ac418bd1539aeed15842fb47d99106c08f37450eb1e8ed3b944c7730864f00ec7e14285187108d6a6aa91280f7052550a1498d4103cfa29c1796159c532ff65b1664030dcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4781aa5ff73992482b4f0549e0039d1b14181ef7ed072179b05f11956a7be2c7e110301125ccf904d8afc8cc7eb1aeac428e1832b920e2ea55ef9a1435309954f66f9cc68647947943975f51a72dd7929ede6e5c0661897ed2b8dd81c98815fd9fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h816813b76dfc1d7db4873840e0a240ee4588b821e4398e53d84ca82bc1627bf97f6f315a588986dbea2cd81bd1b086b342e009e892a2c94d6cc26742ae97404d358bd6ee1064a94da71fd4f4e5f67f1dbc5688316965363392190b5222ac0d4b6a52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff318260cc8d01dc8c9d093306a913e9fbbcfaa1ee59c39c7abef3c1055b858f624f75408a3d8e94a884905fc02f4e2fa10f2b381884c72aed98757631578b1edbc1b4c4cfa79550305a11ac3b01987b6790dc50f9edd1c0557e335c9ee80e6e93fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10853fc1bf4115a4797aa840e6d1b7e4461235a79f95298beacd48dd91e793bcef671ccd913f866386b091eac69abccd489602b9cf2b79f7f8f595f23acd7cb0d9dc0275abfe911bdeb1e8618879f074f0d7127d2c7a8983a9c7a9a54ec0a95a5380;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8aef8d7131498d8f7a1ae8982a63bbba8afd21c370c2440a12a20b6f80440d12dc0082dae94b86b0546157557487c5a5e613262cda16baf3b42443a76ba6a4ec2c4eb803c64bf1ee248edc24519b78e00f115c03b249861d8a8de24a3de9c9964d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc16fe02661db4744364203887c7d3d6f8c4c59ee9643d3c155a9ceadb706ebcad8ecae9df6902ddb4106f66bfc6ea1d0e6de7e477aa13c02440c22251622f2e9acabe5d0c3c2f3f38cc49e6b1009d20933fbeafe3b2c7a1871f2e0e26df3c28044d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5036decca938d23aa954e532de8df26e85d6892068fdc8ad6af6e3f16a998223cf530e3e847a8f8a0aa5163813b8b02a8b772785dc8e194a2acdae7f70473b8d2619916a3d64bdfa594ac59a5be58e0967c393d9c4a19584ffa210320f4070223cf4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4be992ce1502f4dd1732412cc7dcb35bf9607fea906d2599ca395326de64344cc4e98c8509f0ff0f860e141fe4eecd9480b347e287fdf0b9181b056e52f8c07217b3db233cb12986f964dd151a77faf4ea5b5c6222d4b97f17ef9a04459d5b8b06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h578fc85359513220290ed7c4c7ff08c98950383be4eac7dc7189b058efbc50678667ff8dbf2f85bcdc7c00ad994c328d16e2e9b4e38077f73f53661310288673178422020bbeb5b784f8d0d8d39a9a6874e57adcc99e19d27b13ec7c18b99fcdd12c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51ecf1de07b924e4674e3cc3021a7fccf20f69cf0df77b1f35efc49908a93558999bdfe5676d6b7acb6137f13ffd169847e6bccc209a8a1c9d9da60924a5d01ca24a01ec2cb8de527186a64082f73125f14513f33db7cde9e4da20cfd3dd9c15ccf4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e5f9441803e14e9ab4fe16bed204c43a4a16ad52a017be4b14159c3a38b52cc6f81e695a2ce46d950d34743fd69f5c1b0de319aa39f72b3151dd895ac62c0bf16ce0857bc9cb45aa6cf71ea562393fc7beb80a70da63de1f6a01e96dcaba871b881;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5da0ab0f90456fd0646a5194795cd0583f7f37eb5482bbc4443897a09f4dcab9e50975e06f566712db1b7aaf3c4c16dff882ddd6052f3786fb3ebb0c8190dc92c9df7909d055349d049ea5a274411068b6d13450a61a59e40651f613b7b7d6bc6590;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe2b97c5829e88d7e14fe6a7efda2cef67bb0553e348baeb418b5037fe431dfc0d85c3a048983a12523d9f4a050516053bdf04ab97bbf120860382e60a06f1c0bf630371a8618c614eeb5ed7be09ee60c47d451fef945c187521affe680d822c3094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf829227d0c873c002a363637e6ea6266285883b65833a758dfa76590587a1105cf97d3303c52d78de6a0e9013e92e76310df1c38f84cacbab34699ce6f6ddba0b9ddf3e09bec849290f1445ab147ddbd0e04143b8eee675fb68839745542e1611b86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2686b40abacb0836de8dd9c17e7837fabe7cc8a0a0702983824f3e361d613355715c9b0612f4157eaa6ca567a4d472905d0e2a72ed1c185655fc0639eaeaa799a55957be68037a2529b60490be46fceffaa511788578ca77d16f35557f7ae9ea79f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96fc974f94e5fbc2bfb9534eeedc2f24ceef175d878caeb3d78732e7dd6589a7518b349d5bf72ca9113dc6fc6fd9fbad424bb58b5b0cd4f3b45ae8bbd82452e9df7be1059bf524a7e941b40eaecaacd5bd15f3800c1a220e5bd82359e8091508172c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ae7e357433bc52a86840160ec1071c711d6a0de76b740ee0d4dfd56c05a9f8ea2a3f1ef83ae9b653182ddb68daf660a9eeae48e130c62c82d6c65e8f23a0829818606cba71e8783d0de58eb3bca2c70a67574ed0aa073fe076fa40e18a82b9575f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cbe4a9d4c646329e98aced6c13fe76c2996aa72b0619968c97741b78d4f68f142b7d4ed94687c1baa2cf30baa9aaf5c1dc77add3a1e34e351566eefca761198a3198561213444b9ecadf6252321abf2b49a6eabb199b5701832aafa5a5373ac3fe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd788beb034cabf689f2be407bbf9a1b4c236c23f57f3de688d897edba0a12cf0e1ac8bd84ec2b744e33ee3e60c8f3b727d0ecba6e3826d525bb292eb1e6581e48e38dee09c40de864b12e0aec2c2a1543a27b3b8da4c38667b51a353bcf11c523fdd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbf43c4c4a660b551bf87b0edcfceaf2c66197b9e4319e8807c0a275b619990e8b0d04385dc1195779971ee371d08048fe208ad857e6cfbf4ff9acc7443a2bee1a0594eb6918615e7ddbcf438b50a402c16167dffc4009957b301e29491acb0d0650;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5df387cda70dcfc962844c12e5d7873ca6f8e9e78178a73262a97351fc2227b7bf593bdbc2bf04eca2eadf4515bf4ad270243025179d78895a30947c64df18afb5765e4c53b97129d387947f07ce9e80afacc2978f5a4201da9dbf755907a4d619f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h491db0192f3dda824d8e17174a04fe18a255c0ea633ea89d5ce7cfe85e5fbad9108939621b3178389f4b2d1ea13a350de6d8b05de3968c44ce52c3ec7b9020cbb8a2448f211687a687a5d1cccb6e1166150cd37734a871f21ac036001fda3e5a6f3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dc0de5765230baae561e414771291debb73480d67ebf282d0b56e5eb5e08924a90ea8bf43e7ff809c8c2e54c2f7c87530aa1f3afd99dec65752d7ebaa995e59dc59a4eebec3d9c2b2ba7c0dcd3bbf928a1366b1dfd2afe5fa4581fcf6af2c5d0da1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a1ce57cd292976a1d47d2ac8370d8a2dc8db9ef1893df62b80387a5ea32df65b011cea2439e56576e6d4d10b862881fbbf01cab4f2d31be711c769623ff3b7f2f834fac75d3733c92c6b87cfa70e7649b298dff37197a756d9fca4db85378710af6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h478f4fe6f9c6dea17773a1ca22d40258f8ffc8d7516784e99e991ff22a5373b74d2ba7e00341b85ad2d2c1ed0d8ed1ed472fbcfb2199d274dc3f7ff484098b28108bf4c119cbc4fd3650dc5f5f1537a2e72cc028f005af310b1a417058dd9efc24d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93f5aaef9e85593d60510ffaf56e94f4790fcaca73c8a21192a05becbd2d3b50d2872d764ec1312f654685b1af861b4b5646e9b19de49a1da2b96442f0eade7c41cefc4329c93ded52f3224791fc0fb8b043e241b08131d25b71d2b359dc12f68ceb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h469c86da1b0f9f19881511f9502f80169f85efb4f6d9a637be39f98ba0a7bb61a2fc22e3c6747d6474299fff381c8a1d94841e5c8f1ec734029f4251f48297747435e094d441fd406caaa8422dff285b42c6a69d7d0e5318d6e19eb79eed13961a8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ce02a5042d86723ce2b01fde660d41cbf7108cc2ce1e97c340bc37435398a6965a35032583dd736a49ff8acfa04c7cbad38b68cd6dc5bafb93ab07bdd1a61a3717eaf0dd03ecd878c7dba8faeaa9e6207e312147a3e8b32704ae01a04fd0bcbd29b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c50caa6b9a1cd2b106ecaa95c665718e31e5690637a303600b864b3d56c7bb693be4615a387dfcf26f9438c4167fdac6666c3d237118731bfdbfc6b7a9db08de88f8c36cbb6ed8a44066ac38d0b0c83d024845fa668b5daa2ec283f0e8b9d836810;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cbc8fe6a8c40f798c9b821721ada248a25205372315dfbbc0aebeac9fdaba9c917f24471a1500ef44978244cd380f1e2f32896ffd12a988ca63315fb83997e2340acde25b9099d62078d541d4d2b131937d323470592b2394c7ab270f15f8d1a251;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67edfc3cb194b1c988e42783917ca140d62f33a9093efcf66556fbc03b06b26c9b8ccb9556feb4db3c262ffa0395353fe9b492869185384cedee9995dd8c2901e3ac0dee4ef66ce4a7175c5a3512acbf483e5bb9fe793bd7a0dad25e9121dd205fe6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31717059ef630890d05fc0489fba8c53bc31977c080ec9dd34a303b8a2619deb1aa806a1aa85742a05c13877ce78df5ee6b12cda28c00cf6274208a93ceba5cf8f9c311504e3f435af5f67ed9bf590109152e940b6d6bab23e35755981544e5e7d38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0e14e880ffc4749a94a4df659c731ce3b6d2e1ae12ab3de56ff59380cdccbd8637a165da4c0f9a19f316bca25a5237dc7e5623007a0d2b70ea672a6079bcf2edfbfbfc557085ae8aa8e866e6a71b1623b5ca6b4f725e872b6398b3877f14366e5f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc71bdfc942b261b3b3d0daa000e87db1d67a435a9e4468ff72163c01d2a981f9f4e61ea61f88d449c22766d93d4e2912255b42116ac5db5d5dcf9b982da9e16ef552b387efcb97dc11f2ddedd81bb4b10d15399cd30ff3d2c1aab925684a9c09207c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee4e4afd4f1c81b417d58915917bfd85fc6cfbc6d59193a03697add8b356963fda41e11c5d5d26377dcd97b5b1dabddc7240724772768f4a85bc74d2f9f5e002be83bfc947d544304e2d972d6b5029793b2af895afb2162afe58c3d072480578a19b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3b4d1a727dc67c3f4c5c9f0c1ac858442e3fe96d7583681b67aa746d3d1640ad63b176df405d49a7a20391dfa1fcb7f4cce7ae5bebb4b05ad62a3d8868112497915d8909bc032e23b552e1bf5fbf332c805c50356eb4c0eba430c3ddc38d98ab503;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdac61b750f16db24e014052f2306c1d6a421ca1c067991015a540a023e22c347ce2575c849305ccb5b6303ecc45006f6f514ad3d09bdcbacc6bd79a792ae0a44ff53157ccbbe5dbe31ec5b1231d69bf3c09aa3830bd6b97568bce1671a1876c4f35e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d9153d4eaf6afe5c6e8943d67f72f5a1d4682ca022214424708d1f23d74760b8d1f72b0328ddb5117deb821eb6113c24d66d1c41daa31475593828d3d7a7fae4d50bb47051855d5ac2daff67ef24c4d7049a9e0140e893228a4cc7a9b5a2ed154eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4acb8a08ff21cb5d9647e855b6bda0d869ee664a0dc2a5a2ced5348808e764ee56328f3ec5c897c69727b782e0b2f73c551b4cca958dcfc081167d1c847535fbf059e3a2ca28c4eafbb267d9e691de451045aa537cb115323fa410624f4cdf2b2b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1232681a1f04ebe5c2ba172f7e4d778c5bfb1979fda1a2639047a1f73dc555bf785ecce4d85a6f98f8ef961d709ea6e2e3106de6f56907f8dc50726e6d68ce200f83da6eedcb03e9f147e09dc13d03142b0da79705cd66341e902ced9b94afdb2faa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8377ce97036828328d7059b322f0c2c2931958e5c312b4cabcd05a16e5ba3354a30c27edae922b5755b5c9bfe57774c9547dcff3c5b3c98ec14ef8d0adf4095403a4a902f6d5aa916ef7e450e7b9c37dd94de09bc5e695ebf3f032f3873a4a08d51d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecb94bf1723f771f3ae07ca4ed745e5e8d1d368d82cda01c22bf2602fc07a97ad5072d5ded5784ef5ac439a6fe3390f760b338f58f6fb07b33630a98a6949332775fd9ad552eea9547e098bab58cb6fb94ade440c3001e29f0575060cacc047f551b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb844b27191f0faa68ddb7ab226b7ae3cf08901e5915da1e59c17785d9228452aa85aaed6515cd38c38875ddda98ce8a154dd6610d974f1c56a8bed83708d8e24367f532da47af6ff050afe16d1c7a4a6eab8f3dd23198bea76a0a33c73f0fe6a123;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73cb6b9b1782b533829a7e909e875439cce023a7fadbccdfc4454daca03d3b293b08d91f333b0bc2400c1e03e5fdd1ee54b88cd6339ef73b0aa8113a3cb357ecb4b9e2b8fbcf4d78c02cd4771da2f932f392922e13147e6ee0ac567f192744bede3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1849cbeb7ca4c871ba8d89bbfe901f877ef5a86bc2743aff06af3c40b3ccb25761d8af4560a91e8a548a771984ab361f094fe963ed429df39417c0910d60a841ce04cfe5a5c967bef426ed13d64fad876ef60fdda1336f845e4cd48e9835fa592f4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf80c331c37c504719feffc1b9f5d4e579435eef02f053a44d8729a5b1d44ecf6a7a00a122a5cad52336868783460fa276b1b2d65984426c61c05ac3f8a2177435c0700229f678c60f5b8272da75f4343341e6826fa3ab079a2bd0e8a011c3f4c0993;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h516da3d24810e67b05b9a984831380afdb03dee47043d7f22bfa2ffd54e091d8f58ce3f4ba21a4fd1cc826c8e14478c0e6168cf0ddf44b18534e1991fc4f8c4d3ea006c0cb3a0373ed5caf688225f57086e4e399749c02df11f36d385ffcf481c7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76cec989a988e253597961755aa69250f30c1cd5c8d6f76ac209f009c52c8e529a4f3158b8645d72ffffd9a82a354d1dc0f2ce80856266b41ebd07306ba76bdf30f0cc76019ed7c89646a00e70e80e41b997c0ff5a3ce23df340fd8976af24f2d7be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6ace3537444210cc728c990e47101a01b0cd68847cb7873783a6c664734b7ba58f6d01154318c9dac943f7c702c80009f099648aff13e6084b0e6c13c5c1cb55a8e330ec662327c7f5f2bc08608a691c3dc07b491c587577dd5b4c5d57b63fc1a40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha020d2a9db3e2dfe69767cd1299c280eb3e21958b8e8ae149a4f99549f5ee0dcd3a6071a9ebb91454f4ef125a18d9032a0209b80f031064aeed1b835e8a4ee2faaa1ac73bc11096d3086cd752b30b82946c251d5dab3bebf8a9fe541f69d07ff1124;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fc57db8da94c28fb3414cb32f67db7040e286d1e847f58efa4da4a990e4f182000bebea9546fbac2d10a14810a0408fe4696ba09870cd3d70063498e3a6d51db725f794d204647887a1dd79eaaa1ab3508057c3efef4fce3dd0c4e959d2128e67be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3cff9ab9117d5f68a48c8a222d878ef4e0b7b64a44827b96c5dfb6b40c04793e86cf1ac9f10776bb0dccdf55170812bc4acc75f99147b2f45948bfe9a4da7d9b73c6d353ac820daa6b980b3781eb3617a1b28d96cd2156bf56c2fd383c162d1c3d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha10f1a542c50ebb30a52a4f1ebcbfe3455ec5852a3d0dc049556c3ee7d9e29652d435a17fc8eef0ce94f1e8d2f1f6ace8be7b8364612b85d57ce4fe85f7fb8e931ca0a09b7f82474333b36384ced9be96f4203e9c3f677a502257fb94cd2ed3f3d39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h531ea659af6991a3629138e3e8d31a96187d9f3a1d40a904363315ed97da6c4887521cdc5602a7cb6aec706d06ef6ca65b400f1e6339a2d122f722f8ee4fd50b9e3e9a59cf93fb029f774c7b0ddca13627f380d792d9f6307bd9ed331c814a3cbe9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had0cbe2e28d5aa9fbd95b55c212f97dfc61661a2e6afb34a315426fcaed19a8d8dcd7596f79e170fe7b703bd8ce1ff121a17b046a70368e93fa3c78ff0d01d2adc54d143ed42025b6cd6de71c8a929889e559d09d84883d6987c17cb026c2657d57a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf851c9034573f149b671d4a48aab5b7c43540d0a78777d3dee87f1124cb8fa3b84e6557157c902ee5c81c56c176b0052f98ca8712342bd2c2f13b422af65ff9b5b479bd1f9f35536672c8d21a8cd24d3ffd7a3576db9e602677bc3589b200c3463bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42a379eb58adee98fe4d6762e297c5c749e9239d3ecd07c4b8341c0be5627c20a0ca5605ab64feac830ef58e1cf483515c4cb4a287483205510c13160483d28d82fc79b0ab7475807ee96c35356672c40311d2feaae3049b46992aa0e32196b47582;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba6f4f45c8b2815671edd8937b37ab8a34654f158baecf16d535fc8d5ce92b21e130e137e94eeceb09c4823adcb3135ef22dc63be3db0b889c36161482413d603619ed07f1335f44b405adeaf58042d983ceda1be54ee891c1639a96f2b5d0c53e2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcbcb59b43dd6107802e79952e8fade71d13100ad36a4ede1535b597bb6abdbe7f46578775422e23febf7167d00c0de7241cb149966b07458abd21024bef939a22bde482b969d6dcc20c7ee4feb51498fa2da34168e4d87cdd73bf68b011bbb086ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68cd7dcc9c7593456311074edd82b7d499143517f282aec3922f34e2e4dfa0d296b6cc012f51cff0ca8869a1dabf2d84cb7218d4880bd34df29b69270e75b30eaf98e0df740c7810a648fc9c6802bf3a4c33da55ea46185ec1f3bf27e46b4f4485e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd61d4cb8d518cd2d6ec6d2a1e1a60fb807f54c17a99e7b75ed8b48d9532032905706ac6f092cb9524ca54c943b857961a129afe12a235c70f4bfe14c484182cb8d51009875dce4f92fb8a3429ca5692d816e8afdc53fbe17e520e8a3841699ffe80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18e03b8f4562d979327b32f9065ebb005681ff44ff45324451e8c4e2f8c7d08273f6707c3ad05777dd976bc26bdcaa11e59f1431c04d00427a2890d247310124b923fff9210ba22f1146f9dbb674d6ff61c664f05181a79cac1803091d9281a338a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc57752e4248ef9f03a06bb1ed46cd7ebcac36248e525ab2ff5b0ab180d4fc35864f6ec19c5bd32c3165ce75c63f02c178f4a792f24a7be3e07d6c9b2b6e93047355fc9f1e93149af7f88c784b4d451f1e1c70db5b55b6817b7719726ed9d3a8d5174;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc758d50b08798022066e1c8efbb890b3fb7635847b3111769a10bd6e31862568411ce9f4a1de3cd677c3954eb4f9785e9f832b0e7ecce797ee1949e7d5a6b48d5a927e0ed5d75aad4b788e131e29efd47a491b2961991dcae0dcc0fa8631258c1497;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9c74b2270ed73a05e66cb28b2e031cc470d7e2a2bcd8169246ded634e3f254fed448944efe9782b1cf5e8883ea4e7c4f2fe23a089328c6d8620d81dd72aa6fd704651471b86117cb38c52421e3296f9f82d7e535e8b046710381fbab2058cc4e46f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he96cdc83fb61adb15e5c63132142171ce5eb752dbf6687c158b3275b581f0d54af700d498aa6852477c09b7cae36a9fdc47f823ec940d549cda5faccbce5e98898cf20805a77946715ed21f8460f3956e8df300a707287b9779babce556179bc6d73;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1b6c6e78256f8f583736392ce01e4d3545c606f850a18cd1b93aeee60c4ff73780079586db7ce61d8c72289daf07bbb919034b97440ae2fa58811e24a964920cdb216f0f5a24ebbb8c5e9ba203df84aa6021eb708b74dddcd499f1da85f93a37a7f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeed1562b59f64491d53a5d38a022c506c58ab2f3a1a91502e872bf2bfa63296c94df17fa443675bf9ac11a7d2535f88ef81d7f003f2e635cfe2989da0abe2813ba27d9986c7875b4e09f50c6b72b464d962b6419f35666cb3c3e076279792721df9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16abec119872f710fd1c4f0357609b084bb4fa939c6d7228fd13d9487d1555a161aedbc5b82af7ad5c045869d67605443ce60cbcb99111200ace7e97c8f18e7afd232e4b9920267ed6beecaaa9e99224628203fa565fd934ca4aab2b52dbdf9f9af8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1df3417102a67eb20dfc9ed3319d8de5d07e586b5f22dc85b1991f3fb0d6967f8d2b5a746aa8f3d0fe13ecf0abb006f2df3f51c692be13d73d3694b367a62c298a4b26f67d92eef72ca698a1144a600d173aeeb36cd48a58511670d4b4f3e1da383f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b061d5ed503c1a94cabee9df9563ffa42fec820c7cf8d38f71a23039be5bdef76b40529e25359ce07e9699cdf565c2248cba2227f5ee42b62ffb3040a32ce4870952db88cc25276141c8e6fdc5b0261848f2f697cab648b86816d977d86ba8c5674;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37cc5be04672fef2203201e0e9758eac6e28c1189a90295204962e0291677c70e687cc7700a00a1154c2ebc1b0e140d09b67211c165e582f04ff5ae0a289c33820ae4aa9345c9f2a2dffed9a8a07160ebf138376824c26434403ced27a70e5ff1b2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b679a214972205ad93be3bf6afab8d21448a778d35924ce16db15b299c508b36fe71d22f4d48a6df8eb48ff0b624a3572e49919688549cc3257908eb2974e17c22f6c7c4bb856fd66975a7a1c00db9abdc78cd81dc588831c092dc5e6f13c07d89b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h762e0015fa1010b43ac4fa4a4ecd923ce85ab87115246f9378b145d59d7a941f10096a3bebb9d8469a9d965e5c4ef1c6a558dcdef351b82ee056ed58c1a96821a8539717d7089e96ecd79e22a9998b91902c0ada6f2b296be767fc1454212df059c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1ed2e36f8ba9bb367704fa3ab05b4c297bdc5a7ba80cb341c2592f9145e54db88947ebf36523bb4fd8cd300fe6c9de5ed14a9b9eaedc28ed3ffcd1e8a4c715b6f64ed9839e4971ea89f2a7575f80e6d144de2c7b79e06380401458ed3291e05b3e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c8469721cdf3a5301a95f6b6f5aeb60b28c012ee1fa8127a1d48e2ea02a4311d9b0bc8847e68e85c636d0d03a6308d34c696fb7d2a2819a2e55351c4626de47785e1d8128c23b4c6b05b1551a0b674037ad1d9ddbc26b5d10c79c22fe37422730ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5ce600cb8673ccddc2bad9663c7df4e030cbd20540fd05b34693fe4db238ed8bb50171cdfd0b77dfdb59d7e55efb773f76e7233fb33f56cb7a738c1513f7bd8dbf8ee5bb0b2bd323afd688c3e0b061277947577e042864714ff96b161dd74584a64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b4fc6179291fbd204cebd0339cd911f3ae83d8be20a5c1b5beaa8d5006f40ce56391071ba2c656d817cbd0f782b99b4b298607fe8c869f9df74515653da98e4d0cbbc520d1bcae38f4cdce5ed931b7095e761c178f602229039fda925c9f263732d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283136bcb9978ef146ef690359c3097761e78edcc67890da2b194ef2defd4774edd5c55577074bf1d458ed6112a74e299eb213302f668a9cdfefb9aeee827a3fc3af80d16bd3864500df3dd6be16f11f25ba958fabbbbb518b5ebbdcd6ddec374db3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8997add22c360ec9b71336cd3a626deb6c7f445c6ff554a6a54bf0b879f5d0b8c891405233aeaaddcef13893abd80530247bb5a03a3d448ba9ed45daceba80bfa4426fc9ac4ece8d45c86b0f0fc426d3a6deb947395f06447233e3fa486f0b70b2d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h911c23d9c575e3ab233f4b56272b27a33cac8629a685623035de000111fb05c4ade9f65280cc2c16865a6e1762a3a9a5c8714d621943ea37887e678d6d29c436f6930ed71728001a873603fd4fa1da61b19b6333c94c2e305c7d7a5b08f66329b9dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4a7959f55d9742aebd8fec44996b7bb2682e2fcbdeb0f034c37b5896e33091104aa48ce3635475e0ced43a1066a9fda259a1993eda9613e7802fc51a3e441b807365843754fcd478c0bf4f95182ce4668698910a76c1ae9cff67a85517c2dbf2d05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564c4b34394bbfab678622561a7a08d29d48a9249b3009953b2ada0395a0e8ad24c4553fbf96365ab935a6d4b743e3c740086bf50857e15402e8afa9a91a4c3ac3be530f5484c7dc0253ca0ccdbe1746f676daad6be401e82f46b3dd0885f158544d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf287fba1caa763736541e0c58c641d7ef5abae132ac3e52056fd46459dd57c5890de711726c0f6b3ac53a054488b5103db81b141aa3f7f00bff57d6af9285aaf434a10e07a2519aabc1ee29022ca31a9347f2f449954b6e8fe098128016a3c8f17b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14a8059209611d073f05fe04fdb2f6e42eee8c8370445d5ce768befe9352ad445d860bc03997392abca0d35e98804eb52ed6bf0cef5839a4cad4bcfc65d38a82269b132eda581e07fb488be840bb111e7322242e976a6369c4be8eeba90f74ffb92b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81765cb6b7d2f363cdf186356faaa82984771a5ed9c8280f405a526de0a90e420aee69d33b1bd31ce1f35f6320c20ccf4ec59ed5365be9ac1498dee96dd21aa5bfcfd9aff184d27d555e5c6503117680b692d9989386bb6612dada601786021526;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc12fcaff262bdf435367a93b140db0e5e1b02a782fbc6c8fbcb2e0c74f10be48537349312b84b6091b3c2b6c073cc8b26d747b0666b5c7a4604e9161fcaa335a53be4129705e556fbf82ddc9ede94f664a1ce4ba26011a7864cd930cbf6162575832;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h393723874322e946325ebe56c8f06ca1e40e0e7241bd10fac78c1e9f5b10307b03a3969878f9cf4f352e7c9c6f6d12adf444397e4590f797b280a0e5152b4d3fdb065e439099227c88e161beb913881c19555cc613320ae76e55a1582bf2e01edccc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2be64d004b0695f64bc692bbb9f9b3290e4ea18f7f6c088b239f1414144b508af6cf3e220668c4f43a4eae5af4091621fa1060c31cda2dfcd840d93c40770cb4fa1f100cfb08602815a87c0bd69e1a8a479a9024aea44e7d251ccd2d83c0802ac655;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9537cd2207b9d059c32e27a5ffa3d7f04a7c8fc7f1789c55475d5c7a349c13b20d89ab0812f406df7877a00cbb21adaec68ab82412dcf414f1ef897105c47e4f28ddf7223594ac49d219078e6d1135c3120e9c06fb235938b775852e3442172505e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha257a2e9c478400703f06ed78c79e45ef149141b805a27a5e31f06cfe9ee29d6b1ad2d4183c2f46472001fd50378dcb0d963359bafcc9519e9be90ad3318f9bf896f099c3f4d28e3678a177dd4e8f6297b93145793ea6124fd64e3ebedb6708136a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51d754d235043ab3d47c7c9b1fc9fd17b395580fd194b45f5cafd080c523598765640a1002dc0cdc38a10dec0b38d945f3e028295becbb82dbfbe9dd87bac84b7ca6768a3c762bd9732cd3aa2e91e17d951d90a1c38ba56e73ff0eed77e545051499;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab96c5abd044da677a651d3210d58acd99aea2372b105943fd420ce6c83a541d3106320dd3bdb34fbcf521faca5eff9daec5140b0db2204f3c5ec2c9be56b8a1f7a573a2f24591523ac09bc068325930abe217e9fb6662307a665acda2f55a7b1f97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68373b28ea37d0f4be4f66c9116b82f6be0c76b7189585d64f7259678bd23aea4bc9c112e2913b861028970290a74e92ed01f449915ed85a674a30f9a5c2603c470284678c539ef9a352ec98a7e6f1979aa06691bc7cc0494163fc79720c5602e059;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b419d2c42bb500ae0b06b095b7284c8c4982d71e041f2d204cef5cedd893d66667425030c0a62c70d5cc7d6348a1cec4e30227f552bb0ac43b1b597a59e5eb3f1c0c89ae371c654d464da38d831a409de868d7bf9bad8f488af953d67a584f6f737;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecb1bc5ec229c3dee50b179a29f0cb1a13be42ffa18ca83917a28237e7c2abcfd34df860e31e3c47bdfcc133a50548b05d1f58ec1fa1a9820cc94754298d94bb083cccd4d1aee461e9c28280a3614fcf419f6f6aec08fe3b4dcc6f795556eb3b284d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc6a333d896ba21ae39544b6b8c736c0016ea9d24e8157afc15ca9f84ca050949dc86c6a7e5b77ae026b1a376797fdc3f19bcce8ee7e730a796c4a54987dd73aad45c8b14208b231a053d5ab6aa369ecea87d7444f4040cd3a0f8b89482208e50a4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8fbf49511c996f079ef8106e2449148ea5811a46e7663a86b1ee3c5b0780a0e15f4c53883b4d76faa4cb895cd0eea85f98b347c412d7ebe59856853a17abeeb1319e1035869dc5731e8c558a9c3146b6d19d655dba8c91799a7cb76170380585efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49615362d1c0d63e300b35bbe6f1092d43c76b26f3c8579411da52c4a87a102243dd61b4ede771c26510510a3241b2e5b16fdecff380fe7a513b1aec896a2ce1bcf4e0fec7243bb489767af81b4f6f1c71c97eb2436c7ca62951458d2b80a6f21682;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5234241bddd0739fc1c773da6c6fa603b99d43da3133071a0f005e0cf641f08e8fd754d656e3fb2362ebac0352a3ee22552041a05b7726fb94c08edcabdbae25c2cd0afb3254827c9d528324a803895ad74a2c60be828a8790d51955130efe191cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd00fd5d9de6236ee369059030e680e69eadc011518e0cbb7bf22dbd04a81de388c119085043dcda37089e35c56b51e599e8956632a3ffd2668642c10bca397ff4183323b1910ad135339ef513c809dc19de89a0d3cf89e37ab37d983182908a12d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e741f7d0616cd57b2caee3c8f182347b0d7a1291c7eca86464cda3d687606f984b26c95e15dd6d859f532dc4403c781a470e6eca75122442c783c6a299eb4f587c9519de957190afa096c1eef7b7c58907848c42259aeb2c388953d4a65d308b85e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he47e98e1139ecc6da30319d6a53b7777b741846130266e13fe9b4ce207c971ec5730142a2b294750df75ba7076826830f124ca60685e9dc26002a1e94c6982e5ed40d4b5221e1d76304da33a7650d00282c6aa7d3ebc028cf86ac83deb2ccdb667d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebe5bc8ced212c06e1893585edb58836d8eed376e50530c89a9fe468a0b61144177d1e8c019ccb577c4df11ed6e0fdf9e91262302682f7f6a973d218ed6db3051537238862116e836d0ad24760da67067ecc1259a73bd2e22a0120310e8aaf66cda9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f11054e386fa4f36ae78f190ccdfa7adc453ed58e25dbceb44b92fb980df8edb6f0a6cee221616355bb56fc665802beb1a222377c526644eb1449143d138c91539e7eda74013c49d48c2f1383c21f218becbf88a81fff22a2aac1466da145495691;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fe3ffd66c9859956cf53c80fceeac52345eb4eb46beb8c5c18488652a63650b98bdd457296e798c8abbb60bb25eb3bfc8b8f1a989a0c2ddec81a563d9fa4292160aa4fd6c01bdbb26abe88032482902f6821f4c88fead94ea7dab12754e3b8f5fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h718ab6ddd522de55712541a8ac08c81b6b164be0cc57f00eb4ac198a685f69e150268ffd330c9ca2f8b791720abaef48496730aedd408b4ccc637ad05f29423434346ff3aa466e58872a3be4b1c5bfb48ad2a2524453c9f29392d25bbcebe63f550d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86ef757a6ad0baeb21de5e96a202b2ee5dbef413bb413059f4b5c5cec0edcdbf35f47c0dcdd0f98cbc309059b049a810e2b8ebe06e5f313f4f7c59d85f2154babaa64c2c37a11b9c0e6be35558e381ad889727f909a6b45985790f9a2b39fea284dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafa4a550ef912e8a12c025329f19d22b8eb3e54eaafe2efd35d4160c49028a4a7c340e405341207ed8e56fe6b73bb4ff52d3234ca2303bb518a13ea8e61fbf22a30fca792ae2494fc695181af1d6f870610269ceca17b81142b1128d685cfa656355;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c8f8eb870bd85e3a965dc84838301fc292dd1586e9afc2544fed43d76ed2489b1281d1b4ee5bd1848f8056d33185bb037aa768ffc61d000102bcf676e2ce2516628fb5a8b0aa5f2fac55d635a69a0b38bc6d720eaf75aa067586a2aa27371ba0914;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf53be772598ede106ae6850ef9e54a370aeb52fb8b3d476d528482bdef7d663f48ef55a03028a6d2633c7b69d72b0bb40280307be495ebef430024f6bcf8ef1a602da40d9fdd5ced6b24d5f16d745a8f567bac09fb3e464ff214846a552c440ef44a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb426b6285135f55e8f9c9a062817ef1b1242ce49f879fadb689ce4308d8ee4732cb9555b3719696295ad28f0996e58c307552fc71e1f19cfa3984832c55d44406aee6c85712351f88c19fe53d65c8b582e4dd4f5af1ec7105f698b47209729013014;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ae2bac7bc7bad2714ef2240b1a93ce2f1318ea2c12f7735457445319fc698ab599dc8687b0fdd66b6ab41bc88f089dd3bedbd5f5d25dac7838d930eaaf713a07df43b1bc4b4aff88f83f98dde12389cec64d57d4201a915f1b3cf75792065b9414c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e401d54a7ceffdda90b7a15f34015a0462161dac3f2529c5c3c10123e2fd950f6f6c9d65cc0ead8ee36b89f67eaa2317fae53e05a5d804159b996e5d791ed059e8137c24c548e14b7334feee0f10c7ca1370543ddbd6d9edabe0639c0b1379f75ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1556b50b3b731bc63dad84a6f5469b6ee58910a1a7f68e374c4be2f2658a0df2fd17c0af21b97c93a3d0940c146c47db2c0da92a13a5b8c0516bdf52db7576def82fc975a51c30ee8b3ab83f28a8d3d2a9fd9e1cb8f8a69585b02ced49ca75429e8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he34d159ab0494b0890cc8fd338794d3bc4af5c180a74f1a77e1f39cb21f00a3d1ba3d3f6b63c3372a5e98d5a10d4cede79cde6d34c3a82a6b8e6233b07800ac728dd0d4f53e541a2ec37cd58f055a4b944cf2da853096889a8169cacc96bbb1a0adf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3388445158d6dee87de7ba454984b2f5dcf98a26aee061fe9e98a337b13c49c0b30c07c8331c47ced9586d40c4075e5c69108a18058ce1fa2a85b28c51da2fd1c5e1ac1be8d17a96d3fcb5994bd51285ed7dd3b960da0672c7b066a3d449e55a6267;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6d5220b00268f67c54f73ea2e142cda3e5b3a38755f639e9fbe33814279fe6b0a840abc04a11544f07dcb760b3a9dd04166f8224ebf76f7528a2f516ab718081dcecbab340d21918c12ada2321b24a238b27272d9cff82a01feccc79ecf856b0782;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb13982b39b47cd6d780d582d03610415345311f172ccdd1423c8c8c56a299599c654bef2f0a76bc9a21ce00e0a64ef9787762a013007a3f90ad50af5a8c857b73789e520608c29b77326f5c105261b0faf8e23306fafcfd02d5dd359dc35957abf09;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha844928de646a05bfad444cd8ff4597c9b10e4c20425c9fdf0ed02dfb161773f6e4a7e9e807292d7adcf61971facd2300b7518c7df9f76ec3b09942888907da2e0943003f50aa4095fc5df45bbc78efc5e93392d2ef5c2d80511effdf2fc712fffb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ad33b9e7b8abacefc3ccc084f69543c5c7c6f8c7af1ef4a7c8471f00dc25a644f1e3a0a801b71cc5d478353b1faaf85d156bafca1b53ab556a761176bc6a3a6db9fff22619903601da70daf396de0d83791237af4c6e47f0684078b94f349e12f12;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70e9268f6ad49366c937abb801f247e8989cd45da229e4c3ac3628dd79e6682eb8d83e1f2c3dc1eac48f22e7ebc49f3cdd23c32288ed14f74905a56a0967197f547bef7bc1a6e229479a46ffc4aa29d20dff4221785a35591e7e36b698e22b7218f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h498811da4bee5bdc09bb3fc93aac3462822948842c3577b3aa85a5b63ef425c7809ea62b245050427880b647cf34076f739e45316232de9fb1dfcaaea58023f1165ec9d70a9d21c73e3cc5d00e76faad2638e20cf5c62d6f2c7ff06be621793aa071;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d60cd501353cd24012f29c4fac621a6d4b5f45496b2e81fe50855a33e2b2f66b6346c914e1562d38d59a68319b40e3eb75561ba7e62f5d27417506c5ecd8e6d0888e05c2119cbdaf90c1a3e696feee78ca003dad11b6a14a1df786adf26396bede8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb90dd88852686b418e034b19ccf9f0c8fec21bbcafd68e7590eec0635ab07eadc98b522392f71a292e87685946a242a7e52edc3ef2e04008e07f0ec4de8a09ea66e9028fa7a01879c7d4cd17e5fad544c4d41cd673b3891b9aa9113d10238995721;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96bc1592a3543aa9a21969e2cdea72e181e3b931d111a482e413620be2b6fd4ace5bc993261fde030b3595f04871ef81c10ea77fa9bf5d53abedbb65fdbd507e33426a3521780ae446cd53ad11b3f02fa66601e0732b44da9fecbb6fd5d4874e7537;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefdeff22173b63e9e07a2c5449566d7cf996497b9c37cb1d2b06a09e1a69dece51f9fc1517cf72a997578438b63096fed7d80a665598b9e37a41766857c02f868ad0a707fb92a1c91ffe3d6b6dfed3af91f6dba8937eb9b5ea4b4b8997224a7ac58b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h807763568525d755537805dded1a333e1cc6fbe1685a3efd57643d39ed39d06e9120f9c3d60b197bc1157b0a3696c5465db181c3ea9d9dcd476a50d43c51d9fd978b99ca6d4ec55908db4d9a10e91d300e509640abe6a315f84712c8c9606f3280;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc92c3fdeed7e39c65e7c8b5b558f307cddcaa1b60752023475fa2904b770d99d7d1dbb7d02b4efb014eef6dd03f2428f315cf815ece940041acdc06542a15380abce3c579688c9f4570a3f5bb3dbc9311fa4de9301b5ec7bfe3ae10fb7d7e5f631f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d99360a9ce4a37bead7eeb7a942e6068a9d2a58d60920a51a6023f68bc2490197c613f1253b1492cf65eccb31688d209cf139a58a00f504bcc824dc9e8d892b0783a30378980106ef6b987e0cb5db884d097abc6242d6a5c9483e7a9df97c452c3c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha00512793ae558a97b36ab746b35f9d2e4fea9205f956b45b4df77197fdf33c506bb3bc2e9428d790b256e4031788d56f630667f9b57d097efa085cd03e3115fe33a6b98e8890053ded3ba56a69f784357cc2e71641121f38cfd7ab3ee20a1a516d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h748c8d4864a1d8ae2eb5148d29b593bd4e7109221192b6271a5bf782d918d57a5eacc825b296eaf9a8fa2c0e2358e4828d9ea53cacbb34bbe709b4566b8cf0d78f551225045663cc045ef27a45fb06f5305d50bc2eaeb499cb2ae37b4604a416c914;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc65efbfa00a4669d98d99f75b873ff09d745a696c92e7964e18eeb74bd7271d9f7fea71f36a0141e4ab4d391ad565fa6d35627e205a04c7e375dd11f033f82c2f88c1e8833eb40801d8263fa34c9c994cb4afe9f5c0b3a997662e920f5b982a19245;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe248d090919fc626c73d7d2ad6abbf97fa87c663b89789350620806af4a2b489db8f160d6f3d777cba8fc0f8f5e21096df98284c6b68a42303d92c03e4ef428b0ebbba47049900370f486048ea126efb99423bf42331800c4e2d5eb1738144f0b60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37b9b4f85e65dd937dbd98f62e5d9af4f16b587f3e93e1b2b42bb3de0ae9e60b7ca2ecc5c88316982a81aca4bf0242776cf94e769afb7d33c20dc0fb3f45b0d0e217894d5188b281aa487bef6fd17ee01816ea1eca9903c1ecb0d57ed0b4d2dd592;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5786d58c6ebb3d30036252c18a4fa6daf58a843ac4734fab9c9570be5601c8850e9c2c77a44b656aec24e2e970e3bc4b149300e2e81b58d32806a162560885ad033eb129584983073a720a1d0cc4cb0a15bb122f21fbaf8ef5d273fdba359860e3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h931dfceafba3a24304d7707623a2a6d636fae50bb5224e9a2ee8ed849ef5421457518f26d9fc1f0b580119ce9c71f05799f59d29f83e7576480a914ed794a8707ded5a7c4eb2b8cf7ba72883f9435cc12097c7acd27b777f80f9efebaac584a5b237;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37279b9c0a14dbf26df9a20c03c7d99478c8198c2415f35efddf612bad4616486f1973a8e7bd828bd1ba9df0b6de114b79c92e7733c351a241887c1b0fb8a3d954d8efdeea9f07bd647bfb7bdfc60f14a6d617a88996fee930f447d3cda72f381de0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h683c6be833c48838562ba7823a62752cb4cc523ac6229d48e840fab7a554c077d26cdd86db85c42419fa7707257a30808635cceafe0e740d4e1b49173af2e248be419e98a5a92d45ea37646306ba78873c46d38ddebd3def3901790c93141f1f1e34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcea68ca7dd07d677573b1befebfaccc4fb62c5b03ddb12a4b3a7992c8a2285c9bd02cb5f3fd3a4c479b90a38448af0f20cc509b38bc8fea10810a01c58d3320110a33a7955153e7635a19289a6ff32ea4a47bfb2386ee53a3c4a55d548b22a14dde4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb54b9bad94ac7d6cc0e221f0b7e5043bb5d5ccf5215cdc3818a7f55363023eda5310012a820252989c647b50ce3ae27f1db2dc65cde0afe27c0b06a8bd770c3ca4c1781a66be0820ea598353774fb2f871c435fbebfe8e86329dbd1774d01ce1828;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had3026bc168ae53af0e4624b27b980b63eeeae5d17dc20df2f86856e0de0199e456563c92a989eb450671cc6538f77ba286c5b8a5b44e3fa4b562035161ec3b5ef20a6714de29ecffd9799e851b847ff610c69b4a94ab9b3434296b350da46933c7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6d2c9af9c599d8ab60f35eb5cea1cfb3379f6e689cc9825d5b04db6c365383858244d4081f5a7777ad1b65156058cb23b8cb23fd95724e61e3bfccf2cdea7b2fa249fe9e534d429fb3c335ce7e74ea27448edf732107b58ef4f1deaa61626f33f92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d7f0c805e4a595ff99a32252b58616e7ec049b7eade42efc2788a100438ca12c2700009ec18650d98a3f8964ec6296d82f80a24cd83de92837c1f5441f8efd6763822ce73b616ea0c1922a1a51848b5b47f2c3711ff50a4b76359bb4383b2a2bf50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93e825b9ea3a83c0832de9da4c97c32af69e5c964330ddcb3de020829e9bcce489f8c9b3380fd98790003a99b82e9000f55018fd55a331ea47969004a331d07ce11f5a7d9c6143bbf1d7ec2158d83850771584858679c9b5c56addab16daff2ad829;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5bf50cf304622b6e2fc6cc954518a880e6311576650fb7160fbbc4026082cf52ee7593e903c34d60dab779ecc16ad670977d7b4459bae52f36c1e5646da4691623eb7265be49cfac1197fff56b1cee2bdf8f6cdaffa7311442c74e4c1bfbe3f35c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a0e70bad4d2f923975bf43428950fdca13b181f6a89f50e430b7cc7bbdcf8720efa97a0781c1ce9d9e690ddac7ab7652de87ee234721c422ac5ff597e9aee3620e48adc2c317723b1d1f00f323e436ba3708a5d4922ab7ded26cee0e8bd9a6bb507;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb30484d2160f92991ae3a2b6efe3e16b78123c79dd7714e708d52326424651719c451a3a10899244d13f9d9bc81a0ff7dd63b05218e6405e9bbeecd70b762f67bac480593535c529c4cab2031bd66c7c9dbf28a7dc8e9211f5dc1589024d4a54421;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38276af43f231583f6900b22f694285be868a5765af202ae7bc24e48ead32f812fb4f0f233200054b05ad51c0e7fdbab93620ac840cb277e3e303c23f2c7abe98165b50218c18da1b78c3ea9fcf37eae4e5d418b0e0d47e7c47228cb2ddecb7fce3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfae69c7afa9419f5b87fd691fe0726999773cb070d365b6094a486b09965f691579e1618243f89aeac272a1a2cad9a59356d17d42ecbd4a37ba7d9c401208edc723e792014c6367a11039387ecae7d49628ec7407eeb59eba0a70c4b3ec7b6576f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce3021c022b83c23e9fe8da61f55a3fc57e82052fc039a5d015784360ad7f31102ff203641bece5772638e19cb8581d4aaabd9fbc444f1a33c121de193e85f85079d17fa14281d73551c5b48094721365dc9cadcc9c33483db632f6dbe6373a0016a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f3118e3890577bb673834278d5ca33bd28df5c0ee740737a773fe29b8d12e438b52bbe20eaba4c2d14df4108b25924a284c05ae576827f4fe3c57172c147acf88e708183e9af13688a5a1ce566a8f5e19da9a4d34fe77bc84a9dfabaa97f7792836;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ad5b9eafb9793c8b8856b53257645b5f8be985735686be476693db8d46f43e2196949e76557dab31f18ea69a15e77fd4137c06df2407b04b6d3dd11901bb745ccae3573b2043aeaadcfc4da0eacd2f9eda4f8ceeaf9d639034ebf95d5ff233cef3c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha34d99704800680a139a50e989e601f331c46250cf55d138aa3c42276183ee18680e625b387320afec80fa3b152889ad68bb8964e4e48fced26ffca1635bd599b17d3c92b818180687f0bbd376ab71899b606dafb013b0ac95a392ac9322cdab08c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7b898cfeb2d18cfbd13598f4a42d164bcad11a15c6dcdfab47d2c416fd95ba1d80bbf05ffd74667669ec65180a5b9003eecea9147d349af0606d0d0a14ed994ad391084ac86bf8e26ef4532c0ba31228b3b8a2aac70873aa2944fad3e92bee049a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c8aadcbfb2e74525305d3c220696f1f6f588ae371ebd2a47969c61cc024359e58d0ddb2c1f29d78bc01dc6c480ac2492f5fbf6311a656cb529fe1f752e58245799a89f6a86e4833eb841ed047faacc0364e22eab2851442bdd5b7da85f1c06218c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b53cde889568525e5fef54d4d2bdc0b371ad01f74f4b89f4c21ef703e5f62f2cc29d2b2699a8f59bf3b274b781596f5bfc5eea422c96e334149c6e7ff69f57c32922c6d7f54c50e7ce89d36bcab192bd31db7ed0a5e5447c75050c5212b40049c76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68c0b6733ff65ec5dd55768da0882befc69310bf0723f94b8fb03cf1bda6a7f26644ff52c1380e774333600f5d483c678a2991ec194882c17d1a4b44a86aa13fbf0eda658b30fe03a556e0f2786ce856b11f78a9401f98105ccc5a45d1543e0af0bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h376ca6c2479b3faa77849ca78fd4fe52b123b2e45f9a29b24ee68af115fb46b46d352f2b206bc8783fe6d6d59f530b2585c916f34b5a0ccb11c7ed6217a3881bac59b13fbc6c8408198fe57a0ba88664aac1affeeed0184830ce56df22da4887aa05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee89969bdc7dce6bcbe4c95e1d2fe94c7bee3f8df699b24d984ae67d9399063abed7cafe588c4d0446c684ce5fb31a46eccf7122abe5b90df853a49c40c6f32649295b967cb6ef07182854ac640dc59ba0e26b7f9e09578a67ba86f1e32fa8bc3b38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ae4e10fb0bf6553123490d991fb03035da1061d59d6f7a867e1f808b21c1fffee9acd5174ff619c165a33b27163dd21564510c9097deb80940de9491cf5bc37c0732401b074cebcc9c3abe98c9365ed8414c729ee0cbfb31d230300954c502399ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd699bd257b2cad05b3560408b774d8288c0888ec4f5ca8cdc8fc6bab99988f85e2ee9fd3b24f786d41a6c145dfc3046b0d85cc1a3a77334cc66255289edee9f5d9b0f56f7a7946f7633c15a33d0aedfd0ec51b5b43a7b4cbf2e29a76f2af9dcf4a55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8593a67f56d3b11459605ca994240df95c46fd3ace5e0392f37ef3e74893e66ed7836338d34538fb3ae35881e596d605fa0f3104f47bb93905b7aaa19a5f711db8776f96c75ba7a3378e0afebafb66fe430a985c5bf0452a37e5fc42fcf96e104b49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h688be7027d0949d23064d1809401939693aa86b0ffd0782a148093cf572dba22781bd3ad736938b348fffc98f176a8557a0fdb3080727645e92d2e77781ab28fd8a5a504fc4728a030d1b25022a65ca7f2c9a0f7c28e8d772c6fe344a5ed0f0408cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f4217f619796e4afa87dc2308bd80b5c40ff595eb047ff76251cc1b1c3f1c57f01ccdbffad71ee88a9a71d5b016cb79672a68321095e9c03c3e9f54ade92461fcf93c4d73fbc5099b3d3d0e17c2d340a4a3c2bba52180a0296a0a4079aac595b46;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbae0e213a2700abd7391c5a5cccf41c6969e61a08c11106b0a733da5f5e33cb330b8ffcb5c94044e2a12bce80b994496711df31333b2026a0a80ace2e7348adb820de361bb799ccde2b436cd7f094c6b661d66919c90ab00eb50cade8565b3b0e47a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h950c41e9121b74df5a2bea8ac3fda2c949f3070b8b6ce3b3db84c897468d4a0fd0b2b26b9ed945c5b83735cf9964e5897004c0040264a091f84b9dd5564abfd274f684ad98117350facf4edd2f2454c6e309b3300fdaa6f8191c2ddd0cd560b4eef8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbf949bbdece54fdb88e4878bfa76487cc42c53f90a8c34051e2ae68018082c378aa2acb9a3b8ca01ee1cdc69b2fb0c82d627d05507122f1df9c4a4a237d2437762a74e82b0f937c2a42baa34530003a07923e27448c2c1ee844ee44f85b319c06d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h948470fb1ff6978492d4a29c1cc671b0330ec4e59d71015f6b8cc9fb59dff4b4e759e8ba7557224f0b4e09e9a68f76839676ce14e19192660f4b17d4612c4a8c5b36912fb20d6647f2a739ff3cb60753d5c7641a2fe7a52fd4eee0b8cdacb28ab1db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ed6bdf5f4e7eb9221ff0f65c573fba8ce6b808b4e59e6bbdf4b333e71ce5fbc018ff17fceb0965d1212804d8d44cf84a8c7fbafe64a15ef030e89c9e8009fc2c6bc187c236cc97bafd392bb26f2a7632d4fb8b1b94e7dd9cf7dd85436b74692fa45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33c420de43018994c634eb52bc43e111e0eda88aaf379b143588ec07ccd1747d7691764fc95c5851fe32614b0df5f43cac0a6a3584c1f0f6d99a39bea860d2c0cbd39b1252781a937c4343dc1fdb5e3f0a0e5244e7b4b6f64d8c6c21b8266b557e79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h485527f1e4f2267bef7dff35a763974c5d289ac1d6d19a337a033a26cef95af53d65d28129be38982d9c9d614bcfa64d4153ad7b942276dfd4f5844302272e1af5ee0a01510293a3f394f6f0b8a2af8775a89c87abe882036f930e0fd995e03c209f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1766e9d3479c52b99c5b6c67a124ba1dfc2585806cac2d9248b5beee26fd10d52dd9d9b5143902620b0863d2285799881f28875891c40f786169b78cd5c0a410b564501eaf1f46c1360ff845301e3f9b4836af88ba2c22a4a1be081ffd03faf9fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h808d35bc7d8877dd1f9cb7f41305d7672f15bcd201f98e73d13dd75a4830585a2ccf8066082482f0bb55db71444971c3dc4c3bb6d6949763fe9b5812e78325fdc5a1e8064b64b093ec9ad95479662a4c819e78c921b0b593d2f3e9b48d5a71c54f4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99db136c0caade18e9e87217046da4be70f2a35ca1ab4166feae4b28cdf342b8b63e25353d13f080e7cb64256078534600f6da29edbb428d19652d2857ecec1228fe05b2a712760ae5b795d5b72ac478fa20c4d34cf35a106322ab461d2a2ba25f99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ba830c814ba287a3c4198a924eee328e3d836047967955a8972118777e608be2a9b46e01144154cfc28df51b788ff85141d58e37515c31f08d6613afeac401588ed3b19d6ac418df453c318e6dcb7d2e3de202d78e555dc24f3b4a921ce695a02c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18a5c1908159eeaebac7afb4051a832e1e8f599b0f3edcaa0358f2a68fd2c3fe74a22265cf4975f005f97f72547e5f5cb7d9bfcedd46caba040ab6a7dfd85d7ba4ac8ceab1c342b80748f2cbb0a48fcd30ed4b07265fc6236acd1e7fffb8dc85c0b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96612d9ea8fdcb7a2cc8cab16a85787c66e436e1b8ca1a0b8ca30ab6cbc06c262e6f2ee9f78bf7663309b6ad24296fff6713a69935d4c71a3d2bc98322ac87b82f2e90dc5d92bf0b355371506a2f1a69b3db0ab1e75f705f33207a32203604ce39cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he19149184092be2d9a73911e2420c09b16913543afccaca943d78275d5f508903ea7935a7947ef010903662d029290d648a0361bee62ee75fe8124bbd5c7e15946d814a407129cee7c3fe9597be17d0b969e334b96c18ff296bfc0484272ec9fc838;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb15155c5bffe3174fb5e9e300e893136dacb956a242605187bf8c4c8c6da0d0203c3b31fef265e66df40a75c176cc6a2c2630d6a83a4ed155f613421293034e5e98345a23f53823705b28ceed454df6d5b165f0ed0ff17ca64ebbbe92b6d1929def;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ae5f8a60e1a92b629ec9f660294c5e802a488212ceeda4765a856089822ca084c26bbf3b01efb8a97aec5875a9e6b2ddef598c0f9178b308a359c0d4047515a56341c364178b185d6a2a4c358f0d5dd89507b8a16dca05a2b930a270c97d96f85ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4076132db33088da5ecf9bab3439f8efaa78ef9ac6b030441c737d6f387ceeed69c1b6d3fc864db43b2b879212bba62a9b2c49bb71ef2dd875e7fe285301363a6b16e072c6846c3ef5e8170e43b883beea9a47b053b4ebfd1fcd5268d38f9c9e299;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6948c0b8571ad4378b8607f3cb7b81d0dba80b8e6449c29d3d79dd35985f360d92ef8b3d6377ef14565eaf72e6d60d263bc60c68c9a9c0e9b23f540a1c56e1d38d2a81e8c6438f967801cff86bfafddffbce50ad28ddcdb5dbbb4f3bc4a17f61a01a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfb1f7009552bfe7edfddfec3e3d1b5b6863dc66a0d5c28e75d2995517da775f2bdfa0c529fc14fe4a85a20e17e4752acd7890b4c0b4d5e48e19bcff2e44dcc8a7187be736ad811519b792b69990fb3df8f7b2b1d5cfb166b11dd8eb3d2917fc6223;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf1f32925071855abe8176f0f8f219ca02a75ac697b3092c77951c80bb15fc7225bc02f629bad44fd18c1d2a123a62326548953414f8cd894d087f4c3fffc2a00bd76b3a93689f38ba355ceaa96a09dc8a83c972f53cd219980dd7f4a151cd948ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac1fdc013ec0340dfcd28649bc08279b0e58d04d205b8401bc67b17ea011bc2b59592114d3973e7e3e87b90c95fa56bdfb25dfa891eca292f7cb2d1a4e4801e7e3b058b3fd6ddd34025c656ece0d074f84277fe048a7e55fefe41106b8cb2eaaf144;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8a15db4d1a3255c400c40912a978a6a03f92e7af12396d9d3656c0b68f2e5b3e6ecdc1a05e19294fec2b44eda5ae28037b5a36eb1086ce2d6e74c6e782fa950adcb52292e5b8e7eff805772511e785a00761890693d108943ae8feadd9989d61928;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f9257d4a9d1613e14c5756bbb3a4bad1ddd18d3c24d079b81685af1e5ec1ed4ea65aa88ba550e99a3c23a862c51bafa8b6f0f8cfb590a0be1628726d89dc0f81c5c3a8cd8e7d15d5445f6eaf45a9acf0aea7550fb4214b253687794c297fe8984c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f95e2fc7b877e43c30d0b6b265b79bc4505fab84b6a4c058dd2f0c2a3e7cc3069ebe1bd92e44e9055584d79cf95b3a3c65c9a52720bcf24b0969fd032e64c004f93aad58823d8641ba2f2572337a228362d903ed89cd5afb4925050205973658799;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha01ca53b7945fdde18b6f55147a9896ec4d4b9e4ab82f020a6e78a443ae2a0920d25f7b40156f2fd4e8cc66b5aac7b6945c6b8e3efbba0ba9bd7a7dd807bda20fa19c7498b3c885f441b3585babd53c4d8ef4a74e56197bf6a2c104ae45b10ccd814;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha86e8eae79c831ef6e4444ce85b4af6cf93068e2da09e04cd6d2fcfb604bc3d5e00524e2685b8f593b64e365cc2a710ba6a6753067567372a7a50e56165c4c805de4e7a6963d2ef44e4b4df9b37dac9b26d4f1f582bc93e572656fab028b9dd8dc22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9de887910e893702d51cd748bbe77d7b43b4c76d70dbc6d041450070b0618994429a151cac5f1459eb809d3568d7e3d3a5e2f11076cd3c312bf07134b6257f8206addf90c80638041c41791a830f5efe7ebda74958791cf26bac96941a27c0abd96d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ce2c634de8907605ba0af3dbfff483ce04b56c3594b640c8e9f96e0b7bf1ffc8635e34b600a70c693fbaec71b23ee7df1a2e30389427cafff2ca6fca8d35974770b7c002f7e3417418f37b5e852e3934953e137bef8300d241618955dc705b690a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ffd445b866fe79b8958a73a8c671269afd5028da13a677eed21aa66a18a4441c39ad4f9decf150aa3b4f7b2e7821e9374bc77b611d3f58d8a1e5342255ec1208991e8990195d904a34fa0ce716c2a8bc6b231d42fb743e52f77b5c716527e668c2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dc019fad60a40455a81749d0361f39aca9848ced59db20420fb9d4205d40183c588f1cc3977c47b9c0cb061e25e01f003306e58a24c3d31f1313a85a2a7ec4f842d80740129f7f533fe76ecf2d9485d6779867bf8247a51c96ec5d62fac1239b6d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdababb7829d717623623dfcc6a037061f17c72dd19a6b319f4d73ff54cbd458b22e2e6ee666fb00c83211e0e39c36b83bb80123f3cba25648e6844fa57274c57f24f536a53de20bb7b901e359b234d2bf2bf9df99fd7771842d1e5cd6f23af81d06e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71bfd53694b01659c9871f428a5d5b6f26542c1ace87ae0c9b4a76d7b31c4d7531be0a5dff79dc6aedeb7a866ce606531b5ca4c9404e468338588ae7715730fa0704ca757798ecca9dd2d6db9e5ff55f1720a27453529dacdc38172d387d960e5d10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1df6256229c4db82f9d40a4e71e90c36c1dd7bef0c996ea7c9207dbf6481b7a0704857d9a9ec065090d70352cc2fe149403848c146afcef83a29a3f7a8ce291b08d353688cdd0ad5f2ccac912809bcf850acc63303c2b4f00a48998e2083c20cb034;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bc124de20a093b25f3e45f9a965191e3d734d0dfe40815b9a8aa9f23dc91bbd3e562d9b6c535c3387919fc78f1ae78b50207deb5ac33960b8cbd9bd54925db54d9096e1a300a9672f0338cc0d66491c91d37f40af502d8c255c48f9a54c939536a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd074683bae63e430c0842c0447c67c8aadfdb2b749156fd766701fbac209cfa33ee2578b46c16f09bb2490ea3ddc0351412573b457f08ea35c359b44dfeaf1d3579e656bcb7910327345c865d36f50229f468975c501fc2dcf4b837110a57ceed78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haea03a9385562e76b4c6e1549750a30f8339c5fce0da176c80c71cc4c7dbc9bc300a6fcccb67d7a95fa61c3e18408093a90c217ead630ccc358d41784e0b598561c95fa8a133fb57ac8d87e97a0a6e48ce6f2e4f2e0856bfb0e3f402eef4e2df3c36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a85f824499183776929fa29a1aa23dec206dd8d01c5289d92f23c2b4792d7f8c35706755132990300c5ee27567c6096169afaebc59cb2b862749e8a79488c94444aa3b6b10438a6b38011aa82f6f597e42dbc242b98dd38f7a9634c6809a1757096;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76e8f70dbe256d40470b22afbd8a33d4120c13e2f92c14286085ac4127cf5357d576c66073c54462e858a7ec1755109edfaca98d6c3c26096ff3115ee61018f10fc460bd1320e74b26cf2767669a05e057fd6309b012e5a7055927296cd2a71cc46e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h942cb29189833de1d8af6551eed289d8f75151a1711a15f85c7e40c30072f3902bf15960b84892dd170ab04c3b687cfc710ae15accd2396dbadc6d9729cb3329d6f883e5f803ee981e09fc2735e9b50487affada6ee73a098f164174e754624d4b7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d2dc35a4ec441d53549e94c0c921e29beec5f2aba886286331417d92a1640b5c9b464bb5dbb3d6a08576328e5ad91983c0cc5bb951c244daa9bf5d357e5d0dd60da5dde0bb095fa77b3ce692d90bd09758f483ba08cc160c13c6a24cb06a5a1d028;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7f940d55f1e14a22a55121073c8a86fdcba0800e5a0b2f97ed24e83c65aef12d6182b596d4fd82f57c4f8b5e91dbcf40300bf3a8139cef2aa2208c15e8923324890c93826d8165412b8f3f26b21dbba3455366c8c0d2b6d1d28e87cf9c397bbae2f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d90e733a729f278785b6313eae83261c28aa4d995f8d9fa178b85159804fa11bd970e947ead029c23e34ba8eb48ff5420eb8aa0f2018ff84cca298d3e452f97194a248dfacd0b21f4f298ba5c3f6ad18bb771e463be2b9a1065f0991a3176cb542;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5d06d10847015d9070433c86ed2f6e0e8cade5d7144e514dcf2aa7bd7d766fd2428668ada569fe08603549e2ea80074370c10da2974762d7d9b5fdc206739003e33fb41ee5ae1fc39556d5788b5f8e05ca9c5a1801eb69f6067e82604e93be2f544;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f91bbfa7a87e4c0b1bb0aa2702960c9c05a717e9e0a7ca74f02b627fed5abb01ff3ac972487242a3679a067829fdc07bf58ee40b2b1cc5feb372fbced1c05203fae6fc23aa177bea84e61cec71b362b0ee06cbbe6995ac9b5cfc09f0ae55fa2aa9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h747595c0acbbe9a5c24301f8abedc565f291671d3c646b76e9aaef73f102851c22ee94d45ebdd5a690674cea4929243723b370083a7bda7e84c7223a97a71b93d4b2defcd64807c3a93479f440925e80e2bf6f375aab97188ae5f39f050d2debd96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde8a045bd756d0a9e312a21f9b5e4ab0730a0d89911fc8fac5d612be2b9f7af7dca202d51fdee98cdeb95398590525a57496c7585314dbfa1e1c9ccd9a25e5a384a72daa4324bc6a44052008337e9d575a5ab64dcc9ede3629eececa9de8675d7569;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h779982b430b7e1512eb4f33c5d60a80ccfc8c19f758b7fd77aa67787f03a18ca6b164a32a3682cdeaa239a2e74d74533c7453a8e976119d1ee394b9c5f76b77e232b25add901415981dca2c31f1ca270dadba8de2e5ffbd3aacdefa3f7d2c38c8af6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d20e33dc2a1bcca77bcbfdf36bda362d205df7623f41695a6315f59116a3616c42f27d6b891d84fd1ab1b02a0cfc48856f5d86365ba417a0a2672a5d8fe529a7a3c1a50e26ff1edc8a5786d8903d166b021402b81590eae1b2a2da4818226bccd10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf9e6b93f1ef01eb2765f2d77b667a6218f58219be968322ababfbff533172fcb284beadc8d96d2278c80a4a3aae91292fdd1d8aad786054dda6a2ddc1055ee3c2eb9c447206147a95ba75cc1436fa5a5bedf378d0336f53a66b93f2f1658136c922;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98c0d57fdb707799ca3d7bc3e0af0d0870efc28803ac65422b0b1854a5acfea64b5fa2f5c27722573604437e4ed6e2e04155325d1383ef48fe33bc56e4b977f101fb6246a16ecff69d7a7db8f9007db86f8500f6a6267722238b07c098409d47a92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98a5462aebb6213be15b2cf18c6d6e802dfe28e23311f6c6705835a1e49125f76a0a3c0d2571f82c2df561d79d81c6333ba73a0a77c5659efc239e31da46ae1fbbcba974d38d7e9a7d80bc9f886d2991aff2be42bce4f9d246d6d270c0c2a66b473c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd64ee47df01459e5e6975bcde78f46f2f3fe8ff0e69362aff438c1b7cc932de2d81838aaeae65645ace6c826bfb06e967df3c005a103173d315468bfdf46324e123963ba2b25ba6c939cc110d51fe3afd57f646930035fe93d214fa9690b1061c5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h536f8f4e337f097b56ca508d5d727859296c5893f323e93cbfd25424c6f69da69a58a0c282a126b3fa85a65c211de89ae80ac5018e2ef026ce9712006f50f4aa48737eff5749805d2dbd00e7f476443854cabeee270b322742a2a1160c549a5478f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98823a2ddf3c16bd4eb97a59edbcc75b7511fb8734b62038b509384437c00c4f1394160dae1071c56abe75bfa31be5d7d066c0c73a1d4de13e672a581c27afe5e16c3a824706248341ee247d01b5d0f6b605da14f1346b680cfece0aedfa61f7a542;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89f9e80d00a49320295da9edb057dd5d96ee7f79c6c4af6b9a4f34a9584906aa668d3d383443845582a504f1fd9f6874878e4e90aa8df2b457c42dc631e1d25459468d0bccde0c1cd760ae89da9f4a40e91c7e3600f785dd6d3e08876873d3bf97b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf1b784d359a9f7c9e64827185944c9726fae360f7e078fbcea29a42abb8753708d301b2f072d3e635385bc440a70b32d8c2dacad53deed5296064229fb761605bed916d558013bff788eafddf561912ea7042a9dcbe51b9d5e82499e974d8b7423;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8abbcefa2457bd07c33525e1e0fc532488a3b762b0ceba24580a6736af9bc0d4c27c510e8b6e41d44180aa7cb5adf335108f3e0a65c18855b3ab33f64860a76463306ea154b5609aa5b0bd95314c9da138b0f9eb25e9b1af5f9f8fdb31f85c8e8708;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h643863b82e53addf5b91a6d213ddaf0257e1871cd90763e9db0463321bb9c968751311ba64d00711408f7d0219cd39c8d5773b4ee866a7fcda1ac9172be61da747573ed4ff772a45a7f5d8da12d1e0e3436d59d282d533ad675c406aeee6fc9a6965;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h451cb7838126615962d6dd8013a654ab8c88e6e30d9b59b8bfa80774bfdaa4c6975e8f5b5149c861e27b4377d0d81cffeccc007d9015cd74ba91d2c8f8bee1345b5da2e8a19aa4e79c3a54d3cf4583ce2f835a2140408ffba99eccf4b20e8bc025a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a7cb54c1a4694f7f5a9b041fb33007034d061f57f78e68a0e025d142fd629c4e0610f47dae521df01965ffe4c3380ec768d9dfc24d0d00e34b8d610fd4535fd9f190fd80ee05068fcd9f7f31afebe02307d5dfcf5a91cd251579c242bcf40830441;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2689aa1fceb9edf01cb8bf8a7cef7595b527670d82293631aafe0cd2043bf505724111aeb2b018eb177985f6ecb5dde0a9aec0437449f75744705c468a8e5fa7485f6b8f87e0d7af2dc151edb9d8480845fe89673643431f48575453a633ed9cf57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35f0d92453869a290ceb2b2022b6bf1f21be7c4346d5710d6f3f42e23d06b1198233a73e3bced14d7a6142bb422d0fb8a60091c03035bdb0295abc83f05c736ff3c235c044ef8e06fa71488c7e57e0ef3466be9163775ad23916b2845ab00250dc6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52af75fc1fd7748b2b7d1b78b686502fbdc9974fa4d2973183a647e879cc73fa66dd667145d8e09e89fd9ca918f4c99695af4cedfd3061a11057f19f726b8ec1962a0ceab0aa39866e6ec56f9684b39dba797a8de52fb2bca91d0606a8b35aee314a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1b8b1b5629121b0940c96789f4265cabab7a29bcef6d8315237d4c2bccde5ec9ec6cadc31aa7d7307c6966c3787d216f94e5c886141e65824083eec6227d5a6674b762f62928f8487bcffa5b1043b3837e77ab38dc7f6eb9527200a3cd4e2122865;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5a4632ecc213ac9ac8da34b5f12e0f4ffa5a1e6ab84ccac2d25b26b78faaf3f66d8b5df30ab73360143bb7be2c6894bf57dc7b924d601d6be34819d0d83b69862cb1ca4be0ad7f71f4a7cbdae7b680b2e041a8fd159a8d62de0c8b564e9d667c30e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b4f6ee3cdf6a2e4d6fa0d6b2b999ce6c29244074a28b1866811b58c625513fd49ec501f7d26651fcae970fe849c51109c3e6fcd9b41588efb04cdaad4a8fa77d7347fa4a842ce1e3a40957e52ac628ec1327f1d37229e2538d621e553a1c667567f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d0366eabe366875ee959ed064ff59a74710bc09c2a3662fd8dc79c0ad86401c37deee68612e6f4f8ad251572676365c6fe73a03746fb73c3aed41cfe37c6dbc9934503a48b27ad5c7968419ff3eec490668c9d17f3ea452a1a065419e2f68decfc4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fbee9258490aab246617551aa9f236e77012ec59fea893d4a54e2e6d0141a7ecd4c9111ef12f8b274e9bf71bd24ff5341c5cdbfd3cb78f72b5ca56fb5d4fcc4e641eefac51e0eaa6b66325c8fa2b3c685ce2c235dfd16edfb4d8436061af741ac02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h300bed7538ec141291b7642b5f0e7fc29d96ab381b31dedb609dff6ae87fc3daf878ee6c9434716d74fedad7c2640b7f3848f37c18ff599e580dfbde452a3a5f5b029f6929dcd0239bf220da59e02ea79ffb6acd9c1e13a5a51a86ba5f07c270919d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacf5b56bef06b228b056c8afce5a599bcb9a22fd47f9af56b85154d0db640aab5561448a33224e005ac91717b623dd867546e966f3e4249cc98481ab7bd2cb6ab905753237afe5aa3c02df95c0b3cd17bca9c8fe88f683f79339e2c915b3b8dbcf82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfee7656d2c7b6a65b11a50f8ef816729596ec0a473e2ce1f020e6dec0daf21fe050176c48621f9e80feec7ac8392b3633ed6aae7dbb02ae45169ac97dccaa0a504f1aae7e5d9b64fbd7645f314d7035307d273524551c3bff8bfe3593fa5a3d5d3e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5de92c016d358f4dacf25f877e578e3885b031b1eb0a1484d10fb27870290737cb3323a954566a1df4943faee5ea188a5a02c11b9664d04b6da3cb2864f4b1e5c325ff323dabc7a8b2de748d8fc721fd65abafe3349068563687b2aca53191718df5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9759ffbd5876e025a0b06b26bd635184a9ab2a69b3ee896c85b22f4fbadfabad0f2434172d669f2f55b9f47042291eb58420bfa09679f6269d17c7aa44eb60ac32bec815efc8b9aaa9cdd3bbb8c2d4fa54b6bce4b6f5f61830075a62d41ffa0a8348;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb01d4b5db112b8d58c6734796dc4169d2d56577d8288c141fd62a148bd19f39f093a569c98df3fd2909f8ed4ab30de2b017c1623b1ba16a968a1f9eafa812f6632c444706c0a82ba138c8dcb084b8f4297d92bd70ec52dbd3945f1d720f33a0cb9d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cbfd5c6855848f17b76ff807e510e6a5bfe675b8d9b2d0308285c78d69f0f87ca3366a090a0b466d792fe83684cb333ecbf86da6c3ca8c3692fe03638224ac2ffdc0461f85a78a2bf6f543d302f2cc2cf487871b81962039b0d44a2902cec116060;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3868035399ae73cfa8cc3b037401380dee5efd2236fa3ec5f47f4ab992741686a500ce7e7e4c972636623ac2bbb790eaba07dbdff36dbd2c8ba9d1c3bef4958c851188d1cf52597c071576eb1dcdcf182386aff6d8968d8ac070de057c9178b23dd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53ec258757438616122a0004c1dfdbc59ec2d8b889824fcb30b23cf9359d26a7e59266520030325306075ee218972f5ebe98e452aa1f6b72c383a9b80bbb783df68496c037cc6194648c28ab07bd723885986fedeba8b233be1d2a08222430bdf6c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfef229584832402fde41cbaca86a2f1e70f09855eb9823f1a9e01875e089e40f089196497f1cac3d015bd7c0d919156084cc968e83a76df695ba7b9ab4d817a290ef2c5e7776196552f72a9ddb0b8ceefdfb549a16ec0b120994ec1b67c40fecbbf2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7cf4ef5c2526c4dbb5f54728688f07baa778c53d28a82adb5622a8af28fabc108ff834049565c0b8c4ea33999c57e0a2157bd439f4a3a2dbe293bba6f686b61373ea2a7afbeefae5dff83b039590c3a84f8bf2cb19323ee44d517a40fa9483452be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5493e645769605023ff27dd80add613d578eb1fa2e5ce05f48b01dfc41d28ab5ad7f75d85b64af1c25d6bd83d56dc90073594445ce032fe738e6543c91002e3284a21b25ca42a46c3ca85432658f8f905a341e8a69bd74913d494309027db679228a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe8dc4790cfdfc81eda06dca60e540e67589296afc9307103a92accef8c9f2028fe9e8e0d1e63fc946beacba03a8a817523fbc9bc0744b157488be0ee9e64adc370619e0ccd89abdbef15956d482ba14401cc988c5968d116816c741d5166dc443b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc93dc49820512ad862cab14449a8eb2b5fbec50d6c84905006835971a98aec196a8c637cc23038747695e7f54910020b09b4f92cc0ba256ab0f3c47e07458a4f6b65738d0ac6e2345424a4eaa2767f257c1b39aea3e952fb16e3de1dd72a66411b8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h485edc99dcdae621ba3c1d5ff1c82f21d8f581a94c722f7b1f97a82e34ab25a9b3bd991aa0e1d6c0df97bc872665c353cac61ff7761ab9969a10470189d6133eddd68e4478f19e988e9424b136459e3f110684ffb88f681e1fc112eaeff6ed0d5129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84fbf00707cf87a06805cca640dd6954edc58d9005144862e82b057da757b9bb9432afa5f9cd362b76853415b4760257ebf51dcbb4fe0384b098baef06c9f35f8cbcbe42a63a285509f43836fc3ced1b5cc2568aa31482a924f9531f4d357a3fa389;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ec7052fbbd21909035282938d7fd68c88c08f585ebc2bfe81f4246418b264e71928000e48a5ee7ae251dc8c7b5f5d5c6340609d90c037e0b814c127ba2d01b58d6d820a7283fa4f0ddc1b405d8d9a32270420370f467e4f673f01beac56dcef9b4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f3ee90bc4a68418f674b347e7ae32f230e9890e5ca87ed16c31d637393965152fd4b9f1e5575e35c339b4580e514a6398d4db683ae7e5137d3ca5db697f1fd21c249720cbb61d8d74a433309161355a22cba8022cb17747b441635bbbb253cbbb48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c9317e346768bf6f37c8cd56825ead63afb8817f41e86b5998bb8103290e549ae12a5792fc3dc2ddc781c865c6c1b74897ada8f19cebc1a7866ee5111be9c8b094fd31954577534db1439ed3ecdfc167e5bdd8bca5b1a821afad09c3007c1eb4f80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6817a51e66368cd31caf2f73370244d444a379c19d2c348da72f6eaa817038b67214daffa559845d98aa11c8912f12a4713fd63a6fe660b7e6597c938da6e1ad654d1a9f56e00eda14f6390afed66644ad87ed1575838a2aab6668ddd7914b19aca4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4dcda2c82c64b468e8cd65ff128ec473cff33b2a9d308ef0b8ca640943b48ce40127de12b295ad3f9985435c79ef7cea4db6db2377fca910b73a6f15c164ac743e98ebca6beb2805bfd90f67bde9d5361672132d7696436378281c242a5c741d046b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h676aee0ba109e2715ccb36bf2739030ef7d2e7118226d10764a9ac2ec71e3bdcccb91ad680826af80ab66af4887cc2392865c51279a14736e72542400af2d313002755e44d312cf7c1d305d65e899801da6259b038854b806b150441205695b71b15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cc0b13119fc03ec0ee763bfd5ad0902621d89b3f1eb62cebd0f8ac68c91f45fd2c9249e3778a10a6f5f22736eb3d32c9b9e7721e8315f3c474eb89ca5b4fac7018d3ce45a23c05fec3a8a544392fb087fb3aa8d7a778f62dfe04b13d26ba2bbc918;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97ae8b3e7a2560e252ac9bde821169958044b3811e3fe8af741fc6e4ee46309bcaf732b4aaf35d914664a850cf7d9efe42a26c6cbc639e52c3ca75a301ff891f94fa4433a4a7d111e544a829222f454b354b60c7dc5daa1266ced71c02779cfa8212;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61e42a4b452d41da023594f34293120619d728ba41d8c0caa0533e12a4ae7130a412f8a1e5c84b677b96ecd02d4ad24e573c693171adfd8ba8c488691ce40e1a28b364655f557c1070fbb311e979a698124d793ddaae8c76a64d3dfeff00aae340ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h191a9b2720306078f98f511c04540d573bc584d26377d26cd661357489951f0ac213ad9e99251da9f0f073697c9d600a231b03f206127fbab695c8425e2fb6873684d614766e056d1268061f2d971b521bbad29d0d4c59ae8b3b0ad924d91fa1c591;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h495137473a07d18dfe2e0200d6673148337f16e4d8626a7d103eb91b84a14c4b2d780129169ba0eff7d2961499610efb486bd8bc568e621bb2b905f3eb35473cf92224943271a16a306f4c527c6066d6bf2aa704025cb168bf58d22e08a750e43e49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fc3600505cf3dde2fecc986ab0b6c43990d935cb3fef140714ab1f84fa5775114826c1b9fe369f11039bdc56f26c5d2baffdb2029a35c2472a432ab5ac51e28ad6318c76b87a4ff0cd99de05a4849c9759a38f09d86ef5a659cbd64426f2f2fdd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h110b0b8e968c3666d751e3a50b687c3e6654e2565a51dc3aaaf0154d092b42708555e1d3b1e4d27c0294c2e7182fe194534536a2a6d6fd6b01d8cc971dc7f19127cfb0091dab99c7c29721d640b1e3b85e657da565162a6c6df699c0d8470162c56f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcd577c0b5d46ee19fe07af95e7d13083a5689b0f0ba6d881e6e4a207e5c34bc7c47eeee67baf4eb5db0bd56b0f6ab010a30d078408cc046e0d54fe38a378fb12e835cad3fa0b3c4c8f2604d8a7cb6642c8b3e5b7bcc35b589fa16a984180feba6bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90fb3e8e1f4f282f2a43a8db338dbceb16cdd8adcc45080d8899d0c4c794365bfb431ae21f1223df21b2815c96ca94931dc1bf9b7c37a82fbb2c1904a5d7591632051019149ee74816e6fc8c4a625cdc048ea24686fd0b794a65a3ed1bf202db5eee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h675b23c5601e7dd2867012e5bbc9e5593b94cf1b2a1537e14a43fe43af910706d0af9be30c887314047a8d472230d42ca0d19819e3cb002cfabba18ac4a69b549773c6d21988a86810fc5e45e14a044d6a171529813457fbc947ed89160551af4fa3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bb7e4180a6345e44ddd60cf234d0f9099cc49543a3de7ce6801968082cfc0fd207b953bff261d5ad14eb89b591f9b9f5eebb2ae476d26a4757f10369d9c9cfcd442d1dca15e24a2c329170899b35bf94cf664bdfa8e2ce4ff5f4e200ab58ee390d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb75082a9efa9f0d64b14ecfac6a43e7ce99bba2ba5063050a8352931e1f1d982aec325701024ac9932568320645539048cf4a4877cd9b22da64e222b7144e906fa5a4b7cefc832a3284a79072c6ba8fd55e34cb5e70742a53019e9e944bfac7e489;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h436b0120d50d2e5f58b48447f8af55872c5d81dc19f2d8c47f6382d339d813a24830873ffa4d812d631dd3809965357e330eca9dd9dee3ff1f677185e974bf8bfdc4a4611bdce00356d06d59b82b5148da06dc7e7febcfde338c23a913ddd1bacff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6af3c1623d26ce25b4d11952c9c4ade6005c6112280094509aa702d559c4802c38a001ee50422ff4e2adfca8f900a7f2246def24576a5624658caad50ab3c737b6bd0b3761245a382cfdfbd794ec1023ec3a1c04cddf98eb77b6a0eecad32548b2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fa9e672ca32b3062bc32b8ef0e9cb23747d5648a58531f09f14cd81e4b243a9365996fa2fa3a6ee86c1cf82a5fe3dcffbfd4a01eeaca387616d335530a1b550a29b1f5f2cb59e812be8a8a58db89c4ddc436d0d83e05fe0dc9f4303cdebc7760582;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fec4cae7d76d7a27c6a082abbd7e2eff48e33baa9c8f9d8a53d097d1be32e740db6e28d513f42c13f49eac5d3fbf46950c0c851223445dbd5dd318609596805c00ef9a3c2aa26e49b0de6112c1b464d61c2a5d1d6a599f71c40fc71efef9f7b2783;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d2aaaa81bfa520aef95e03cecc3217d068d84411ab4f4f9db7126b074790bc9a3fe5cb6613af184409072642b8d7ac36fed77cb3faaf7104928a54d95176670eb022b046b4e795890295358b3b0145c3ed4208f6ae68f1c126b45546dc6318e842;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95dc343869adbbddfdb310f372e97b84cd9a2ddc8d2cf0b6d1becac78f84f3d2d1d8bf7549f03e7769feb97188f817018f1ac185fbec3e04b25f8674e3c12a1905500ebf337092adc0b55945bff16ed04d124754d05d52d4f45af1d786b438f34795;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3758883026d2eed6ce5637b8b854f763be0efedfafa0c1dba991e494dc44b43d58e50a6a20c4fed0d080f31a3b8d940471c49bbe206d8c34ffa3d19aab2ec873cb33af0cca93733f021082e4948062a45a42dcd101310cf8b7005a09f3295696775b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcee37463fed16909fa505379ecea2b1b92e850e6686db8c712509087c41f130c68bc48f2f81cd82f3b65c53bfa67a04e7c7d4fe711d0172ea6f50bf3e0f7194ecd852b238270ebceb5d52a72b481cd755ba15226348dcd92a27959bad26aefed0fde;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39ef5784bd1f887e4b88a505e32d7f0c0422a55aca0e36d5646e21a997b345803fc73ec6ecbb974fbd08df967afa6b0ee39e15ff8d5a236e3f1026f3a4719c7c3d18b38e5c76296fa683d8a518c478af4d45f22a9f1bc7a99bfeb0babeb3b567bb3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6b17adb6efd4183842395b7881c66dab71f6ff71f4b86e830e1debf10b39590ef046d6b5a3260a89ce8b56afcfc296d1f30aec8d271a94d1e3c2e782d11d8c9c96a3b48b9b51e317f511848f4bf0432a4194bec317f1c72cf172b5a90b6ff8eb784;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe848c5b00a9f533266cf3fd7bdaea5c927df7aee39f27d265c3e2100841483d316ac421cb103e01e7a99e52bf34214eefed16c688e983b9031fbba21a43a1754ec5d92928c35ef79922fdd020b3a40435346b2af3946f2fe80c0df209e222586821;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3e4414bd9db869de384905501b9099d499ba13c0d118d48c6e579ca3018b0d39779e1b4c018d3ec2c55f1061abe7bb278070ac49f6ce6b8a8ce50b8b11da0023d3484ee48c3ccff752a420f0452cb03c3be1cbb90fdbf70e02687dc8c60bfeaf253;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35a5d5275afc979ea40ff5b58c3dabc89db5e6a477784aac327d4efaf6c49a89f3f31f8c8d74f1c7435333f6099553b7f9e80556ce9e9b33ab1ad98b28159df9956d5126f071983a8393522f62a2e9814d17bda0150ab53a72502546f8b97d80955b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c906da40241b5a3872865bf7513b871bd3bc439559407cf3d5f0aac19402860391fd7bcd007ffe7fed1abaedf5b6010e2849085612451ad288168b372f7bc4af891cd78dff98e77c5f3d3083bc85d27234417094fe2daabe114b0bd1d921eb14ad5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f8021ddfa3c2f3b519d795ed074db9919d014b29d256d11963bf170bb8fe54e1587ea49e8125afe6e9837b375b367203104998e5c47675ba4899a8d1a75ee9770fc367d916296ef2fa9104f207c92f29416a2acb5bd4a48db8d8103a060c4df8846;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h298e760b5e66de0d16106db28741f919e0a7ab6bcc580ba8e213c447c34b833f43e899e37a4dd4fba0feadfaf068583f10d22ac0b554279c39d15787daca2f3fa34c00fb04ee26c9307d6ecc1f410cb96ae3450066c73cb00574570828544c491e28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1da824c9144e99aa4e172891dd61001a20432408dbee0218ae2a3765cc601c200a33709cb504fe07bfcf4be20e0fa222ce85d9264215d000b0499ef4f83ece6455896887850893f366b5ce821900e9cf12a98df59a3521bf19d60a53a10b344b9ea0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26fea7eb8f8cdf4d991e2e6ac6f3911ce760249c93b4c152f2b645a187b86154a13cf179340351ff677d8e5e1d08b76a5434aab3f3994726a45c60031cb707a45f925afa0eafc47c5da22bc8581c265c4e437732418db642562e2b16548bba57970e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h886fd3e62bdf9e89185180f1a65c556c448cf40b2f7e441cf15b42fc29fd88be1c28021bb10a3d3f5e6c2f6377deef84338fd866876c2534967a4b23e1d18d1002e22fb1831b61e076fa04b68be91acc59616bad1f552caa11b58f5a08049c3e2dc3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69d98305cb3cd82191e7f3cbaf37a0defa0cd95e6a556fb71b38688eb50db54690c1e9770de0c8fa766b6e0aeef282044940942f90a5edc67b55ee3731307784bce4aff96b85eccaebaa75131b48dafe8f8e3e9d0fcaea4aa053d22e8481aca3bfb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51f0a680d8b229a785bc2642c7eab4b9d8221d1df4beb0f4a997609ebe7a939f9ea5503fa86265dff47f89ee7baff033f8ed2ad0b12e65be57e364fd4767615b00e0602c378a1a115457479c5ef5a7dc27a54e8cce379f46f18027e6ab7e3a8266e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88cf6b5f435bac89bf460748ef7928e312425717bf40d9ade252ee9d2fb7e7a966eca8fc5eefcbeb22afcc8b9729234d56c29ebdf75fbfcdc330b61720a82d90136de5c24b027dd5518480a5a9b9f7d1e60171f7fd84117748a6607f99e2f1760a6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2e6f692c8c25bfed1f7594c95f265f8e94b592b517f60f7866917fcf7f7cbfc01c36fc8e78841ed605629276481c6e8d3504def23f3f6124162ac6db5679e4cefe4488eed038aae8331104a7e3fd3ff119e7e03a61ec2ab5469f55e7c5f23be2688;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52c9dff146e5f1ebb451e6a9f34a5364444bf6a89c19a30c8c129a5a927bd65c69fe3bdfa4fb1546025105129444688ca6b20013aec3c4259f0bc228afd631d184f3fe5d0bfa337f74118262929a54ee6a9f9ffabbadb30680f58b050835bea93ae8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f8bf4fd0138168542cf79a627fa93abf2841c357fc810c077f256a7915cb53dc33d35ebe6446f765886e8acd6d3221dc4fa509f63b2a7c55d397a7986aefc32d52784a81b65c71cd156867993ae88f03e2f90001fe8c471acb6e14b100ea7b6092e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bc498a86bf28c9f0d3d8dd0b69367e480c5ee540e23c9528096219c539ed205cbab0669368a8a83bd42750361aeb0e5ac8725218a1a1027806a473ab0ee1707ab7fae22866f96334d51e8a4e97af5f326340ad8194ba802ce49f9585db34dbcd45a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0f5972a017c5b554a59beaabf0c2a3b6988d2efee2f2961c6301e9cf0fd2f55299710aeaa45e213275477b39bd252e74d91e721db95d19c4a7b8f057e19c2a84eda61889b0e1351027c63694e62b2ae23c1bfbbb489903a0163438fcb607db2744c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61e97d5871764c4748f3e992c751c7e82c57847be26bca0c8da03d108f9b5e7dcd6ad383a44eb1bdaa4abd345be2f6f2b3d6b656c120003aafb8a9da65b40fd5dcb4ce22689011226aef23740cebb76dd1ed83d3f2a4b3ae8d67abee28c2e9db9334;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8b7987c879e254aadcf358efa2daaaa105a25b0cf2d70175574eab764483acf3a726c6edda3a014165f9036e22758b62c9cb74f77683a2af0ceaccc4e7055a769349798ed3a1eabc122f1ed3a82b50bc43a50bfc287dda5b089867e749f77e3bc81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8700e27de07b5e12e43a2577adbdd62bb61051b92f6b8ea3c6c9af03120d0e86122a9e2fc3f073ff823bf28e7e52064f72121f6cc49490da5d05bd0dd5bbbdd419627c901f65a00e34799a2b4d1746d72a2be170ab770e89dfec9747b3d9a19da539;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd309ef98aedb1f490ef5824e9267d2fe8c3ad9c673019aed746d57ac10632503d193e94d784a5d312d734474c1712cf4b5204965c114ac37be3c687a9d000f1f2bde19db95795755e2732d0662566d8b16cdcdeb23e81061192220a12d4ab5b19908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57ba51be86b038d741fb89ad10d4e914831aa4871334419c4f10848ac97a7564b5b36998c28a50d7a334163084e443037dbfe1e7a554c6a57f5b6ccc40865b81e5554c5788ab151c47783376a88bec540170ef20b3c1c100fd6540560677af390c41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fd4208ad19f2aae37265b23c8062c7a915df5491c22b470896021f9cf8da27905d1a074603f24a608d2701d48d4854a627c7fe65d36fc981d7aef5df23a571f35eec97ddb70a5d9ec4a5e1d31df3b713204b032d9c4731c0d0442049edd6815ce98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h348fe253882a1405b9cd87a59d8161f8acf6f16e055bd36b188e476fecc7bed5eecf66bb05fda3346993abc19d44178c5ed9252572d53499847eabddce8ddb5119f0e4e6f022dd44acf97d2d7433e2cd1183b4e7fd8afeea4554d38517943bd10dd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0301332fec5ad8fb2f9db72fbb7e35e4a7a7ba2b98c7aff2d37e33460a3ae05a7288ffb6351ba35b85b20602fc0425dbc303648d8d26bf1c7eb750539bf661fd338cc01f79db1c9306121afcb2e57d3d57427755685f67f5c1ff54460e3d14088fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ec784759348bfadf1d09b93ddc5489e11a158ddca6e2bc2e00d7a98e19cc8db37d9f5c552984cc8ce5274e1c2a9d9a064c66f04dbb08a46ff8f00da4947253c35f0cb32e39fd328f384fff0b75940f1ed3c1e15529e5d54fe185265b064b7d97179;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heba8480e0dce18c2d2804fd69c6b482349354bc3b0d71b1b518f1cf93c4f6a6e349915701c8ede4345a66488e7e3e36f60ed6aee9e9c7a62f8330ab02bdac68469d784ba2d4fa08fe3835655f2af63184cef7ffe3bd6b4ae0f9a418628c03928404;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa06d8f92b0d463340d15abedd4df46ec36852e267d109b5df21a11b7d67ba2cd1440d2f78b5fd3f288908c5db00702fc5bf956922285ff6d340535fecdf2c97215e34b1f198b5a4e7c06dd7f60b7d84a5f6669410a5261f57665c44b07723618982;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a8ef60dc1c834d0cc3fc347aff0e9505a05a8c513d7b17b696662560c278620236851bf31c8731aba1fa89cea11a6d367f17c3dc8dac88e63375f6206cd83a403d1df095d37985945dbe8d0aa12927cd631862b36b3525a14d498fbe674f365ca1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fddba9839940dda089e2472349b1aa081cd670ed7d50320723be39059fd3571701daf2375a7011e7d9af78355d69a58dd117f980ca0d1d92d927584bcd8357ed9803a08cc331fc389693b482bd0441e04b340bf3dfcfab9b8341611de28d18cd299;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73a28510d6f70e76d2bb6ade143d833f66f44d4b815f8ab3ddce4221aba1cb64d9ede4074236ee591f13f037fcb26866c7fe8c1cbb0219a5b9e597e34d894531ef8031a992fa5d9052e57f7d359536171a031b0b6714c7c4a98a456a8dc6a63cddc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc01c45dee7a63a4d3a5b4c145cbd4043c7740259a2b7d72c358aec9e6957be9e63eddf7edfc62be5b33cf7a513593530801d3695d2998100a986fa56ec561209d33d21ffba4e5c869ed40fae2702f3799f73b3501b4a7bac6ce1706c74ef82698a2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddff380baeb400efbb959bc7c26269d6cd7efc82cfee39e85b19ceeb7e929db207996361e8612cca99125e3d4b7747f8f3f91f4d80318a7c3539f6c2c338f33cdbc2e0c6825677ec92660faffa31d6e32ae02677982c160c5d2e69918d21d0e3063e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f1700fd9c78275e671d4be6f22eb30bc21e10ff72b4214f2794718dc41d23aa55a65f1b1504a364f3a4b3f24bc1d11c52096f76e29fbc11de8ad8f0e1bf60a842c9d095aaa9c093baf7c5a1af2fd78443ae1a63825bfe33cff2d66e70d620d37cfc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f301924d7859264bfaef7916c7e574554b20fcdf222e8445419b958c5df45e6dee915f728432e2fe4223824d5b72cf078d00e7d41e1097293d16af9528091cefc4dfd4ac72786d8ce33925a688a4d643002a2b85b5a0182075b08d99b9a8741696a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed4844538ce1152f6f401bcc488144ca9be47835d89e3ae196a12b2117eb08d286f217df27ea051466ca77df9a27c05fb37c4d1e079475e992df65d34a9a425a52ac4d0d0b3f0d57c12228010bc2779f9feb790775e4cbb2b554adc0dda8de0262b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283e48151b355d1e7ed0522775f33e4654336217e5d3b2ce57e05ce017aa0e8d19088bad8a98ed1b9eb310c0118f7f5dba9a83112f09445676f9f1f796be36e27bd4cc518a0ffb1ffc1f054610f1c4cdec29e3844f51cd0c17b7110bc6e9b9d2606;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fd0c2b70924107ca1980670498c3d31da23bec914e3be29136893dd7de94d5523f769cdf00d926f0b3f8f819c3211ed659b38a4354fb6520806f10eba92d4060a8433ce743e6a733a08aa36f9889a916e3e846662819ebabfc4a990aaba78dca6b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf95c41063a851d7b48c18b48c5d33c986251af9340a5e1e0dbd6c0d08f3688791ab6e0fb6f56b9af7d576f4a69d02e4884399243fa69f9f2094cb01ecd3f254c68b3d74d76d18cdf15d9b2c21864fa45a27695ba2e2fcbde737f39a33cd90d5f6c4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59f3a19df1b18d3bf325e5d77336783269d8169df5b06da2b145eed3832e34fb9571a0b27626486f1c9ea2104b09e82bd3af450db12eaab49d75f4ee05d145712a30bb0a9b2709e528466e310537c2b5ca46761c02df9d2a0478472833ac1f29c505;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc881f9ad8dbcf10603b809fc7a3fa893724ef02f1229ba55986bf52d0723f3db93814b3beafeab178f5184a0ee95663c02f5dcf031821482ea844dfbb809e574df8ee4dca249cae3ae253a5f990e191e746ef6e2bfc9ef31f8999bab0106390cc3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hadaae21391aaa344b53265a1265c97444b9c96d6bca5374ac62a1f711ad8eb99ee9a8af3dfdb4f478c049f43bebda57bffffadca0ed775b38679e8417ccfd10ab64d4d7e3289a0ba56e9309c02a0000032d4124f09e5943e3d624395dbdd8d877ace;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74494fd9c7304a19c723b83f29b5948bf590bec89d22611f80ad1777413b507c83ba14fc84cb6bfc021e1fcf24288d01e8d240178f5200b3e8cef57713d1e672c435a41b7b2ed453466a87ae8617001f2f7bdd6b03025c4eae65f517bfd3c337df87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aeb5de76f20408bc649efd63736771063309ccf0f6c9249177fba62c2880e5c81efc268786ba70f052a4fdc19893df20c2e3d18bc76b8e32b6caf8546d88785cf540bc100438d7198215fa8d4dd228904599ec03f40df03c97f880d4e082369518;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h507e616ac3a8d830f0ea4964609107cb35fb7b42d17b6ceaf5139947b87a99833c62dd2b32e47dbb4e511fcb17ddd76841d139783ec6130b16b1ae09dc594c9759d745861042f5c4fe9f3f1b525ab96def9663030f75421ab44be1c570ab296ca7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda7f209f7cea54eabeee0510f6ae7e4979b5a68aad5e305dfb330da1f66bfa502379908f6fe564228b792cdf0cc6de8f54246ebaf07d6cedec5802faf61436e9cdeb3c2e890ccc2249bb0610f542c360b144a37ab490537c75715d3421e26766b4e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84412e1fe368d39ee4a3e725899424ad93341f71e38bf3d7f0ce064efa43f25221019d90564b109220f8464659d39cde34dfb6c940bfd1c7a2a7a445e12ea5f6079e618f24b8750eac5b52ba0516987df0ce7f11ba3a2874e8375c8f8d23bb7fdb49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc17482a7cae1c01ee3dfacbe117fee690dddd87906f0de7df657a34d3e97dd5be72b67cd4904dfd792ffc2d12c681ff29ec8431c8da1fa357bb910acc0b79087a8f7125138590fc990e4e0e003680c07f4d7d18547c0d6f0bf06cf774ca64374bb07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h575f7fc124a735aabeddc1cd155dd508115aaa13470e7e55980e053c05fe846d07ad4969c952aec06c7bf008a14b6c62bf26f5576c5fec038eb061fd7bbf665f0e5f05a25417fdac203d84aea0c17b942237c69e129251e7055b4454be04aaf3b47e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94de47cdeccd3abcfe43abb8e6bb371c7a3719a76a8f6d7ada8f27bfc854beebbdad774a9d54379c6826a0ab743c6122dbb2a1b5b34f73900cbd83a4350df2fba44f80da0070a686bc22e7a584a1ac56a3dbb3ae7768e270bb2814c52663c5a75744;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96c593588fa39b2e695f1ec1bb5c0eadb56a982ab7627c0eb83ce19b1803f755ba440996ea9ee3bf46bebb39c986088f90a07aeb64e2f6238859109976e0637d6cf431a666b30432c3f1b2727f70ded3dd4d0202112131250a5faa24c5beccc45c1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h461595fe4aa5e7a34f771d13f6a1a3d150078a1de41c610eb338abee0d7e18874a85af2d35f51edfa53d44aab1df7edfd24eaa0ac4c7abad6374862acf8095c5cda37969bbf4a59090078d29e2ea4ef51cf94e0f74356bb5750392bb9558b43b6083;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde8a57b7a209905adc4bed9d8721a716392cb090fd7ecdcea9e2f5f51aa68e11a84f93161e36b1812d999c51c3d2048ae9af55d5fbc80be79a1c5b686a3dd2e0ecd9771f476061ce98ade9d9d0c5406fc6d07521e206a36763892bf860d2639e3ecd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habd60c1d41d4e8258dcbfb17d35f2a3f00fec268eb422f3c50648b756f5358fc94122cffaa72f70c9efa015885e44ed4aef8d2db57e0d828d0192701a461c4dbf66773b95a7eb24a7188b74da50bd3f8639e04a246a33059794d3078c3d41b76bd1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57379ecb76ff52d86ec3dacc8b6b56365d6624a2bd9515c2588cf476aaa5397e13b9fe2ac26c7404fd16ce9a55d5320b1fc9d54db4278892551ffc83d0ded09e9593224e10c0d229c5f4afb8293ca67e719d4864c5a59dcb42ffff0a4acd376c2534;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b19ad1db37517185a6ee0a10ebc72a9dacdf4c7fc27e42184af2afb12126529e59f12e294545b7ccf94f6bff645a3e9dba636e2c7e8d533ff4cf266248d8c8d01cf9e06391d244d09482f3c2af2d62e36d27965efbacfa1f36de57b3cbf22e744b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64d66375fc9d0c1668098e8fa4e3ceec2932b8917e8d9d3747c5a222f4e85a2270dcb2046606a92ce184fa39a78ef8bd86fa87ce144b9917cc458b81248947528b928942a41d9df4832b6642f571cda63da6512822fe0bdf683ee70d04e1df5e332e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fd1ea9cfc07e9e8b762044c4215d8d3d1dff0924471912bc13e0c195a7fc6ccc4d24e7e2f616d614c3a9fcb7c191e5fcecd528bb2aa45f92864d05832cd32c4c986644adc2251571c3f2ec7c8fddb0062285ddb2f8f6b80d2bf3085bf373ed7de2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h639a42049d1a8b2ec577f51c3f36eb6bb2c61ee6b913491b8f36ccf81bee4ba050cb9c97a9ebb034ab76d843fda99f9f9f8e9bcf3ba9d8af907a05c4063b04a8f6e358301947b5b08b509e916e0a970c89cad18e4039be1790dc1ddb783a5ad7d6b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h535d41ddf133f8b114c01401684e3ba0ba7315d05b461f453476ea5f03340453520b79979875a9b7f728a88d8b1b4a731c054755b5b93956c31fda7b1c50e8ab841b6a5977ab1e11abb2c30e77d1f87d45c1b1e37273bad5140286a20bad895b092a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf49a45fdc4bfe98bfa4c3e4b05fd47a21dd47ac8c7f2a3cb109cdc3646f51bbd23a8e58012e77baba0c0f7d893e5ffa47d879f8977c87f2068f66c5e4c72ae8a28d30d8b49bf984ea5301ac4b8bd9c964af3875d3ec161c5964290ed1c08854d4f00;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd064a6bf60538007c5859c0cd6bda511f13902124105ad42ce30caceaa704a554ba6084ae5421090e0daa1ccf222388548ff8c417288c842721cf5566937020dd9f6149da9d5ba54e524220c8268ae50e3c4d15e97a20a5b0926213caea9d419c0f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb27c09d2c1ba2df04c11eb1f6d7d03d410d44b5d5e0c64c67a5fdaf0e70ca4a7b3d808fa4a280e1061aa2ee8219b8afa367a5ae5f5830db2f40ab74f63bac42c4d1ddf0844604baf19cb266525c44b788eae40575483bbe19cc6e611eb38b7acf07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95a557a42eab6e690bb108b96fa5bb2f5a58001ad238bda25f304bef8e394edd8a3c6b8b8dfaf1fe3a71c740a9ec0d984f0a1fbf3f6212191416eba681e86bfedd38659434645639e0a516a3b12ae1d9dddde315e8dbf6e213a82bc120c7ceb9bec4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h893bc97c0e4c28abc9897e0bd4c834eb7c7184ea2b2906f9666e8446921c59d7a0f6aac0dd4693df0166abffed34790745fba9455248550e1840aa6dbff35f1cf6882cb36edbeffbbf2eb5e0c16b8f0be19cdeeadf41dbb047da0eda37d5c0004423;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9a2779655c449cc82d96b290abd215ec62a7c090a16a6b3f3f60856b0702c332056ce89a0477581ee58a005cb6996e456ccd7fa01b715d7a94bd98ed33fdc2a2eb04d3c5d068b1aeea845f6d29bb98213abe56dd17c84a869521de47d93fe9d240a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha15807e8324d1510d7ad49acc441d614fbd3427ae7c9e0c888e2befbe564fa4cf4a518e81dbec419ffd6169885988f4c82e04fc1d0d419c9a0c34758802973c9f373d90a5560d3a1d10494e8eb7b6e012b170c426f827003bed468d05ce618456819;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc71f0eaa17a212b31999016cac5dd3e45dba919ba937a18d5859189cdface83e264b16c4d2b436ab8ae38dc3a2ead15a9237991046e9879f4c5884785fcdfb529019137cef8bff76462e6e89e0c7dbf75c226d05dd1f42f7cd312727f08b0ae50b97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fb0317338563682c4807181c7a8078fb4fab380c256d279d3e52876d9aeccbb32c6116d77a5c48fa501c62727fab324e42df0ec044407c1749d1d565fc91d5f9bba1c1dc3e1ead7aa9d99465c13fb2c95ca9807608d9b77f00ff05d011448b75659;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3193ce8bf603f3e3a0a6e5e66f9f541cbb929acd884b146b54b081ec1ae9f345f424172864ccf8d20a7681941e01d8e9216c8ca5e1065fcdc6c57228f3a73d12a5de34c92ff003ccbb7683375edee24cd8b94a10306c4904ce618b72d021c216b677;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9394ef7740d693396498867e22725c7186e521c4dfd5c18d0344190abf4fcbdb4f220a42b6ef0c0bb29ac2f19e5589b51f921f9c048230ffb213651186afd0ffae620afa857924348a4d1522aa0d30304f68c6b0bf819e2ab9ebae7b5ec65cbf477;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha541b9c4248666506a63ebe35a1379bab8f3bdb1de3be3d3ae056d280359dcd95927e8209b5fe5631c39aa141618ebadfb447fb74ab3a216e383f782eb8f639e5e318a451dc0b2523da4afe7eb9c240e5ecfa3888ccf3fff8e610db54e4db3d1a388;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bbb16f6297555ca755c2c767f4bb745233d511fae4a1172dbe3c1337f1207a9107ff40fbac5a73cd70185d098414e616429c55bcf4a78d4ba6f848945512a1aecb140e8388a7c6a1caa68e239d326a8f629221c6b82a4132e1bd2664d8b10a12eb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9166ebb7cb30ddf6e8ac3ac8e0a64fae4b34820172c5327ef94586d8e7df4eb51fcc8c822aa85aa878ed17619dde1b82dbd5001ca2564412afa96341bad5c8a5e915a4a78b7bfdf0705ee835ff7af500607d2c49ca6e0b879d1910d1b220aa2ec4e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb41c7be007b935783558611bd954fc7c58f855298d966ede2ee3755c5a8f3f8da4d6ff9d26a19abfed75b3906b5e37a629c507de55171947298b4c44fb22b3e439ccce3b10ba67b2ceb056bb4b8cb709c738d1f180a152e096e18f605da5d042fc1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e9e4295c9f95f71a1ec9b7f67408201f14b2818a3a9e3d70c0a93ce6a77836cf0ffdb5fd97fcd386ecbacf13b93df28aad22817d7db79e01135e2397df37bb28ab8094731d58ccbde6ec56aeb10c83f32b0e9a05f3eb0df055daeb5978b1af46d7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25b1682ed9e4c13dbb1b9ce30a453562b35d2404cef636cbeaf811c75909633c705928e20f83611c2e3d8926501f8caf6f5e232888ffcf3b8b72d767909ba0759f03a6689018376a33f55245e5fc09647d362bcd20f6da160bbb929efc27331d96d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde06fcc0c8001dc57889e9bed4c81d80e27bc757602b7cc7bb0d48e40d0c8aa8ef9a720b0485c5a50672907f0d08ec288ccb835c4dcd5b52da5038dfc8efc6641b28748c4561799b09c4ac57ab7b2de0a877961377dba5e309ced860b0bd9f80a141;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefe5fff066ecb69dd8dbeb4064c550c8813d0586a7ba2f2a889cd083f222ab98684546f3e9c815cacc231d5135b741ee1b4a457b1aefa4dab6f01aca8e842af49e00744fffca6fe3269891d5f26dec6e0e1d49e3bc1f7e9a6aa3519ff3dcf02bfdb7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2a7cd59145def884258d5df9f5a7f9f3b18f1cb9c619373757f4494d01a48b848ea164a99a457bf9dff3890eac204f3ff0965157ca5d747ee883c9bb90f1a0278abc2833527c2d792c055e7f4b00a957c26d6bd884939e26ac3afe3cf9c3bb4ce13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77d83c09976f98378917477aa77bb77c1e404274f0536aaffb80ecc6618e783fa39d45b5d19929cbdb58f93d1e5325f05bfa4aa98a8c3e52cd292d6b30f2aa1d0eb92800e99ee03fd2e9a39a664eaaa72614d6a1ad0654adbf9dc5664abe9b5121d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6df14408b0efb2b27bc91495775e09aa47c49bc124a4e11c4be6b7fd9b4c7e83645a4f11b9adbec92d1e0e79b95ff689dc84c843e409c21a2c87f9d780fb15d9a8c2806e40a4bdb41ebd0b3de8c524e412d3fd4e7a298d3546433fb0c863aefaa86d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62edebf67eeae635a6c53ab1109eeea3664d5a269458994c80e6a28c6a7f8ffd9b99890ffb04cd5aa92a3b8fa7863afd00aa6e87bfc9d5fd42bc633ab43adf72e38849c44e18eccc4f0a6fc347153eb73a461211af80482ca16a73189475c6f5066a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64f03018d3438106710bd00c329962b8f73541a15794c926cade233c07682e4aa0947b7b5b844366af51e0fc6feb0904eca2175b521fb1c64f0029ef68c87f06ff54257387a9a0376b1814de04da1e5ddd8666aaaa964c5a56efe7f1e30ceb0f5579;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4df40d7ea72c6aaebc25e44b0781baf32d7b09684a28008e5e1193b59f32dfaefee88bc530b6cb45bedc8bb9749dfa4e6903e709ceff7070c69b92e1de4d5772058226bf9d31f717ffaa65049006707146f4edeb6982a5698590f07576edded726;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86923d6c3b71fdb581a3d2f1ccc9916d740270583b55dd6fdcc7119f9cb16831c9578cff2bea380d1a84225360907a7b36d35fd9e219fb9ab3cf6f0e0772fb58257a7f25d6df2812c51b5902b04fc19f0b005d34b5d89f60af7ad522226cc457e5b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ef9d1de515588edc92c4a1415dea0173b959914a606993e0e887351d423985c9a08900658d82d0a7bb763ffcf5238bb5036e0de6900e2803de692ae4f2f57af2f27c29b91a6667901a4e6825fb0f9fefc23fea62a5d9149979cf80e956e5058ff26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11cffa0c6fc5b6f03ac06e706a6044ef5b508ff59bc3e5fbea27ec331e0d7334a4ae5b5e98d40b0cc15c55ced631032039ec2472417b78e9e8bfa1d68e12bc5dc8ca01540700cfc88d8bc3cc76e6d0adea925a1e02480664dc06a6604fae4f4b8139;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ff3bf117592a508c3d1a050ffc3506e528dbe07e4dc8fc15e4b844ab8064b025873e33ba7860346b1189e1601429bb264a5c5f51c8fee4b9e3509103597f195f04086d2d426002e444cdfeaae673ba79e73944c8274fa68392d36f0abc455abe281;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5d4ec843587877ac70ce17f76c60c79d5d0d7c9feed38153c6977d76599159540c8d607e21669f7eab7bac64bd245934043a019f73529324f15624314dab9435be2e31310d656a37c390399ffeaa5ab1f671f08b6c3d73a8dce7ad0d93218b8f272;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd226cf3980abf4fcefb85d799ccb0066d7d6c79fb39a1fbf660d190fda20200187f40da0144738fad77764d50f7e1bf915a4cd59ba7cd8e65836ba534a0a893cbb1cb0b37340d5871cb7e293bdfdf5038c93b7788fb8f96e79cfdb7acc821d347889;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cf9b7bb365efe1efca3b3d74e67de6509eb75c27e5d93675bc20d48aaf4355b77f4cb0552ffb44e8cda1c00fbf4d6991ae41cd948b0d1b30500ae63f895e4c4b300a66198e456e2cefc2225f49525e38cae0a5ba505bfd1f4832f126eda23608129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dbf4f584cb76f21354264e1baed64bac32b8a72648b12176571f73ce52abc368aefa2afeded4a0e795b253bc586f7975de3fd475c7a9d6b57ee43c92cf84507be2c0160d05e164f075ec060a71a3c1bce0144b18d1164c260910172afed035fdf1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2261031780bd676126400a3d3ad5a3bf4adefe146ef67cb7d53f361e2ed9ae21ee1ad67688e8e8ec777efad3a21cfcdc6f2f82ddb2478a0250218c2e14a0aa310fb8a8f3f32d34602cc00aa070aa63ec4c815a24a4e2ed17a5d1eef456a70483b0a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1631166a0ca9fd7d778251c4c71361f8de51648ee657fd0c3a0c3cc2e8aeac6729aec4cdea969a7e18e254f33a9a985eadb0f35556750f2c36da54cb1f505d48b1acf9a7207734045532d9d05d4d7e752e91afc7c8a3546bc2b1eccfa63d983fd29f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73d7402ce8ed570d4d3607f4651b31c03986a9c1d506912e7c12fd920a720d7a29c4fffc022cc304da3020bddacaefb15abe13177a3ad332c9fe578a6eaa37fbe8d2002f976db87001a91d2c63e501b3cd474540c37c8cdb68f2b7a74db772805b7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2412fb7033c446b75c2a3b3ae093e4180c3d1f253b1b19cb9358b7bd95599486ebb8c723d868ddc5900ab255b1080d29079a076434a945976e72f25cd3f2858afb9991392790400b1f9f862472ec4a2f98fe7fc90b92020e89ea64c36c2376f32712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heecae2262838584acabb453ef3a003e83ee658fa1856aec5e52e0ef69615c51b5894ebf69166d7815f234279147e9adaa6a149f61ffd84ed03c7b61c0f8b2de2304625e54d5d41dd109a70e420a814fdea9c5a78e99d4e63ebe55ea5ee8ccbc18a57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3b06bd94b5332783dbc38076ac661855ef14db8c19cdc78a2218018a8051045e2b6906ba3cae13ce86c87be210d8db7431854864db1f6a14cab5f409efe90a0fea854dec038e65b2e2d1cb1fe8222583d7cdf045790e9f79cc3ba87cf872417b9ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50868dd2d39c6379aa3881739ef240c0efe2a9efe43774bfffa160727a957c1d57f72bf9c751e2f10fb92318a1557584c8f4505a89774ba61da8b9344c011d8158af31eef9356ef50303da8fd80da0bafb66edb64118920a96e9f9d5d8348998657a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44cf8e9a4130e0b2934284566d7b21f299d814a01b32bf189b865df779b5452463174fcffb17f72b8cc5c5da7036a0c0213ca23226573865986328563e05a820ad13318fedcc5ec68b47f94057ec11c46a8aa55b4b05f8eab1c179af349309b964d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc5880b95c516ba989f0b28a8beb8dc80b870bab0a6350381dc7c78e9f04359cc07c95dbf365a0a0f2a7c990ddeab8e19696f3720e17d88fe4c70218599cbd74fb685a7578fc48b81fad855962f8f1cb7ba79ae5a43aee5a0714c22fa73e2f345db6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d884de35f2b1cceaf435fb1a4c3361880bad1f712304ef328440171656fb7f979cad5255e24568beb4249efe72c8a841b1f6cf0d34ad5dc1179d3226c832ed753488f62048c604bc4aae0b37020eb3d42b21c5c4e77e49f791b32ae7271a5c13de7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha389efe2a9c0ef8fd43505c601d31105b721bf529d35e9c84a7d8707b58d9bd147e63b528fa2cff345f431b05227ffca1092ead635ba881ffd4c27e74e46addea0dfaf6d05c061cc6b5b84e69d3874a4417be53e296d80cb9472b6d8e4b885a25e55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14e9d1a20c9bda98d431680d1c5afaecaf4c31e629e84f241555e7f0390f1da7e1c51146ba8d958c4920d3dd12176299f8bcd80aec239fa3a2aa5c720f345a7b6a3cd50240cb9ab435225ca771f98a5df85fe4d54c8bfb76e8e79f10c3611728ba86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ac3c21829862c3be16f9b9be1606ee221434af0f3fef10a531e36f4b42673e8c77cb278f3ca6867feebafec785ccdf77f373737be57136c71a6e3bd085761db754a83e6224c0563726a6ce358656a242bc474b9d6b8a0f93f1f86d55832f0fee628;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc48d91a0ffa9ae6dc7df6f9368b89336776ddf7fb12e0980004713963eb948b18307c6b48e71dccdbb74842f18f8ad91d312822169de356d5e876cf1a66bfce88c056d2868558d4b9ee5ee351e3eda46842303ac6a3f7634565e70cac1e2f979ef56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h872ecfc394a3a5467ec8f9777c241551426fa3a60a12593412fa0b3fd50c9d0fe9a8326e1ae6c6208c386f6326042d4c82ed67ed302e1f8d2318fd3bf5b0ce58b76bb3c02422b5d5120c9352915922478e0d34fc3a76f108a9728bae73eb762cbff1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h972ad76bd766147b344f3d5d16d5e8081092f034dd41318195eda682448fd89cf56011f6fc92c933129a49940691089f868977026a54c449e2d63aca00ef9d4b9a19dd448ab115d0e108fa5bb6f5d193dc2d1b4b36680efe8b8ec705971e53e0b35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h784b1dcb9b175550c0e47a507989f6130952aeca692f78685ba20aa2169d14163e1ad054e32e91d3722b941163f501352a72a057bbb33e4410125f2bf1b000b0c9e83b3db3a4bed15188efa36f70914be5af5b9c77f9fc8878148abfd1ffc75f9f1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe84f3302ed9de18790763e8878ce7c75f49a871a406408599aabd2a7007977ef01862d6c2fb7b453cf2c50bb0387fb73b376f32a847b2a78938fce3814e20aa0363f6c08b4db62680cd214b4defa0073a832c228e33462d4c5682bfa44787952f08;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99aea1508b9d0f4031debdc0ad99373f69fc71d84e9dd742bef5f64b9d7a5cf079f423cc13d46ef223a39c147f5e65483a6641fd17586578cfaa97f6e56b0d08128bfb3a0b7bb670cf31e8d82eb960641fb5c096f7fd4b557ccc8fa00338d9193b71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba8a465696a8662077490321fcdf98a9b43d1130700204fd69d59570fe3ded437fea2f6f96eb19310c055e22548162249807c985fe0fa69a24aef9fa3ebe834ea717dd3d3888be1706853708473066532ad10a880b551c627f65c71825be9a912b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb62d9fbe5073bd5756bb38a8b02d987f174f43fc1d182eb518673c4448a6ac034cc89cd8fd737517794d8b0dc18fcd2d541bf7778be8879a02e74a7835554abb31d00c0b815f06d8214ceadac200d9a01692d2846c8da162040291be44f053fe15b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfb50e8143fd5e4dfd6aeaac9f0664d7207de68332eadda60225c18d0186011b0277fd7d5aeb27038763169cbb8e8103c42597eecd3e6204062c5d6cf64b1598c72d04ba55e781289355f866b4be81aa0b0048fd278107e651051d50fe75ceef99d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf0868a3eaa00a41d813a0f797b82ebd48b6bd9ab2226c1aeb94092be4f242c4a507da8af49d0441ad8375bcfc5857ff7c61a091a16cb24ff4cedb902740229e689630f18a0264ae2e175efd7d2b8015e2276beb9d2d8c4b221cd9d78dccf08da770;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0dc6ebc66364d78bb4b69bdb13ba431a3a11c50ab438da2a861565758da106b7f30f2f3239a460e23bf830e9657a378c4361207f494da84150e229d50c43b4c0469fe8a818c22ea1237799f3dfa82f7e3f29e57b75be7ed77028f1a9c305dc1d05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9e4475a8e79fd5440e123a757bfa28b144b9ebcf1646e304acea467edb85c6de4ff788f7957d7efff50107edecf952cb59846c6be997f3c71cb60805d40a899bf4868ab349b258b728d5450acb7e9b3a2785b87e71caef8db8528644471b506301;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10dc8efb98041545c50692e98e34b63d84808c7bf9d547e7b96c99e7f1814ce878a9234a50bf30ef4197b2d5acfe9f9c363ee3e1219441d5cf1d5bda55015f72b99b9a8006e98f1e894abe85922db201366f4d09bd124440f61683ba1a257ccd59d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac6ca8964319483495f00c464886ea93a4f78c6d93b6cbf697b22979ed5506c81f2e12090d7ce16ffb0b81ea7bdef31527a2fadd1acf291b207a52957d119ff288cae395cf39d6dabda9035ea47e54cafc6479a8784c428a04bb6c2dece091e6db3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66a0ee1cbf6a4f87802bb3a6a8a3784dfb3315b57f90ac3ce09579f4038fc251d3cd355b215c20cf0ca495aa1195e206236d963734d9a952b5529aafd5909cabdcd14a5850809c95dfaa8c99426bcacc55a99bff4eec023d9019e5bc06560c46e75b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1fd4e588f311e9ad5bf92c96d12102512c04d54aa27e00e78bb13ded271ab31be6a133c3c8df318cd589a7d6a0b67c794e91a0b6a1686bf8964926eeb18b5b589b81aa6d101a185f9f1a86527ee6dd779638883a7964c211748246a95c7d302495;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7151d4c2656d6c22112bc614466a860ad0883f020e61f8d919db93a70bfdc991dc74f07bb33a5b67d3b742e0c01a05a8943073dce817a97ca4691488e748529961cc5af8dab6a7b81679901f729affc54819c64814de51509d442109448cca1d053c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f29a23fc7f7606d36c53dca128bd615c4942ad6893cb39d7bb7538509540cd764d252f4a5487fec2690417588e53912223feb007bb4f67955a0efa686fa451e96b3ee651d15a2cc417b6aa3804a6bbfe7fd9d5d5fa30395900b343d07e1df1390c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f32fbfe310d8b478b1aa063066cbf5d9d16cf3b7d2f3ca6b388e4c438dccf4d4348aeeae50365d72f37b2ef2e2bfd93c727cac6649662285a46bfeb74a46d63c8e9afefc002bb3a14a341c2a08a839978eab616b1273fc50e8abb213e36076180;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h239714c4284693a93cd15ba3c1863e80ddddb4197487f051cec7eb3319eae04298877964de82054e656703907b4da9117f9a47c42c58ae4fa293cf18ba16d6a543911675490d4cf2282324713370b116a9491420181bbf9815eceec74ed084adbe35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h916659ba23fbcb76148bf1ff2b870f69604873650ee40af90e9535748f6dbc7408ece93cc79bbeab5fb3ebd4155c63980593fb3b4d44c36a7ff066bc34df9bb60d8aea22c78ddedb43452d14f91567073fe28be7b8298ac64532f8a55bacc0bfbfff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1726edacf6b529e7388fca7e0785b4aba5f44b30c75298cb300bc40669d2bcc07fa4d28aac7182f3dfff7d59ae5215abd3e60a7d90e31157b3404909cc99a4c0fe3a237193b0b969b661921cd720f8750aa137fe4769c6327215e2a5e3a4fc42440;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f3be36f162de4e8e33399314daa09239eb66314f77ebd33915e757664b90820655d0440d4ad0830500035a866a9cc09ffff1a7ef2da0df3e0c32e586363d5cd296f7dbc81d42b06ae4efc6887291d4ea6d54116228700c0eccfa780af4dfd80d9a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a454c5dd1d32904eee98eb2a39d6a88d0543c88179763fed02e7df7f366d0f220fdb18ba1f7be22b182244df77b1593cf1ffaf84006831c341fe510a61e571b02bc63f117eeae29bafc38beed9199380223afb6988c75dd498aaca4d0dacb74ad16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h673be2cc97bc3f0fef474d6c1accccc3a764d1366e8417d57bd553ca71e21d098c6eb0d3201c635042097b0e15e80e1b82f7a56719a506272d751b632957f0a95d2816c6d00f1e81ff3299292074d116dd2eab6d3fc79c6ef1fe835d9d96f072f182;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8134722a85a621ea1853937a4bb2658a0bcfc8b389228cf0a3b8f5d5d80ed2a219770e0b7893fa2f729813f9e8dca11b747556c219f9e3692089da6f04771a2a1f95633fe2fdc40e8a3d94f5d46257648225c9220c97f7520c4d2039b0beb07be5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2eda669fbdd601c52ce1f1cd2f5e520a696ed734f83b1673879075db6dd4114398c634cea78f242020f798ddcd40d046c4109dcfdceda67481dd7272932e0088164197a9c78e26f98fb4af0e48cc51fdb5ba6110ea612d6ef5c20cfe89f0e00af23f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe615fbf2eb54991c699c5c4a04f8b366046fb638d67209396720ac4091c6787a02a20a5abdf8236234688c5605b6b4e2086410702f0188eb1b8424a426c348f198abc88a4a80c802c4a044ea3ad59414a5ab1c6bcb8b23cee744b729d6363ceca3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha78fb84853e7c87deb2e87cd4976839b5432e53a7e51b5000f6d2eb44f78bb8e4b5a5c1576cae0e48c56fd7284876997fd6e614f5bee52601a82bd87587b5f2553c5f01650b63ecca46e0020949f55b54e330183267ee5ccdf8d283e661d01f4ceed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8658c88d9f204048d6f390f3e723f6a9ddd425f8701b50db21e2f33cc45d16fe02dd83d53323f786fc24f81e92824d640a95533cbd1ff6e6efbc46dc1ae5e14f6bef7282db32285eace77a8ad0ec477042c0e4130bc963a8355aa31743f6aa110bfa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90812d18fc45f63581849789d673efdba9ea96372b5f268f05538e2ab38cebcb1f3d6e5560a3cac83ea8b313cd5acd460c4697177a335c9484e02a71e6695cfbb30f85e3e67482a54538eafff7e06de3ec67a86081adf832c545b4eaf058a0173159;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1f2645d64fcfbd796ca0a62beb01c7fb0fd726e2f7691258253f70b685cb8c6ef6e325f2b09accccf773ce6ba9a52e6a2d7d30c645e092dee9744fc3e654a5452f9ce1def7df594b0d2e82c3d4f9f58bd9a832b3023529eddd22bda487aa044dc85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41ac4c27bfde7af6d097f74197c6c624dec5e0237ab8daaec71f257311b2f58b6f68cf8ab105bccc05c7dfeb687291fb73c5972d4ddc57246050bb8ee14edc07820b4d560e920fb423eff64c5f30bdbc9c9f206a80d66a8a30cfc58212d967fc52cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8df8ba4b09d92fff941aee0d8cea42f565fe924d69a87c28a95a378868b16f724e31bfca13bb6d6989fbb7981fa1078dab04b4ca622a4796816664edd7e6bddbfff8a19c2f611c71f9f738046bcdbe6523ff50a087e420f9c602910b77e96c7fd4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab55ee81a232e7bd66f890a18596f037c9b2a3a2710df5d8651fd63c5f05ff34a229a005d448c1c33e1499c6c0723ebb4219a7d38b0c0f21df735958aeef19188d3a971e9163ffb07c1d59c499e2ec84c985ce539eb2fc957864816e70b8e101321f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h746bc01afcae48c6d315970696dbb5a64063610789548396679b9032ccd21c6274f4a0e09e4f717a41c86fa89a5f99c19a96952a52dc0a477d27022d373c278c1c6bbe766bb331d66c8ceb1234173a6204e7fc006d2675c05870fd3c3d4d4aac2c4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3e2dd86c995bbf92557d0de1006849e0e7f3774273cf06a2bfba5c7be6ff6db85b35b2dbc29d33fcc077b7f1fa1b676e1a722f0a26dcd4a80e016b1e8ba4e6861cfcd8002df07fd132e3ede005819a003bcd74bcf33006d79067ca5774ac3b2ff5c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbdac80650bc6610d0347b5e9d13b41f826cbf528b46272eadc08f9d999ab9612547d7799934b82f5ca45b2e3a075d6893ccbf8f369bff29c4dda8aea43d319eac7054831bb031ffb14110ef7fc0cc14abfd49ab7238de6eb0194d2b035243f52ee3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfaf17314142a489b26fc73e8c6bc5db2098374560cbd686491df06988c8f6934d8ed070dac45f86efd857922e5003d686b43e9ca64ba6b3b599c42f579dfc93b2ea484947ee89489798611c7267ebeb894749f190a9bc31fe2a251f0e54b61f10ca4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0da3ed1a03d5653535864d3207115e57ed298f395a18419f62c90576968b52a8566b7cbc5e53dc3f9a55f627bd20c27194a28529498ed45553388e0e6141898459b33ba10fc23cd5094b4a5935efdaad2f0621ada759db4f9806dd562bf3ecbd5d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c7bf398d3fe0ff30c6e4296b16c54e7f822a79138d070be5671c9925be9b6fbc5251014db1de7b38ac1ed8dc4942c56bfcb2589455d384d398d60a135f13254d2a35847b17228d46f06045faee0d0d2bc9f8f0dd0c4b135256ee163cc92167a6225;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cd2516d93290965d54bb981c6df497f580fec7f70b4c82f538e6f29ebd9cc5141cca541edd20ccdbdfb25027a9f046df7ab960dea6b4dd4ae967cccf90bf6742b95a21b30ed7f7060c2c71f074c767bc98b9f52e533d8e488bcb5acf510eaf1b12d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81f5aec4473bd9d5ab32d32fba70a14210aa808b0e792089a3d111576d14c93e3afffc25923cc98dd6d355bf0ec8fff09b013591b65e9ef086993dfd61f71b45301f2ea8cabc02c6a6cccbe4d910b3338192d6d6a4c6c3f415b8cae558b78f5c4a92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf8d3d1f6257a3fc21b7d333e50768590e9d269b2f2602a977178f3845d659069f7df4dc58a11fe81ec21cbfaf22a2c4a84474780dae96cc2a7fa54085065191996a9c9917584ac377972edbf20542bc8412cad521c29ee461ee92817a1580bb8895;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef07de04be2b274ecc74a2e59fb0f88d3b60f50c11262c39678323d80213f72b666b2ce3011b32051f5583b8f4af5e873d174d972b9741114998c4c3bec3ef2779d0ffd250e2f0f678ef06ccebe4234b66a072d2cc9ef469a50ea0021ba6647afdd2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38897e880c4bd0afb1fbf03e90c3c9001d93bcb19afeb394e0a35f9805dd0169f11dce419a4bb5cbe3c557ac6299e10ab6a0a1b2744f9fe4bdb81c94cc9455143d2683bbf287bc543421e6ebe606addba26a8bb53819f08ff9884ca797df470cb8e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h896f0f2ad9c8ccc690a998728619f626012a75647715971802dc79c3a6e0bc14cff8175e5532fe62dbbfd4b1648b7f55a0556a1bd1ca9d702e0d5bb121c07be00e4f9102a87d00444b236b325e88d809f3f83aed1f66847075dc83f433642e79f10f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee99006e59641f95e5820738762acf6b554d5e9619d6879e0aef8fcde76640d7573d66d39751ed07a6dd39bb3f50807138c11e5f502a76ea5cd0f8dc8688eb6856677adcd61c53f947f326a31ac36ce0de9d4730a6046d5ad84f4b82f01440afcc6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h714612940201ee7608f4acc7aa0eafd0daf56530da8da49523028afa32f7bc2cb54a405f7bd183c559e4a23cf2b483319ff9160d37dfe4aca340391ee18f32be331adedcce16740009ac88b37cdb7d7689521d4743ee12196379065017ba0d49ddc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc32ff025d526a5802c1a59aa3425968eded2585792d728d06f284eff23b1aede8f108fa6b52a8191c32332f98ba4ea9d980e04e9d9d36043d168bd14e42d0dc479ed80a219df05faa5811fc8a6984208be5a7bf5bf089aa3750328419459f51599e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96bc26bab57ff3d16a5f1b62246fcc36fc1499c588803657e40adceb15bf42cbe3a3d0668fa00398da6f2cae42299e7e4f5509a89986720fec65e300aa6080dbeb447b398dcf9c8690a3cf2e48c5973578af71d3c69cca26623f7f2e67096a34d864;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bbe24cf33b9e61e6647e96bb90de7b4697f508115d4486c9e158bc5312bb598097dea70f598c38874fa67505562ad12959d4852bb0de62827f9705a61889d44dec2370ac3edb2b267aba12abcec69e42d6a672c971eb382e5c996fcaa5ba8691e80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7aa4313e4178f534745b76282fe7119027b419f3f20b7b2af6b7f7aec5c7cef709ad3b4adf92d00119dbcf2e5fca6404e8fcc2f8af67c5893a14b202e1de130acf84088c868ac34555f63acf1a33cc426316f60b3e4b39b3a256f0be35fec3cdc9b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haac282d6a030522879fc5c004424a9f4a8c4cac08429fa3ec5d0c98694382c2a8932e7fe22fd728c712fbd0e5d7c28ea17e353100344254bf1e1b959ee218d759a0c976bee60fcb734adfcd1f099fb53e0140f1fa2b817fd68e1839122c0af9a74f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd360fde97288986500073f3f46d770d11d342584347e1a771bcea4895da1f38b446dd767b4510307278ed6fa7d00d40a9244f13cd80931ecfdd558146c09157426531e1e8d6572e02c2df8db0aa7f0ddb819fae4f8977db9110cd76faa426fcd527c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he74cbf5f0b4d44b730616669017812e9efb13b72458b52b758e9a6c9a2efbb9378672748a3dd2c915b0570c8230dfb13d81bc92924092262426f0a197a699fbb4ab067b2462c6384012216658c50ab19316d153c53bf866249fa27a90431030a6c67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h484aef2eb423ed9e4919c2eeaa81641c969de999deb20055e2bd1b0a65b58a00bf77b4d812caafbecc62dadf4549fbf8cc9292bfe0f5882d0148522e941beb5b18e4adfc0ba80be68c10fa3977211296c873144e447b350eb5bf23b53e4e1749652f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbed1b83a6e69c31f2686d33beaac7761291564db934b218a2867d4840659d86e96adc3f6f9ccce7bcac70a793c122a0f49a300143f8c5cb34a5eefccb02f072aedc56360f4a42b9f32dd7dcc0f2fb3db0a04c28638b8a7e611003960fabbd7545b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4fb89c4861b26c5c235cef05fd6578d02ac9673663c9c12e938a371eeab2e2c21a3f88c19b9e1a5fe0981ca70c819880cfd00e8748aafaa24547d421a352a284f5a7c95d2388a41f09f09055c6310c6764e5cf44892099f4675bddca83007634d21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefe90a3aa394d42b9e61e7535e17de51c7db98e21b9723b2b3bfb314300cd086f771fbf22fdb84ce787227d2c71da7673728a869e7246be9a4eb98a4eb47e423ea78f29a3bd42405c206052af8a5bcfe2d91d6dcfb29d9bf56d14272bd957c44606f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h154ca5c09ef7bda95f415fc8b58c887849919f4a9a83e23e43cc5b835c50a3f3bebc0cb10ed9dfc30d7e7289e9780aad4b48060ecac7b33ede6de4d9872232b92881a7d4a97d5b4e2bc499df9cd0f6b5ddc7f7b40b3ae29a5251deb3fffde1d5f8a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fdba902de5435e5b0f3d4177f9ea6f19587ff9f2e3fa98eb42806ced9ba26839d5deccf1a6d78a9f13ee18bec2fc140437ce702b0e931e92a267d62fedc0855eecb0f67b7da9c2c25a9151c0ce9fa5b6d563117df9eca8027f9ccf0a8ba904ae3e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8c78399088c9f1b6ffd947469b542019435932f56c110763f3e24e648dd9a0731f6a8355661d172e677ec5e9d440d02110c99eb9d1c89808a8ab16c82d7c1b4c2cc68d79e365bacacc872855c5c0e71d4bb6154cf9c0f674b8ce0b885d50cce87b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b04c755442cb312f05e7d0cb3de63ff4805eebee9e337d9e3c36b4e116c4cf9f33fe865ce295d4013b90db8dbfd1bb13c9850e061c722b75e74a209efe803948774621a095346d0dac673ef56545726e499e2182b9df43d9916ed34eea6fdce7e44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5005b582c802f95e71e323c57954af4ef6acf436f20f337496c59bf8dcf1e126846525d1f50d6af3b6d7bb2f354c3b7c459ea06db4128472cb11243e85a326b96fd861ad8b6b98d7c4825a9f7b131d1fd23574b33bf6dee7f89a8230818d97ed5d87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8644dca76f4b790e77483f0030eec76afffd10efc6361aaf8cf68bf3b3a7bbdc1b541244ea9344b5703d1a53198a17075d871a8fb2486e48a719d74e975fd4b193f7d344b73914def0b2d9b40958e6bc9b9e4369b4d8816aed80e287571dc1f9076;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff29e377b54b15bdd38ade78b2e922012870381cc9d63496c55f0b0577a078ba703cdf26434b05450a4b1cfa446b033141f3c5b70e074202ede154e54805b65479099c6b2505b39820cbc30a52780a67084d7d367f19fa3ceec4480a85b93718fc56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d7975fc3fde256d8b8cd8f3e0ae26b33d3350857e52b8f0216dcc9caffaf79dd85183736c30c66675ab49ddd273ecd64c6213bc8d55efc9819ae0a8ada8b1c74515cf4fc591d64bb04efb998803d56b9914d7f92470126f0abe786391c7d2534b8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedf19c9e6ffb87af6623e449670d574707b3862568564c8d890fe63d3d2c31b46e1c54ac8854deeffa3c5e6167a9277f54d52d37ae262bd7d57b6a5db64d657f781edbea35f90fe6d3fc3b2bfd7df51ab7bfd41c9dc6c4d7c1ab637388f557a7536d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50e6d564aea726b607fe4e64f4dc60f1fcc6e04c8ccb1905d7290e9d9e5cba9272abf7936d336557a13120ac15b6d8f63c441f639ce458d4520bdc38cca9140f85244a59cd76bf06dfa66a961e3fb10f65333032914f0eef6e52973b26f136ca6603;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72e3259f7893914edc1e9edce503d4067bb2886440f7cb82d144191a8915365318225afbc8ca8ea4c3cd36378be45f81edb63fcef350ef8db8340807bdf729269a587f9f8748275ac275767f48df82422803487cf9093eddbe1051b8c953aa2e1253;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ce2c18e84cea0443a0a7890ebab6506479be9b68805ca9df83ffeeaba86e647c2f4d4002bff8c559c1f691131fa4423505035a99c35d7fb895c171fe5ddb769c2597fa1d2ff16cc2a5c9a94b4e51026c2eb1624f88ed8f54ddadda8c94394fc0190;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe4761c4b1c5ac61bf0df3debe76774487990bd1c49db451bee755e3857f2ed67cf3871664f3688538fc32395cb489a76dc9b0da9817433849ac735604fb7bf59bc8543ae9aef04260fb0fd4bbf26c1492ae43c30c75b38227df320249d8a9594061;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9262eb373b82cf91295687768db255d875dc843d9706666a1e111422848c3e4654e51bedae6a4c7d41c956edf06b359f52c49cd717b742144f3a10ba3780a43ad45f667f025c90dd0357495d2fb52577559c0740b2e4909324e22f9fbba2b7d8cb6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d57aef4e4675a155cf9728343d8e7b0c254afd3bf261e244a721845fd29de5c1b0a04d4fd66219e285c55bb7340c76879933c4672185e08ef4f384fe9ea30eeed20b556c9cfaeb24a7023ee251f6c8ba71a0ebb6a40e41e3ffa8b90e765f7b9f158;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e8e4b48402db4f61886e350bc51b27b026fff3a37fa3461edf07a142a62bd0db77a7ac686f23686a42ff67cf2fc825aad18ca02c88333c4fd0930cbe1e0678d5507184b6b166a452d768697402aed4c0fc237df356ed7c54cd610932b90741e2d33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2e8eed4e882f427b23b004b33c4ccc9a9a993e604647c1af4069e4a941ed184bf56d4b87b13c34ca30d52f0f4b12cde0463d9aa8b8862a9a9c9120236ccc566a33a514ad59241997393726c76eea90a7a31251ef575b46908bd115afad77c62432;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cbcbaa8ff170d254f6dfbb64f08cf0e2f7534d7a11e0723b91250a54cffbafc64cbf12f5910b143c6748b9efb837b39c53d23406b131ea5673347802a04bc41144bb0f29e10ed48014a69ad0f1fe33b098b64ca6cecea03e281c4ca756ba4d14e03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h636e72db639f7972b76980838bee3b0f1f67c31874c70c8410cd510182463b3b0730ea846722cde765cce4fbcaff40cc4391ba1ff7562057d7d3e730ff19caa83bb465d787cc4556967111b40d135cfd05090907fd6965371d7b0494c4b7c1beb754;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d26851c0a533e9661fb5b5ad5e080673d2ef2f2f31ab17d15c98a13e1c125e3a0fe056501d0022446fb359ef31f5dd9dc31dd5e2681f5adec6aabf0bce785644890907fd9d97d8ffd85a74af6e729fbca5701dc5c36b39fe5d4416d2e8b6cb3e062;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc39e26e30e85fdd051bb1d8525f5076782342014b67a6945b1bebdf216f80e3607598575e53ff0739335cd987513a460e433ba9c6619f7a7c6be81949ca5d36b737d75b050bf1971f78472e51f44d91bf3d5fad9409731e29c2927ab62c8babed8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45dd86ba150283734b0c8448cc10adecf87ab8071804183950caccf4c512023c19b532e384afcdd0b13d3d3648e511cc30b9ad2d585e68f7baeca15dc5cdfcedf20ab947ae8458251e0293665ef9e730d4514db3cf5c289017e1d389c347c8da74b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6772f2a58bf8eaa1d90461dcba9e4af00bbb4fc7759bbcdeedef3a2b605ed591767fdb30e2950f10cadfcd6b40777cef16cbbd16f94f69af7d7ee3ced5c75ac6a0bfab82b69e3e34fa81d40afbdc20972e7d5f4e2ca9ae007d75a449f7954b532678;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bfc626d2ceb4c3231fa15fe2386851b6affc7e7b73a175a4d267c5f5480a4fccdaa6444917e3d56e21959a6df7a5c43739351344cafbcb8529ae2b209a370674d935925d0f04aec82be035f79d732d6aa887d87c442c43e6a00d8ebd9e5fdc65a72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca4b8a195ac0eb3cd43cefa07e508536d0707f1d2dc874159544ad60ef59df3899c3ffd79864c3fef2fce6ce2ceedd0188f2ab10d673da54b71a652e035ac01a03b8aaf5b14e47bf38bb116486c5c01a22e15fd933122a7eada8c5cb7c54d8bf1d97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66dbcf1ee55f05c17d3be92ed3587ee79869006d293410bb51a74f2c47840069ce5f850984b9033888997a930634a73c7efaaa7e5ce5e108d12463c6c4e5945e8101a92c00b585bf5bf346c7cc3ac693d15a09915e2cb0ad0044ecc1061f1f0ce207;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f1efccaf0d09515eab438236877a8c87c9be840587a83f3fd1beb50d69d3aa9e28bd657ad49c9ba3faffd98344c792abb105b5e2531a2cd31588e76a00a621c12cb3e35b99d96ef4359047457dc1b911a2751c5377c8026fc03e1344d73863dab2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b87d6c4543b9d7c00e9035ac4bd11393de3990c8641daca31ab07cee51852125738ab552d83203940e817ebf812885d0d4dd406637f7626faf876e29adc45ba14edfcb4eca0b17f0a91a7f512283402c3c0e7c735a887ca9f45080ef5fc32682ed3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb66f64e26d65b216d5ecc0e4cff04f21a220a55de849291952f4eb007943434b2bd27bb56a0b92b8cfd4a5ca7ff90a83837c7466cb1e002253cb741d811dfc845b6ceaff459b53f255f7ff701a0cabf2eb480465842545fada0379b7bc17db5302be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c40970b128aa329149bf3b749630eed5c9dc06a9713c7882b679701c9fa6c8cbfe47595d3e18a8eb1e07d742831e6cc1bb7e784e3ad77b3ef5038ec85989c66391736eee69c1941fca26bcaca6b37283e2692da469c588e4b9ea665c0da36a1d6de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h228cf9b761648466f622d7f41d4617aefca6ca27b42ac70baf9b707e9e9bd87f177c9538537f60f07b16e81a627015fda3b2f09d08f7f12795bc3ee51539cd11ba0029ca1d343a3dbb0500718d30a39faafc2111cf6139c78b0930f8f3c1874be1ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb34f669134a234d34a6ebb9535f79484e17a78afcac774173713d982bdc41a0fa5a409b05474192a355c1db30ec329141e240aa3ede5c0274031201c26e7d4d4f46259f9b9eb2dec98a9067c01cc024ebc6bc4a42df12aa2af96700b5a41c4ed2d9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf793c0c5d7ac40637b49072e26cae5997575025e7515349d3fe712b81f436812be558bd126a8144411990077e2987ffa3d59f2b13e2b341a43aefdfb49d91e9a57ccec0f59d7c93dac6aedd4be2a2cb264943896994ffc43edbd763cf2f2f78884ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28f5006d4a8ee3441fc40a0a1d0bac44ccd7651a74dd1d727eeec0653652f84f2f7e589ee8365ae80b86cf68f211e697a19ce6d20fbe1aaf0da67e40a5aa5a67ff9a7d9d22812ab0990631c1708d9c0720c32ec298c649c0e9db717771217f89fd6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3352e92291b19caf8185d2711e98c6b44367800ea2bda0a5b025a78bca3441cd81308bcedee8e3968e5a6e314580ad8a1cdea22b0a2065883139c42c0c575f59bf2e237dbcdac8f30d007db5124c1eee97f6f06f8fddb23690fb39558eb50f404c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89f737ac41197be64df52d082e8c14c1837a7bdf9de9c2b64d58e26746ce503891ce74b6705417995fd5ae10277507bfa82feb8874ca1c2b84a88de9413acd78a54323b9d121d1eb764f20549743d1a3377e0355ca9f0e5f5fd4656e01808a017586;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3198c4d74bcfe2a617719975c9d3a739eeb831822b647478ebae409dd6f13c52279a69eec9ffab5e96380f26ba981cc2bde8df91c681602fc4bb61f9fb5575147a282df13d2d559d1152d6d5eca4a34d8a5dfc0d1d09164e0922810dfeaa59503e53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h479899ee99b5e5761b18cc6d513783aa93239b3db45521aad40c04d55e430c704ee20879f102d3e6a131f378edd17e3432941feb78be261b4176a72a67082e49d995b8d89fb914276f5b2e13f0f31e56f687b36dc4e9f642e0c852b277a3c769f8c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13074bd6f1de619931133e86f83f67473bcf0c1c150528a0acad5b64c0d63305fb79ca203ded13179fd71712bdf312447e7712bf16dd46636b0852e9dba811d86fa6409507d2f55ab856ad2b90c300b063c9a1c6eb08679ae3dd1f8cf60eddc87f18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b5395550fed3d3dde30346324112aa04a43caba4ca34c770d6dd2909a14ba9a27679f72fe7c3497c4a168360c45fcbf7bc25f9eeff58249745e69576c92b862aa92fbcc2011f7a4b0dd489e6c303b6f40b53dbeab0afc6f8ff68daaeccad7ce9db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f60a502c1d5f53d445683b3a33884ddff0883f7757a6ca71341e32a1ed19e4446dc16174d4e30d7caaf7836aae86b1fba655067d45cdb83c80558984979bd4beea778b913e9ddf5332bd27f145301faf24723b8401f7d863b3bce49843b2cb2516e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5516e0fce85e21b5bedf078bc44ba6cb62004f20e2719ec5172f3267abe40743dbd8382944d9c1d400de2c8d06e8273dfc9000369f674ce519612c1eb8294d4d0aab7565567e6a8c09f7a42d767c10e1805357effa5cf81494c703edf89d535d3497;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0c490f18207267c375a143639e627920d496dc7d767ae8c81358b0a77b39fbef6fb9fdb8b883059910fb7efd7ea5590361e1b521c7ad1f7082a670fa4e15251a66a8104f188cfd8ccada4be29d5fd1f3613592f4298b72082ba017c8b0f44359fff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8936c9b6f45ef52fb74cfa6efa035400e2f44b9e279aad562ef538c948b29997dd22d859103bb17e7f93c2537a4a52152263e39e156b6c1c40187f8a244a976e5a936371ec405dda13926f418f783e2e82d885e29dd2f2b09ae9b6e2def9ef12691;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52dee3ae3cacca8bc8728caeb9684c781c2b01b63eeb203064a7a0ccab6999e41b8f0398d441f2f8746d78601c4c7a344c348bdd995a0b2bd45029547cb36b764278f1a864af30c6bee33503cadbe25f73c1fc5a072987164b03af6cd907a38d3dbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8081ce4ab240afe165e8512943217035538907797e86f4c230393609a95ae5ddda771e7f35f362ce8d9028828275d5fe13e79d21f028946e34b2cf1ecaeb7d77745ebda9761cc2d58272ba808594a573b041467d19f2b828eee8f8dc6f54d9b6c1e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf67942a19e0a7cdc6d510207e10b8ddce87443dc454c7b92cfc374212c353d203ec38531fed2537fbf939c267131aa7d141cf3833bc58e732ab8357c8d615c076c5272fecb83ce33a5aa85a1d7dd09c6dd37722fd57365d75f4d872b88351b865;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fa97ebdf91241359af6cc2476d38adbdd889838150438c4913943e389737acf8cd12b26b79c0c420053cd0bb415217eec60d8a6b2a6304becfe26d17ed58b912ac5f230ebe056c07763f4302b3d865c7f97f42c876835ae95357c1753114010155e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6adddec9a09f919c81914eac7999e2dd37f06baadabe70059fccf7d8bbd314c81ab9ebf43b0b927196ab8eab90c5194f977e0e795d901b1ee24754de1949005f709d289754eb504bc0fb7abe89f8105214c1debf98f2b872cb85cbbe684282c6c445;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e9f14080a1f07b4223ad107cf9ba97bb0f163a7c864c5c0e0ff0957ef1f3e682dc9c6a69bf4120d94409357b2b64f78c306cf431efebd6bd484462faf81221adec7f9e6dfa1d75403fd6258c37888fe4e02494a3682596a50edd3a76695b00b2552;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1048af91b8807c93a13d815a16b26b6dea2980465dd3eeff9097a0595a8d7695db54fd02a7e0fed761d2f457b117f7572588f6d7081595632aa3ea3fa94b03402468a957196fdc343691c3edaa4654f0db8c09bafaa669648dc0743b081b430a04bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69dff97d4cf1449e6d090745cd472f2bdc57510f0b533053020c386ba4d6d763f86bfe3d181d4ecc399a7b5007a14ccf45777134c9f36a6cc2e6dc2bc78add72b94fd012dd63636d999304a7216648a255703984f8f6086c3d97fd943d13f39a1130;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h872bcc40e75397d1562a2fdbf9d019f7c73f4aaa23b3a355129f5f336a34b7d1e070da060784fdfe450a2bbabd520a87b77813b314ab4a35ace34cd62b86a5fcc14aa58a073f0558531f34bd98fd61b8487001f4755f9783766e664a1a1fb691df68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h553bf4410e77492181bfceadad7f705d91464885240759d770f4e7296e78a9a87ee33c2fdba1c3ba79af89770fb5fe8c44907ec2d381704ee75586e62368f997d1a65668361b35d7445421076c648952f83274faabe8eec0fe49d99ca64a527ee4d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha081141e45ad7ff447f493678de288ca97724bb1e69f821b73606a2ba26d3b353cb68e4facc476d028b1505dd0e2b457a7273de3af606425bb8b242676c0bf989c637cd9750a6a56fdfb4c1aebff11077c8d66500b42895cf21c324bcac293485e20;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10d747f6da77249d920b806fe90b3c0e0b9969ab1b390e0525d36bfd1ee0319d3988fc0f917dc26c7730c026384f49f0409eadd7c0c900394004f8c769c417a53a5a29419650ab00296174f0507ab73479cd57be2e73d635fc1b65089db26c4f390e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c0d0d024715beb15ee6e084befd013a61ba7ca532a6d25d526765702994411782d728fe66672343492a00443f05a1b10f52880165cec04c966ee439e81e82266526fde6941df4532854b2ef87055a7a9f4c1011a91c7297af1b2b4c53e8c0937ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h620bef7e8b28ae66c9fbc2dd1ed55b0c0ee1158a934777ac922ac3c617415abdafd7d497f470df2676d06206ac3539011d49760285a1cfcb63a96e88b460e01e219ea21231c181820a1d1eb22e32ee8aaa0268790324d479c727ec69d006ef6e8cfe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b8e16f86b033fad87174f5c9396b6c3881de9a11bf9cc1d25275558163e0a986628af15215578afc530eb98dcc3ab2b85b7eb87412c397eaa353c0bf1e63c1894340ecf621f0690151404da6880cf3001d26c726b978c02ae5c7086a145d795a009;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7150c0790f15214e572e3b8796bb91134ae3617782ce460aeb7c1d3c5ecc17374dfe9da143dfbe3685908f51b72e3c6914e3e51c6b88c7b31be868e08d5c74ad972d77facfa442faf3be7ecb742fca15773ed83f85f2091b4b2ba8b14428b1cca2d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbeb5b6a5e62122c5936b5242857138f2d322e9e11c15d167c54f30513942ccb1e91371e97cf87ba6b33346c49e5dcd0630f1d20ea5f74b0e4157bf9241348d57fbc906e92157fba854b647462a19f085453041f9549029aeb667480fedc46e79592b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94ef900f700847cd10d710f5f9d326e13c7feaf081648be9c50621c441bfa5d68fd1e88bc77a6a1b25f0ce6952e95930fde0013754e383693a38e0a929b52554291b7cb747efb6f40e1acc41f71b1f617234b71e817069c096431cd7febfe64ecdd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he46bfa804f7a0160b0ada246e53c4ccdfb0a1cf13aaea36c303d26f615b735556dd8a5254839331bb7ada2838cc136a2dff1aa522666a5f9361b8d6a05885fa865679816742830f0740fd2419fe446113c503deb3f4e809a9fca82f4dd10834b7ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3f120d8c537deebc531612983a7392188dfcac95f66624b71ee5b37946cc6c7087559972c2ae8fc87e76f1a61f8c86bcf63b01d5b61a810de3be67980a43b881b902332170507be3cc81bd4be624958160963446e96a783ca302c500f69c562f46a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96abd959b32318812cac636f6925dea58cfaf1d80b50ffe11116fe1df6768e43bf764099912297050d7af42e20fffb92d6971bb13f8437d11c41c25fd09a5a437d252deb1f88c35834ad8584372825187fe9c99675986216160d9a6134ee89d15103;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hceb23eca6e113de55c521dcbebb765cee2e17b416e60a383473d7a63ce930720cbf10fb592f0c6d93b9136657fc855c405f8ee10acee96bce90a33f4070de7ca0ae047ff9e6627ef4e61d0bd529a8ebc63ab1ef8ddccd6c10a6528ee007a3359bd1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1036c8483f5c59e8feaaebba70d7d97bb33b54fc71eb57c4299927d9d56e79ecc0f7126321691431f22126f879436316d72949688a9914ea41b2a4073b1b3144166212d96c356f9aa2bf1a820c389bf5de99123ce550d71c305c776e1eab312d7fd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14f7e4c960ef5735f0f2aae08b5f657806a5231129ce5fd17dc23f89adb20e523bef3dd315f4a6cf7e3daf02aae6b7be88eb1c9d6d7134e4f9097ca38386bf9e13341a3cadff3df2243c92694b302ba4edcfa80779fc51560f773b6eb067062ad1e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c272d781b77cb6b3567c1a0dad2b986d98274c7b9d44419520989b2b0d8c67e1c1ea86727179ec3bf77daf668f7b2a846dd4bf3d882d086960d1229113d568535524ababe0a46d57f9879e5e19acf53c222c26d9798c2f9ceaf52a5a155681e8fe3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h997c5f114e08237354577c7d840678ee8861e152770a6f54e71e52c4b530c325a9406f280af9b9deb7c01a0497cbb3d8d087ed07b32f9fee1c577183339fd31c2d8e88166c88cf97317d56b4833fddd781d5930b659f287d25ba0a60f9af45d22d50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60edfa69b4602cf98a6bd7ef9547e879041cdae2463bb744146c292bba77c69fbc2993cef16d7b63cd66ed67b3c539657ca0e1bbf374df5215379604e78f34a3ea37adfc6e39019f46339d72332e35617b1d3fcd72913bd3953c6fe61933b17bf2dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h766864eea964ab25b54889461f3f643b79b91b230cf7c1386e9c1d93c90db498e9d96360dbb04e3959a88ec356dcd527cc5ca14dc7fe3694cd6ef05a77db69e887d853e01faaab00fd773de71122fd80d8e0b224ca0fb6998de4f0e6ad7216a195e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fff7aff5a56be8ca2d85b77fa75705d0d79f4f8b2bb79bbdb51c9ff65ef13748708bcbdef217ac0c89c8dc0bbcdf53fa11f375a1dc426ea0563a365fe1995a00f38704ed2b1e082bb6edfa03773cf7f9b7b47ba27c5bf079e18eb5c33581c44fd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd713fed90996a00243ed6a1b24cc8eaecb2abfbc5d0f7b0fd40c91bcc3f6cd18b9fa415e8da499ccfdf1c4493aa20c968625e53dae3bdcd342684e635535bb6d0d7811aa4a574ddfe32bf78d33d994edd7b624fdb80f1b7d2ddaac9fad3803e7a78d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b52d9e25d7e4034bc35e2bfabeeee6a6e2d3498764675854882d04112c5976b97c027ac264ce9b69c6d976feae946d2f9a0b0f1194d08dc4f5c42955fa7020b2192a876431c9e92e5acc0b7c51e3fec923245dc7f77eed6482852cba86671ee3aa8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba60a3e3cab286d33bf0fbca52a3bfa521e209423c13c3ea8c57a4ac71bc94bde1b394805ac3c32f8fd2ee59cb97473a88c6644d833fa3b2c97221fba428cfa6290185bec448e769a5a2d180666009e54f2864d368f01975800f199bd4bc61a07e14;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c663973430bd890f11c24bafc69f5ef68e2d61540413e19a907b02753e1c0b28bd07b958c1bc95a807083277b12515f14d9e4e210891d0b58cc2d565ba9792ac19d451d065d98d24c76870700dcac87458e95609f3fb53f2b047123926238f2ddbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e16ab51568aeb816af62ce871cb4375eb01bdeff9ff48aca155d0293ece90e9735b1e54a81929975674e8a1cb4e885b4086e89ab20127593cefcad3ba418a67991c40a8a54e3c42264d4921d59648fe617c9711aa144123c16ec321d9a870a4bc87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41ab3d65aac3657272e02e974b01b0a0d97de00e3ad240be3650be94f08f5334b8deb3e6ab4d56c582b0d1d17695af44e1c7a913ca03350d237c7c597ad42859a65652056c033af9692009de44922adb07061f2cf32f1e42126e7eff8489d5016a87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd488756bf7dc40bc545153dd4be6cb8eefba7fe60d9bda1070ac1e43ad77d1e9e7b9c6ef9184b71e59717979a6ee51880cb4c1d9df4fe9bb152972312dbf7bc9e3e884c5cb0ee9779bed55fdcd070bd2a9de00a7a1b1ddfdc187f314928b387596f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d22786732ab190e7ff2a992fc5c0b3f96794937d3bae5dd476dc4208af7645f88f0e9be3d98956c84132d814696807414ecdca3f542d056c848b21e56b3ef4843818bec7b79c852279d87a5cc650dc5b7a135a80fa421a90fbbed8bd4e13496f1af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd247e4858a778b66d0dfc0c13c739050b7bb9fd8a84a103707e06cce9f0cb326bea10e7a19cde864062b016f3a837f19dae23d7b7cd29de67f9b46e3d516e80cde25988aa8a74d8dd35f48d4cb99b542e14b7c9b69ca834d3c70099dc402c22e34d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc468e9d7c73204918717700719eb2a703b6460e9e1ebf0382cd487d700c51d15bfcd1e6a2a4f6d849cea3404448992bc28e3e6539b302baf8e15c0256c34c92bc8401059bb1d3e2a5bcf1e376f646886ed0d7e997e1cd7a00a9b3a2d01bf9e580aea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2c862dca11dcd383ee24bcc8736f35308121f2df6012d08f954e1440264ec0551f5e5a9d1488fbc4bcd94b285289466bb820e638d45a84f581c11281e78f2fc61f462352b62604dbc5433547ab7ecc8e7c4db14efe1977b24a03203bd87ae22673f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b171589321ed65bd2c40638426693f505c72b77aaa21f50d6e972ca0c1c276acff646f8fe787a5521ac24c7ecaa37fd5fb18426cd2db17550579ec1fe6ad300fac58a10a6701bf045bec2f0b9864750075c7975075b607c6741456837fa76cae4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f46927dfb6910ad6597923ecc2c85c147beed04e0315d5a4c16b5d4cd56bf4b053e68f704a976ec77d7bc8857fd53ce87f6f88537a8f27ffc256ca8a50409f33fd8b48b80d836134a71b7c196af1b1781712545839cba3bd86e4f1cfcc10c3be3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55921fb8f0ce3cf7a86a578dca39f724194ab8913d9662df01adbb3f13dc3a47d0a3c23b744d2382ce2980c6c957cef54fd1f68a0b6482f66e84c72ec4594ac0cf9788b0435b3c60ca8367db68b47337ee26b4db51d57affd58c51a51db85b6beb2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32aacc4074353c662d0b84d696a6a12d63a2ee1c5b5e5b57dd68c3c80ce9c77f781330789b9624fdfffa46028d642a7ca098eaad1c0895177a8e3986ab34512e8aebbd43266de281e80e4546c22b0dbe3a76b014c3d6c6d2504c7a6c2995628b0c08;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7bc1a2ca532cee7448f2d811f7a680489a9085636087b75efd1b97bfc459e647ad0956465201ec7af33301c9b6afdc5a6764f136b4197749b98043f363f575abc04b3e5c499fa4d17b8a219f6f4a2eff0fb912ae108d75acff5c99033ad57950588;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96b3cdf1bf3676a4a91c68a35aab145d24ed388b3a375735dedeb8825d6a95ec65cdde303d5d4ce44bc5a0ad47ae9f82aa1c23a2094a31d264c24309c551f88007b1ba969f7f952e7bd287a3c296a19c7b2efe4572e338649bc4ef32ba592fbaafc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5eabf0790953c16899ea740e4780068a882906e80296c54dad0ab197678079e762b7563e76341033e9404ec8876df5ade5ebdcd8fdd35b9bcc66d176ad96f0fe92b40c9f99bcbcdb719c5e2535a642e4659a514ec0922dbc643cea3cb059393841a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50e2bda1eea802a782f313978736bde84fc9e226f0bb5959d273e238299ad76e2efb3227bf67b0faf9b920291c767d2076dd9ff8c8cf32c26fabb1dfa8d106ff60736a7330ca62bd7fc23ce59c912843717c73137002fc8acead752c60f6d856f2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h861e95634ebfc5a654b06e0c42d969055d1f8e775def878b7d89dd57f1bf75f2361170e718bd5e94052f834971faa2898cfa849db44422f8802cb681d6d05f1de0a7e773689ee4f7c2e1d3b8e0158967d686a0d03e4cce68f9ced44c7a642cbc6dc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde9e6e334af42f265e24860c7a0e25db5dabba069b8630b963f5dc2aca48a37f3bd01ad444ae1ebcdad2c02116b615756ef53f98e3ad2ad37017064c1046a9569d59d91e0d66e8923fc4da296ac02e446e7f23499eddd463cb1d2667dfb864b089a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34f959f8d0c3e328053867748e911e8e51a5c32d8643673bb18c63f21863d9e289f78ca89edbc168d6d3a4be5dd06f926420f55a233036a6e5a0fe5afd62f59524e5d282721e9253cc302a24fefd5efb900e350df43fddeb516a5e5991c32974a581;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecab3dd79054bfaa6b99ad98a6a8223e2637a612ff665046476903f2e9510997bb9fa6030a006d117540e9b7c42d64892a181ad6d3f7a89b7af1395e8bc4bbb25ec54cafe58357db5beb67c2b9b1523584e900e76c0d06eaca879a4e36be934b3d2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h937daad6cb5a4c4b68d3f6f732cd5a8e7b3fc7743d8a9ec4ce6bc50300250fd51f86ec986987274865a74c4a75cc036b4d5afdfb2037b88f015f6dc8bcf0551bd2760b9a78f99ef7ecef700624dabea454e9ee499b744a2202cae1ec0ec67b9835ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70d00d1d84f3254e6cfead99de53743b81107ec40129fbdec4443ad556aa67f7d6234f55d4f3a4ddee40fb34a3773bd9fc19a2945bee5700f9f553367d5f44b820d7310c4f1ea5dd82fac7da5830d6961f95ccb3d51190456b8c5f529f7cde5ff8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd49804533a2cc29eccbd4d6b287e76237932253a27246ebf115880569c57adf0bdfb6c1a6567d5cc933024a25e9aa2fa7646a6a3b7af210a5686738eac1bf279b4ed5f69f9bab9ac537da64b4c91cad5c2db19a97e50659ad89f319b338c1b7fb9b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12e9d5d784f33f9b8d0291e69e0e290e9799896f5f1fe22b91215e9c56762c9edd9f58705268e3160a492002bfbd0b2edf59f4318ff27a7c921740431863c16a1d755fccbd7f9971e405a92a7c205ef98069e465d4f7a12e5dfd5200b3e0ba814b43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h933e9ae9c5e55ec03d61b9aa9d2e4867c829d01184ab714a2cc3be580e4829bc9d9e24ce493e0a893fa0868b468b24ec17fcd191bbc91fbfc45297e2957011d06b5892c09309bf508b1b7b0f59cc641200a17916e213b480ca9be884c61a5cfbac70;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87dca9ff09b48bec98b599af58545f7ee4fc57dc98be7cafeba2d8ae64f46fd2f08d717ce45c0eadc1418bbf114a9bcd235735046034d23de6db290739aef8647f21e7b4d12dd42ea78937feb6e1cbe87a783602949e8ad9fd152c687f20dffa1e96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27924f7dc823714c97877e5476483db8d4924e34f6acc32f564e9589a4b0cae6e16723de887fe0bfa28bfab4c2127ee517bd20b181399f85a019ff45c93583aaa03259ea54037819be460f04375a9c075bc373d74e42c840605ae7516594456b273e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f47aadd525be835186df6900263374a4263818b8a6a692714bb7c3b7dbf65e1bd00ff03a35798be88365616b86d60de446f0b508865b3724cda9ab9a31ba49d3c6046cae269c4389854a0cb10e65dd9f470484619c442d3da4b7bc23c369cd1e405;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc6627cdc453ff6eed010c720a34ed4e99c2375bcd8434c5e81f351a793e0dc33d0dcdeb4fd5b4bcde6900c1aebca66aaf60018b9b9b4b17d5febcbd315463c18a0687a315b032922f0fe19601d136afebcc5cf7a042d773eda70d7d7cc4bc138217;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ac6f9131ac28ea59d5e1d2c320b408e799074ed989c68b6b4bdb8a1445e3e8b9830d23c130b59b626cd087162dceb65ca9f82fca1b2550e342b83ed378c7154aed912d88e56c1288b26afbf821f1799c7c36b3251f2151f0abe25c8382bda067102;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e76b69da2b46aace2839ba0de27cee86e5730ff10fc81a25a92045515774c303406cb3b0c593b615dfba802706662c08243f774aeeec12f83c6c2d763cd4635a009a193e36e352470e6caa9b3b4922c1b3783bfb33ac92e018daf3c100e9d75b075;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd9db76daf1a888cbf9416e776e96f450d8861fc94462a7c6992c64d42660b397ebe8d86a8e7f45d7ece678cdb6f13a3d85c0b114b25fbd3b2c53d0f21aa71f78db995deef26ff1edeca0c01cfddcff914913bf76bc268be645c5073a97a38befaed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde1c83b2017f117585df4db85a0770449369f8628e19c0c73d36241d28793a01135f85374817f3b06ab736ba488cea3649dc4453ef6a2ecaccc7e189faca0da64806a369c281d47f3a484b13a818c2f6ddbebc564192d8c07d7959ffcb5cf81c0bb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92b1a1df1f12f72bb006b8c968096d40730e0efccc6a2b36589a3ee6309701b1388022757e80d623d06fb2920557b0dfb0bd869291ccf4f5ee56556381bbee8d2779f22270ad016740efabb00c51fbb8a9b61b4252abb220d55f263a8a69217ea389;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3faed2b7b6474fa5e4b3f0f6eba0078f5d8604063420837d59ceb6bb85455ab3bc46c71dbc6f4cc933c44fa02428ba93191e4b02f4d8e1d62a0d51d43dac876798eabe1f9553417866011e16816a62256b49bf303e8f9dd8695def00d4643f189ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39c539cca5a1628a2bbddca4089927d0da2234e1dbcba09efef85c8f7d3faba7140e7de79b59f938c14252b58446703cc8e4a647f2790244519f8a403d71b5160f57119f4ad7377abbf4b50d66e9204e977d497f441ef5a0f139faeec4be78c0d89b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha675092a552c4ac6234e1649f3a6ffce9dcefd2378df9ae331f8564562250e9bc5c5912642d1f172191c58280b18246e8c817705e59c0eee6a9104ad3a54b941f914060cd8d8e6e39449f50fe89180f830a3313cefeebc1c911d2130f85e47f58112;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c6bec6c2fe951c2567ce547752e1350e473e3e0c23e7ae150a9824daf6bf10bbf3d8a3d53164d1d07a6742fc26500fe19791641c1d7412648af5b91d612d52825ead7afbc769ecf652823547e9df945c4310a8d0264efcbb6ac980c8ce71d1805ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h359b7fd50cb0615cf16df0ddb842a9448c4e87dd2274664bbb9c72b515838cddd9d2f7cc09519fb4e2ecaa076f936b92ea26b3a49728ee9c4f9af12b72999a54f5a5d984b3ff136df18e7892568bdad273098a14c808fb36da33314e0aa3de87ef75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd354a79cfc661d736d37cc4e347ca0b0513701b9bee0e7c54c82912f7a97ee17897b4074ce579a126da5c3c8ec6abfd21d1b046a8ceb865ac5b14535b13eae5c83df66c1e32f7c9badf863f1a18d6dbe797c43033884e34cca86c7e045a67072608e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca8baf05991628100ba38e9f3f7d59de865df5be8154fc0f2426a0d677919a1f819a094b2006f8612b288ffdf944349b1c475c329dc16088fd4359cdd24f9bd2bb1cba61d3805fd3ba083985f90d1473382bf2dbf59235b7e34ca304f5ac3e29264a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4f95ce2b6770ee98a42f1ab6f918e7e7878c355d5be4eccc4817b659bec87bdfeab3a822f1d89be7b40bd4e5e863b6f6b4dfedbd45b519628f328819881d0c065ebd56520bc6241b1d8c6e49678fd443dc38120c8550ff4429adf4b5e2395809d77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc595dbef33f919073b4c413ba9439ba221fe7e231c6873e62d9a8696589375ba6ec68d1136cab6d2fc318bf636be5dc7e76ccb2834fc9e4b12a311f336348eb1d1cac6d9e53ad986d56de7efc44f853a7be0bdcc285fa0c1f98747bbdcdd9cc59cbb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h293fc4fb96b768bd722fd54d5bccac702e3e4d61dcc6a5bfac1bc3cc7f908f0374e35e3a045681a8da71d94223526735114284578bc97023fbb1632d6e1ec10865bf30f33de933b797ade7eb6c0671b61acba2a62441089bd933d6b30c5d33ac1dad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a953296a5c530c2b4302fe2e5f77a76ad446d470682297f2a9192c89e0e438c7367b19907603b9b2f63e4d41a70cec676b444619b4a19dfe34ce0b9208c47f66f69835af048885dee954aeccbd96caf5724af6c55259143423e554ec3283613c4f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78eeb0d8fe9e02566008993243450dc9b68e9d2b64c4f8fb698b566c7f63b1719a15d9970e85389484e7db1c2a8de560a87ca133e6ff1208eb58eacb9eead96a8bbbc4318fd8286137e3f4f57f89831e15c6500fba0b7ffdda30ea6182c9eb1f181d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ac7e026ec0d9ee23f46db9f8eb57691d0d374ae7a6eb5a9351b541c8846c75674232771e294de8651b12a22a4069c05e28592957596d5846bd3ae4cff72491b80ab8c3f8e1e471995138e056e844e06392f558cee69e884f996189ce1d7c305e6b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c787e6ac253cd9ce90f4a0e6f0086f3ff0c84a3344a83a40179aec2b6275bed4268117092815c69b53272cafefcd7e61b772dc9e9e2de5c070026db0eadb66e4359c6243815b13d9c92674b02e9af2b6e8df4065d139152dc6022b0e4673c167ec5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha183cfac111b0bb663481787f3811c1e580665e5e770d58fbbd43fef5f276b7cd14ea428a5989024aad55a3f66c3a711a87bc1396dbb16129859dae48f5f6edf5e883c45f04a3f1eed101fdbde633644e7a859fe0e52dff5afcee0af86d2593fef2f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcffd84e2f17bbcf6c25a6e257d80f147e5df145053c2ff76639d0f447920e02f6d986b2eef0ed11b821ea92b547befa97fdd864ad6b0d71f400e3424dae5ff6fb881c758da24a77b4e7138d87701382b69ed9c10b142a4bd9fbe25e1b2ba1493caaa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38109009bd254ef3970ceb60d32b49789b9646acd8cf6c2964e58b2a2b3ca101776a6d9b5d6435611ba7d7ada0e0a7e7270d11abcc7df1b8304f576485fa51b164a062ee9669fde866fca50ddce5ef89db506ea200869ddff83679a0578f650deca2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h419d0c4314203611538aceea26cc8cb8ab292d92b57662042129fb15338693e84c03be2d57dfbd37e4712a3599bb272ac0919b816d413bf8ba5ea6924ddb2db4f3ad290ca739c20875c7a9e4c91e3a734793b7488102becb218db527f98104b9172d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha313eb2dbb550b80735c19fb31c5038a7cc16cc1764aa38a049ac8b8762e8fbefdddff00fd290f51f8d484111103e945d7da142ac48f2209ad7c48b2553a5ff2c98fce9995a4e1d5dca2ce87afbb79e8bee79f74fde9c0b648b903337c126872a2df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h315ab44b0218ce0cda887fe25e26ef8e7212346055fdb03982e2d9bf1257363d84d883a3455448d444de2bf29b39e460c6fb9166c43ab5ab9a540972b14d790ea7b2228704ab63287d15d52179b43c747e812d4d577a6c52f0f13a929ca39d2fc963;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37f30dbe3a2fe75c524c1bd803dd9c28a6643efc1b3ec63894586d16641f7840fe0b5b67c73b27b797993256ba991c75d6b69c82d00d5fd0bd488fd59ac7f23b69a2b71bf695888e8a6368682ddae208cad78f8ad1d6af69b10cc0d689e69070626b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he21fae669d824ced1e4c744cad8abc5dad7874a9a41fa62f9faaf9a6209c57323232426dd94d5df05fba1f5ebf48b028be0b5432c478fb2a5dc0911272872078fa4d250b3d1821b9b1948a2c18efae000a350103bbae93ba9fdcabe7b309c2db2f10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h998318ec9eb937472486dd5e48d4bd216e28fca05d92fa6745f96c2e5d42747d3313b06aa4f646339f5c2f005949ab0fb777c21fff7267a71a4ef38af6a1642ab293dec9a70bd9041422a12b68b614e048c477d763e42c8071800b7179d69659049e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec046cdb10fd9aa9ff42bcac0c7322ad0d447bcfbe4fce2203a14b31b85b7daafd7d979d94b31a37bb2793a32ae773328cfaa3ab0e1c7852cd86f9214dd94794fe0037f541b332a8db66ed15e76bfa97e52046657d787a7f5cee0430d5d4d3063474;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h499c17132c3cc92b183ec621fc06e6d2b92ebb997f6cdc735080faedcded87519f97562a4bc779a6a09486565868b2b28173d27eba3377301fd5b2c749164bbc605e9e38d8da7a37586965fb267b8686a5c955cbaf7fa8e6923535669b3f273460de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b1ecf2e848f13076208fa99bf5213e386ca199d48b6f93375c01e529a92156a4049c887698298fd51a98f2bc977e8788c1099f7cf4fa6e04a930f57fe8723119ffbdffd6c98edf4aadb86701f3af98e69a6a51e111c5c7926c42385cb6d783f04cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64736ea5288b232ab1b032927ccf8dab23c48d01e77bb55a669955d213588e03d9847ed0bb5c70cda9bb7589aef4b61453f585fd6f274f59a8228ea48bc98ae0728b19389c04403011903ea0aecd4912ee4ffce24c41913c154968213e8eb8e94574;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67675b3c560f287189dbc86ad2ff2ac60dcd7309f56c12e95efbb6f6d83af81dd73630d6b8bc32cab84a29be9cb39dc47bac70a62c95f592eb69cf8d60a40ba54b9a10a5535cb829c5cb43ac88add10fb92fa61c858e41c6d86c0144b83c34108ccc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfaec5bda34e974e849f543c34793b67a27588224ce100f462a0650e05d95811e66142c5bf3dfaf928f2fd88558be0a10851190b6591c2c83ae5348bf8172d1d5f8bf0ea165f15baca6515623098ac1383b81cdf0761b633fc057779f9a33711e3c27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h959e21eb69151aa9c3730557d66d33e3367922e6ffeab61f71a3284e8ef9b123a9fc72e148619b3cc40c89845b22450b751ab2425e8da3e4ca9ad68aa95a709420947bfcb040f30a8891c17d916d600bb8b1f789958ee581ba811163ac0b1079c7c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c868c2279e6918cb6b0cdd2e1a94286d1504b8ab1fd9ffe3c18434e19b23c2bd8e0ae91ac2ce923c8e986cf07a73c85fee9439800f1bcc04d71a38289d92891ba05096a52a4542bacce588de0d34e5de08b3b632f79260bc498886b8e90de23e8a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h129efcdf142baf22387b4a3d3a4511ae35073ea42a1af43e43523dcfdf1080c1ce11522b36669e38a1e9f1d71bae9bd6796669583b6f3ddd435e6ab117afddd7f4f270325359832a209246868bf153facab84ed6f490a163ef6b3d784a339441b436;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ad34abcf0562df748c431781fea05084c70a04fec76b1e155452fac95daf4a76a3054d9e0e6c2a68c7f392dd0c79c775c46d0fdc830701160de0b58bd54481b9c2cf6dbfa1f4267231e925e1ba30e262d67dbd76268d50e7feea52cfeb3296dfce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15b8aad2c3b5683d509dbbe9d3087170ef75061b96f1b87914382022f2e68a30eee6942b052ce42eb00ab689c370896daf54e03ac7c913a4a278062f79d751915770524dc1f9a17cd1309de40725a382bce20d930aedaa2e7b7611188aa8075e37b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9efb0ddaa8009963664ba00902f85a4fbee30d5c4aa62f26702472ffb845406896631f84029c794626117a4ac11a85f204d3b4fd8571c0b3ba1d28b24dd3ec2b2acf98990666f7f0467c4ea57b21f10bc1ae45d0b622f2396b0515b0cf159f8a5b80;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h529334ddd7dad18b033a53a372dedd1069c9cd758647ab5a76cbff56250a93ca9e7a5cf2df623aad67bbefeca4a124310d3197572fcb3b4c85dc951b95af43d4363efc95c4fff3c11795f2a31ebaa39a95151b4122b0a590bcb3ed07807abf19891d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec25e3dd3320f5b7c6165042f31289093baa71bc3f41ddc430b093849bcc92f24bdd259e15ac3b0d41f27b83870df7215c02b8c08918e8b4673ce1980d19de98309bd602db177841d86cead5b4f55743a7f8aebe4076555e1cffa7c3276c2afddce5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb22d0f7a0ca3bfad0d213feed544a7dd842b9232a0da9f05647e4f7eb5487aa2a1f0ce6e9d13bf8faf6f878011688f55377f0b03b2946afb253d942975f9d57c1cba3fcb3117aa10b6061985a82527914b2fe7c272d1489df5a165c1ca6ed9dcc0af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5609acc18dc8eb0f6572fb0cc2160d1dd0031a7edcb04ffc27745c2e7e00775898d778e7fd45fa47312951a5737dfb607657da562e632b97f804ec367b12eba00eeffaab60afede3dc36f88e15d4c1206a704a0197d5835a98fdc19c2657deffd709;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4150a4ca81827143b5b53972939b82c2caf3b381e2546ecb988f4cc19ea72ec72ca8b8af97745de48cf85fd7f48536dfe8b17854f0c4c3b85feeeeedfdb5cb01ca1382eade44eedfb0c89931ccaaec3f30cb69fff889b9d4214caa6f799f822a1c29;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17ba5ed2bfd601a336cb60eeb0036c753e32fc222a32a203a25b292ad4be965e8fd03a0994257ddc21ed1d3964640a1951aa1de2b21a8d15e2e5f5d8f1242fa0a01f4fd2d95f93849d43fa24ce48d7437dedf7530b5fb82b4677f67d1a8174e87d1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62e4623c168b7458ca29f5b50ed3d0447195ee23b5fbc7a0f77218a68a370f0190f7c3704880bf5d5978cdc221ee69e86e537a49a629bf755f34a718541084d828cbfc2fc3d47aa4fc0e901be930362ad0b4f646624e2fc4be6363c6bc66dc9c1e86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1609125d68861a22b67edc52abd905631863f221ad3b155fb2fb20425ae16243f2991620055597f0631a5b56f88ebead4cab3944f6fa428775c023d988dd4ae6a50e3412e3d502ad54d4ad8ea6bbe519afe71bd989bcb870db02399fd4049ffee046;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf15ebac83fab284952e67f82063c80d7e19428fbb5a8f8aeb822acdc92378c48be5b690b48330f301eca480b09193de26c616fc809142d6d915fccf7a26cbb47470c43e69b91e93b3e4d9c067dc47662d3dfda11e13e0d2e04eb1c5279bfe669a44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4c3d5c6473989ad81ef87059f53b4d1d404c6cb38344aca31792b9e1dfe0a098324046882ce0ac141cdb8c13ecda9fe1d85e148d2796dd0f09f93bf6eb506ad280b55f0c94844183c9d01fe19df3afdbbd76a4b8d00104b3ee5d399dad0188421bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3763c37908e7d4fdc0c0b1f73ffc358768e6d56526c81358b8b50cb79916c3f8a4f53cabd63b6f8877622e96b9dfa74ccc1e8b6da2bf25f0245d32594b8071bfcb6dd552bbc79eeb18626128e1a85abbe113d2d1642e8fb1988d0651ff879e796b57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha80ee3dec2b7d6792d4d58b8227474ce6b263f44b330c9779299d246b1789997f6d1b0dd5ae36c76b0e168cd68c036aa41c12f3db6651e199bbfe6007b6df38db2ccce54630b47c1d2d58d4dae3f991f968de70502e3088aad6beaea6485345fba5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50df33bf6fa639befa660176a66c79f3491ba1be5fe94267e7984794c59a653eb62d682489368e9ecab8f37274fa5a19c962b1d88b21417f9b2ad4d4242b9c87d5bb0396adfcf468c5c072050d21121950b025eff426c634a7b2c9763e1a5e34e996;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb6a0f27ccd9e23e336a4619ed6b7cfe958d49b13634784f32ba08e04ab7fe899ceefb4bd8edaad8edbb2d34f2de03f21348259eb8fb1c7cf59a8c1149258ab0fc44fb6117bc5ba50fdeba0ff05ba62ee584b6664ef85260ac0407cb9a0b7406ced5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec23cfae0e692f47c2c1931d7098ef0efd48e526a1d3654d0dc86989964cc13ff05b7242d01c00c99b6e969145c54b0b07771ad1cc06f59d5898e0a44627601147c37ccba54190f824535eb4dffa0512b8ae74a570729e3a1b28cc3fc955bb1b88f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h897381fe40f8893a4d7b8e43f3413ddf86b01dc0c21342d1e1722c6ddfef927ae5cf3320a594fb60957005112b17a7c0b38150e8ce5f9e3a8e8414eab5b5a60352f698c77ff0992155a51b416ec7f782a75e9de6c7cfb66d27fdab17f4df3a9bd6ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a4675f3ab11b9cb7d7f9d351c7a5a567205ec45b7722d5d5f6271f1c95e3bcee3086a6000c47952701a0100b6cd4e70766de710d1cfea9228a883105aa56f7dbe9c8597426c8e11aac010dc94ff37a4af87377c69b80f85a1edd150ba51d380cb6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd0feaea4f8e02ed6ca3de97467af6bfe805e9a4218a5864c944a107e201540297d86dcf2a141aa1f819a195a2a6ed1c1712db13d718bcdbac6678563696ece22b137094107ea61e1f1ffebbf037539eaee28f3b58e208d75e0c37530b08202b06f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h232ada9f718458e40a39993eab4e6bf754f29627e19963abf276220e892d83f2a02704711c8f7c37f35a01d0fb40c50815bd5a564b3417437a5b675abf4fc3ee05cb99fe9e4b4047ea40aaac7fc2c0203101ca0926eac67c8ab01b69581c7199ed3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a59432b51a512d268ab2fd50fd7363929b618bb9bb5aecec28504bbdb1eb3369cfb02870db760d90a66ba540e6924d7888239b7f5a92474d7eb2eb9a55c18e43b77f5f52d4b95954efff22002e4d7db3dce12a1e34839bbfe9850ce8c6b146d9845;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a6427230da6c24ee37f75255280fb1b19782630c4760a2e10a326e36638c75aeec571072583ae7216429cf65441f9d0a8cadfbe29331cd656f860eb3674ca34292d9a17634203d55b182d247f01e30437cd776b45d25a29abecd702eb9571315173;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bd69f454124e09919cc0f243ac7478185ad77b132d1e72c48020d219a1e47722e1848d582e32802ec6bbec1c13fb65f58633d30ffb4d20828895e96c6f8dd9b69bef5df31840ce66557b029afa6d298b984b7c54272ef5ab42614cabaec2743dc9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b4a10006d1cae5f80e8813e9505b6ef7637109e23360101a0445f65ef62f42a419098adf8890012aa5db61eaed85491f728e368d8e0a5d4a5692e37c1a62c8bfca034aaa9fc6a55f64a5f8afc10d77dba3096f653e3f0323189bcb513dc631cddb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65cdf3aaac399ce07dd7297221fc0c014ee1f47386fe3f37e1bf76c45c296f78f96fe5b68e6617e50bb37109322b8f83668da471dc9e1ce1a4bbf7199529aaa6797966304fc235793bcdc8eb2ca2dd2ccd01f11761d54332a239cb64445ab593d28c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6283a89baa166beb512d8f140ffb83e69fb4a1fd66aa5e8b5e836677ace7b8b01319ca962145ccd2b75d4585aa055e06b9fa3d370876f7d15015c58ad18ad24ff8d828ad70dab237e1ab87458fe4d16c7ae4cd68a5f02eb33ee147c7b92530c854a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h138ef25911fc4751cccb7ef22a3025fac1069319bdf5f3606f8c2516454fc12a8b0390c1ae0aeab9a1a9cb7363b8596051b0c08000de8c96c604551699d0b4c29698247477aef238357760d4a1058586a926c3f0f02c68673997883544a801eeaab2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf97d8f5968869b491b94da4c511b16d4c786d0c53d6594949d7f89fbf9a140db26e1f9766f9f78543dc75704e09c78a0585c6e2ea7bb02f5777ec451e9ad3b6ccd473843ab556ba5ac6f96f9850a8a53f0baa6e3e239838b548bd50ee20a169e5c3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h577f4bc52994e1dc23f1b2c571b722a357544e5dbfdb214ec8f7f794750359739282615af5d08fc6095d5280baf53999a3cea6c1df0cfcfa0abe66775c847ed506f02807602de27ef1298459dfdbfbfc3312e3cec1223e88a4a4150381144f5dbcf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9399b54f62f17a6780de1a1e073280cd7187fbbb491dcd85c331ee21666f6fb7f0c6daf7abd768278b0295d98d56eb4825be08904f68fba407926c607592c8554d56090ca8a5b013e028441e769593ce0760971c0a6233d4fb2a35af8d9303fbb1af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4517cb325d14f859f5923008972fdec38aa365450a129ebee25a3517f39d68ac43564280cd9cb6059641e3097cdcf1b7ae1f9e53aab203d272e501eedf6b14b7c02b698351c3fd0577654ffc8ef0483304f854ebaec434b0d92c5b80aa237f553360;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h984f961d3b9daa4adb624b3a868cb108074d1990d077c7065a0795454782dd3d3b9a82375a77e8e05a130f5ed80477df89e022108b018c8126b3ffb0d852a561ffb634377466e546eaa26a9fbb9422ae64bb50ea9b789d2217e074d8599c426a970c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e911705044d130a9380b8ab160ff6fce6a4dbf98e16638589f85393554895a51c61a96ad994bcfedfb6f9e8b94d11a2bec9cd2d8eae1717f1c59155272884937aeb1a732be746c7e9001c8f8ad9538f4a03b4f1e12311613950d2289fafc57b3521;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8bbea5332e1e79abd4ae39a50f1fe744d9bf4c78890569f76f6d43a13aeb77680d0e786276d1c9b29d9ab52eccc7316a9cc147049a5317c6ea1361b2b838271b8e6288ca54e1c1ecb0cd928e33a50c47c84600c4683e5818fd0cc63a2915b47b169;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3da7ea059acfade2015247860e9c638f1b90cf2292c838b4c94c8684a3d94f9d913cce7d43d023c9cf1b07489ab6972d1fbb5cf1e552dd8eaa3713dbc3b70fefcc6d4bf6640b7302451347c3fadc111c010a1c0468bd023ea426d803dc5457c04ae0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h126956bd44ebf397c13f4028aabdda3462cbc009acb130c463eff46adf241e8eca88d51a63f415cb59f167280c6e6fc25457482bafae3f0942cbe824e16b2e299b0d63aa3279dd67574bb0fffef9038a1f028a3bd621f4b550bc342b01c1fb876daa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6e162e81446cb0684748ca09006861d7ed3eeaad4b21ebb048116a30326f76b24530085a00db4d16be8247b978c5752325dc3edd0a09a9fa5b82142ca2ee1d6cc08b3ebbacea8c690acfec22b134b2fa7448612653489c95e9c47653f80e4197cb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82a511e9a7c078c9e5d326a9e4ef4b636d63c648cbd981ef77a7a7b3da348ae423a6321aebbacb71112339b8fc1ddd4f9179c93df09536fad00503724e125927999977195ad69b866c284854cdcb2059732769eaf33aa72c4d63112bba42d28921b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d6f856c007639c277e2eb366b7cc2b93f7a76c9821d080b4d2477f96c7e470f87b1902abcb37dd19b28f70c619245721758d1c22824a64bc24228ca56151f24a0680c912e86e3900a062ab4fe7a0a16a33314afdc3c1c056e57c300ae3c2dfc7c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e254ed28f45335ad3b83a694e95973cd9932a671da84fb34977527c7b4ac181894e8fcf5f543d7d08057c99cd7aa8d7e6b562e380b0f123504c5a330419a1e4bdf2fe4aa23f12f8df6d4d4611306e0bb37ebf5b1043e6a3c93ac8eae9e2e17f8d06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96367b2d36ff1e6dceb07a70eb9c87ec097ee80171144228ccd999a4617c832f8a3f0487bdc95b6bac06177c73b1f6e3c3ab728c02cd2e79a955752f29907642c770ee0fedac33d8a35112c72cf2b9e468c8b21180dd3a85cb579e6dd5ca91c860c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha38a1308e5851a8f4c3de44767716c9f26a6cf1f9d01020f43af7033f205141796127cf0f85125b593b1a5d74005ede84b72307320541e4c8783e4d6d14b9186e90b4420eec2ce386850cd22e7736bb601d63f8da889c5cf2e00bf2e06544951da7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeeb8701de3045c763061acd316ddbf05b94a4b5df62d97429aa4666bdff8c95c7118ea4b25ffd9eee78c45ed4e259533a2f74b0f412ad9c5cd427cda5b81a186d3acec0cd6ac3999d2855a22a2fd89737cbb1c1ece036bb547859c3e96b545a8a0e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc77284a1a9eba2b60718d8d378f40d06d76a91686e8f3c8dabc0f0eaef622029e5de6d6d60adfc623439f57890631eef684ae5b4df8400a4e51390340026162c0583c9cd706352b61d95a4fa8305a4d1043b2f596d07eb5d92e26458e717b03f5b00;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7d317e3ae37983b9e957822aad59df1249ea1e84f3026df24947f0d7aa05731ee2eaf831587f76b6d49bd7c56cd54ad028f319a957959eda1fb5dca04f22b141d57869f22684c8a64137cd70cccf0720123ef6870fa820c17c7358ccee8d68ce3e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc41eae063c09157b939c014c0098939dc70dd40ab6eecfe49f1a394d76199bed54e17f411d2ceb68fc5e0b9ac6533d141fac2f2a199c8baa8d4d3d4f7db24336803d3157c09caebdd1fb4ab22f014f6e4487121f72867280dcf32c3e7c8ca6ba5b8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfea004b71e86bb7ecd779d54dbb388ca3ba0906d898b3d60fbaf8f464e2244e3e953f1b3d89ecc26583e94195c894aa223d27a40377357fed842d541326f5d06f3f5f939cb6825a5a04b58ae495794f041eeddc7c2a753cc6092cd9c01dd8f6fd6b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51d689b5ecf9fa46b3f22c340d41ee040206e88107fef0b43da0ae59ac6d46a436b766589c38105375429dd50b51997bf3891590ebb5534f78172602f1626e15794db0f0633a36affb1b0d093509aded0a94f772613e620364eddc39a6d11742042e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h984a6a011caf0b42b8a1e7f359fa400e0a194dcc7144883667ad2f82809b6f92b4ebcc05f621b6dbf67d99dcb0bf1c7a2105218b25e2c49dd501d8fe515726c97de9c8a6d7d7f7ede7c322dafc3b735cd618385acb45dd22c6e7f9c919e077fb6a63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2caa097ee1d851bcd7d490bc80cd4683e3595fdbd4b963afdadc18199b35e8790c21514fcee045f8b20b2bdf350805e1722c7f4805792aba8c6b68579ce84593695a4739120312976ed49c9e52a5f6b1cd97214e218aed61d750abe8e2d679acd8f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a154087812cf7d68cc833d244aec257f83d391adb385e22db69665c4e9de5bfd7232bafb86d3b10f9565312b5227c8a8d56c1279b9a70005d350a18654b16f13da9014da6cd505935bf161cd79c44ad70a0272c2c82180b6ac93579c3a1169553e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h241581c7a7c3957a607eb7aa135b849a2875d932c9e440a2912f229892f655320d268350bcc44e3b6628499a3eae31e0baa98f60c189cbe6acd5e712f5a9051ed90ead7fd55c5d63f3ec5d8f86ea88660227cfc48b54250f7ff20c03dbe891af75fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58f3df53ce5c480072da0322109a562b33fb9ab2045c81b7e0a9d962d2839dcef09e89098e5fdd0a00a0113099e557630dc3d6988b55231719ef8272457dc0d6b8938a3d6744fc10720abd8873f358eeb8bb118751088dfce8583ea1b5522e44ff5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd6708e55d4f53b48331e882776e947e9d20616035e2f1e6e07dbebb6d1baf26e889c68030431192aafabad8a057941c65f5fd3d7752f61f7f4f28fa64241e3dd68b870044b62de40e27d13160f91d3f1e4c0a92f5713ad7ca5cafe822f719807d4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea5af8e93409183144f23f798957d414a9a10b58683e48553006c63bb8ecc97d9846bb2250704c4294619895fa0c80446f7839a3e8674c2b13f325bc71f46530790b9ec2b30268970ea9b09a89ad704e5ff3b01882ec078789c27d2c0a1ccc62839c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc23ec953a6b7dc19ad6d5185125fd08a24e7bcd003c9756e1b0910aba2961401d9678aaf265f87e4fa4e1c98603788c38d22e068d143abe46dd4542beb36d9a6bb7b7bc5bab6b735ddf50530785c7307974723e121691c5bf7f8221d4a01312f9fc3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd89afa4a4147479900f192d5aba9736487f2b5865f9be5ac1a5668cff5437f8ae67eea9f96dbd2e9af946c99e7f97b07a5231f2f76c8499b64d80fabc3d97c7c6182f0edc7146a8d6aa1fe3f01c85dcee56848ceabb70af53e771713febd2099443b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c71f8a8c2db2654bd6af972c98d8c38379e2e5153e0242f4dcfe415a5e421239b6d1bf2ed85378341f004592908f4f48c152d8d45251a78fd986c2db1e46eb06c979cd392727eda103af04cee221101a21bd42c424414b817902ea416f3e4298e37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8865cbf461bd3c9101341e6be3bd4c86dcd55a8b9b0a4c484c578240044134ff876cb08f390cb638d303bada6c440aa8ae403df941ed8dd9887bfb0a6cc925e56d06f3a7cd73e1c4e5ac32b59bbe94059de26e26ed6f1a56b78269d1d4f2be12a1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b41253080cb0ee0fbc2ba20f27b0d5b8f94cd40cc2556154e2bb48d8fccb7c526c0cfe1efc57b752ee26edd97079d0a1650cd4f2ecfd3396f437bbce27e79260ef7e33af8a57ef843965604e4c45fa1faf43c7f207581a61393a54e7e0d84add524;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78ec9b1898ca7ff8eaf19e573a2b9e3e7bee051c31ffc4222ff5cf1598cd273b470e4f22978a42d937d746e6c99ce4190400d256e157fac9fdccca4166e3719f0a1c29bef99f3836a7de2c4de8c69ace788b7fee28f2dd9c4c11e4deca80564403c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9ee705cdf801e37939aa70aa497ccaaf05d9b58e80a323de5de875d84ceba5d71b28c14f5df8dec89520a3806dd2ea5102ab83d15a229df81e0e53098c79f3d057525899e1dffaaac908fc35cff659aa42bd7b231482d28e67d46557caca7f9d78b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h441178b73af7cb87db3b0fed6b184236fb0b383b351437848a2473f316a8922dc48831d6d175f3157790c413e3d8484ab633bb694f5905b7e55e4b1a91b2ccbfc416509e335359a76f76de96ea0bf141ebb28bcf33b5db5fe73a874c3116db41b972;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9beff6aee54d3c166cd35330a4d2aba5a9309c66ec92dbf644e5f1820830062b2d00d64a49ba301e8a22cab2fafd6c43c7af2627ac36a13a9ff2b3afc2b02b83fbfed2ceacdcfa94a494493c69a57b299053b91905a3f81ef29752cd4fa416a743e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86b3bf31aa4930e11459177d6b4fd98270ac663f15e4a4b95dc18b3f08f20710ffaab95acc0d8dbdefaed5a28ad64ab6847fab593ce49ea93f8f187bd766ff8f2c15d1e819faa4fd1e9c5fc9169f99e9737a1bde6cb363e12465ea54d7f37a2b8222;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h365f06a2bad68f5646dd8186a08afa9dd138b532eb69ae9bfc536242d876e251973251e2a1b5823827db1c7db013f48edb8bfb4ab9272acf2dc0c84504ba41cfb7c8e07477a54f897013467ee4c37f66cd3f1725fcd8e650b93c6c82453a5ff777de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79d8cc06a432a2a69dad5a06175eb2774a7b7cb5944b2837fe37f1ca23e1a17d1d35755c4365f5b174075646e4a3b4ae677bbf07228d5369e31c8423b211f1c5e5d1fab56c0a2c9002c90cbc3d9bbc4617ef1112ca5633442b65e8a1b2739bba596d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1eeff66036d06022a56938f5674ee7f6dfe3eae1956c133aa7e96a4009804d84e4845e9704202a34376f7d2af39a7557bde491742ec4d4799ecd403848428e4b333d38856b52d666421e4a1da4b2b936947e429d68e47333c67ea2b1cdd2c561198;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf93b1d937927f392610d23e3967b02e7843f6d1d8e6ca9353c136b35121b5d49b832f14bb4cdbcef17506b4a04b8f805ffb57f5cb602fd4dc9f202b5506540912daa5830f23f6d953e0e8844d394eda159c75f897949ef27b3ec03d4a1fb01d30bd3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h676ecc46b6d57d64cd432e8aea468c96b3790034c59319000b88cd4e312b214180d1bf6aaf7ea211aaaf4fa43d58d330a90a3130b5da62f2cf44dc73cfef6ebed4cae0de5ffc38fcff3779bf7133647f2d5f6a04a8e6d100d6b59c813916be5312cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4feb2dead0d2bf4da995f79d2b77786a2d56b3fd5290fca5c1a140cb3e958d1ae284e5495322727adbd3c47b35b804d5fd96498a7f698fe9cd93203aa2f059418f02c2419d79265224a57aabf0b3b299360455b1779ace2c8885852589a7cc5f6ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e2028f02a5971b45a80c9165269aabe6289fa1135d344b2b4d2c1773c0f95e8c32a5a7a535d3647ae270263f5afda16afc61bbd06eec85fc84ffbfb4d229d6d7ff988e3be4ebaaa56ab211947f58fe59edad2f4738f92093146b77ffdcdabb747bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf96aee22c4677a4fd96d9ae28f9c12c720e03ae01cc8c8c3120be657ab8a4c39d24abb7f1278d97a00e6a7611fb7e8768404b98472874280762adb8a9315ca6b6117a82efc700db4a169fc1f806bdbf3d840645a25edbb012e765c6ad938b047a64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda91c650d763410378e000c0400abbc5d85ac41ed20b995a5ab7c9775523080a8215a2d3564f3a90e15668a7aaeb59268ac7a5fdce98dada40718045f842f9d5233ac3dc73ac7ddbb64046413a3395ff1c8e4ebd300a3d5a7fb594758a26e82d1e15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89d46dddb04e464a3edd38e47dc2aca427dbfb87f35cb28bdb156eb88b199928cab4df1175f61a62936c77a5b2887a9b463b4d7b94f133b0176d7f6947a910331898a357147d0f693295021fc5e6d95b24bf1dc718c4bbc43c9b7c4f6bf367a55010;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb09c08a5e67d6d520c87d45f08e131384824c7e2d23d5603276f64f2d6e16dc04999634cef909c244fbf9e68bad39c64418a884b65ed39c2f384a0bb381f4b989e560e90d1c08d56ef667978b8e2fe1654ca063b7d5adb8e2b9b4f4913052bf1db9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3405cfb6317c88da107a44085c8801dd0996102b668fceb67eebc1c8bc734036bffea68b1acace9433a73e28ebf4c51333384b692b7e3790893cd5d879f8a1f877a2595be3b05946e9e3e6f83bafb76226159af207f782ef1980bd126b0990182175;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h390d103027f4bc4d5c57c44d7fe7ced231440a6a2931d184f08d71386d61e610a024fe8c0a477fe2d2653e5b654b1d32990cdff11f69948823f511de0da9f51aa21725c6d8390c1ce6b1b3375202342cf79a1014945d916501818a06fec6c140f753;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bb6917b36f293862000c63003c0bd0ce68fdd8c6893d408f1579db3ad56aec5ebbc8ef046bc49e10a61bf27e9851a806faa6ac27e7ceb5a311e707fe47819f887788194ea01b09332666510cc4daac637244376f50724ee595a4a5935f199d5aa06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89409b13478452853cbe0c743ca761b6e51021ff930dcaf15f0007385d43cf4c645eef561516a59382892be6c0c39d5996ed0e5776f944842570c29bbcb48db5103f933d6464da4bc4207b3b38881e91a7a4ebbde9f7eb741c29e82e49141d55386e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37fbca2ebedbb57c16c01e750195b1a4129f8989cf31d783d0fe69e7a046879b3c8054bcedab70be78217e90fe71c70c476a8273f1407446109d9ab826da92ebdcf1744f91b61b2b218eebd8c24d059de7e4a2b12814493a86ea8ae0f4fc2838884e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b4d7c98712a2fa7a9d6965a90144b7e1a7f7cefa437e31393ee1bb018fa1832c934611008ebed25b07069354f4055d810033661b49ea0617634d680711ce4d1dcb1b6856ed60842d5aa3d432a8e8c02e45a353bfd5e299a130e9ca0831f7295fac8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab49baa23c63b2d994ce2374b2032546cbbdf2f27050136079397acde984e318928d9e64689eec78bb5343ef619bd64ebab79be28ad56238ea224cea83f44a0bed023d80768e6bcb8f9778e119fd82f248a8e999cb8b61b07a0abfa03effacd0093;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h436cb352e335236a2df6e38c9067d741aaf572afdf8fb935ba98351fdbcc3da2fec3fde738055a20a04ef4199c1108271d09338faade297d1adde52b733bf0b042c6ea43267d038da1e9ce60b13abf0937b6a1c155629dce7f16f49ea3d55b5467ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf829a40ac6d48e16bf29e7f87f58ec2aaf5368ef5ac9a0bd402edda00b2813b794fc7174e230847f0561b00e30941130435dd825f79b81a1c0cd8492925aae89a7e6ac01575da48e7e25b4e01707e0eafba1610877d55c37c1cedd5431c84104968d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67964669a68ae1666f117ece9e7578ea480afd7e35144dbf34f0b27faacc4526c35c1d89a32cc9df0f2179af622e13ea3e8c87508e50d386b0ed4dacc0904f46ac5ca3b595e6d83b7bc7c43f52aa3bdf7334ccd0aac975a2db552782d7a7a446892c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb4ec91b9913d68574fe827818d1ea6dd163074f6b5170e317c9ac8d3b0a0b9ce28d4f639e24e470e1000302a124c2ab03c3d8f0908fcbd536afe16555da69d74a7319fc033c3358aed85853e4b20066d7a50928ea6949060944c40c9f39a012e2bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb06c53cfb4b52e06ae5b26d5e8f7fac556034f6d91044331dff74c760d9359acea0821588b8ea43c5805fd5046b3ae32c5d0a0e20fc77a1be2210193ddc59ea06a3e1086f809329ea28319494c7bff9e1d874503769e8deca133c8cbd6f513d6a759;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb00f7b87c81b6dfca3e646d0d79852465d2bb579bd90516e3940fb4389aebf373b61b9583c48e265f9e9034a675bcf7723de694a3f9cdbb4d4391e5b3be0bdc62d5e0c7053306b458d023fadf18a753c833a13febf45ec4e1e8cb62b58a04da83fe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8545ce480355c024594b6ebca1d7b9149e09ff35c9ed9e80f35fde3d6e192666805704235ca58c64e4b9b9ee6bd225e391c382011cf7da2c20b139d2535a53708a7d4a47ae2e03b3cdfcd11cce20c65a66c05be7d0f200488a05910c48f2c749a14;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97b26ec7aef36e9c9a7930bfb6499dbe18a1a9048e3c9603dcaa447424a26b8edab6bba4cae41bfdfd3c2c6f5b1ebbd6c67cd1807bd76fa8036f5db16c9846db6e4d023589179f63be2fa8f9b8257ec00366bec9518d2112dff82c3a3e2dd351dd5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bc8bebd265f0dc82d58603ad23d817fdb74d1f8f634edd99900bb8b6945c030c4b626d305069a637c3018e992af06833a0f085ac962e199f1daf522eedbfeb57cd7453d4f953516edfc7c3f712be66a4c3cdca9618d6c2c9083cfa7a8774466bb23;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7b05cfe9df1b2d0219d45f10dc345f0acee7b1433066fe7467ad8ae5955bcc9cd260449a79706a5257b0a7b441c2be4a3e2e81b11962f3a92ff6639ea753899de78bcae4989b9d6861ebc7c112ae3e3e1d23ebca2620b54c89a67f5cf28d34d33be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2050bc7db5e6ee05cba22ad97672445b38cae0e8de14a4cde7229f14c9a6fa435db4a07be15a5fbf6a23366cf1d6cf25c927f332f07e9edcc998a815a2b0bfefd7ad17ab08246905b8abf46773aa866fc4caf540f8d35282f3b191ff22109f162e32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2d65eff110dbdbb78c0b14a5f56c7ad7ef37f16f4cdfa9158ef8204e2e62c82cfdc5176588aeb1e8dfb0e466d6d5d1b4cad02aa5afe480bbf9308802344ef74d0ef25d19c33bc3c0a7a3bc634f428857c3955f2871b18c44d4d07c4475a12d6d6dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h125e64d3765003c2ab139169f2faf6916cf6b3061e0edfab8ec0f3bf31bb8f9df21203b66ff6b837535375eae3e28bdf934e7af9a81e0584f57c4a3ed723f957fc36e3fb25030e55357877c7e80bc75f31047d9edce43a29ad80d26d820a13a11f28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hede704f30a55081f308c328c23d4561f1008c668e1bb5a9369a4d7a46a8be95bb980faa82b5e9a51f9909965d40f49a3e2a826bb5c9808fa7aa12ffa0e3b2d9e322fa69e9429abd1db0903025952e925ba666e090a27a5e45c6e7b9d84093ded6358;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24202d466f776f63f9165df33df502d5e5eb77966d0315ae962a3beec035bb5f3fd3ee28abe60eb9288351e0a668a7e4976be0a5d25f13e650784d728c6f11ad73bed719a09d2703185d532897b3edded9104317f6a2d66ad9a4d03f57a0fd5e5037;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64ffec91bd1d9c34fa85a34e4383d85b50b16a0ededee715d190285dd2ce4f34f12de13b061d172286b678d4ea5b77c442d3c33b211558d7fc210c1b97c817bdf2eff0b916015e8a3c8cc7f74f8c61e5cade94be1e8f8b784cfe7af6611378321c1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44825bd6619f522fb4731aa06d01b09fe7d1190550cf19f826d64e0f800a07d58aaf5b903dd500b500eb660713b3042ba4a7958ca0fb274e02f06ae409a76d2ec2880a861e10bd227fe9a3a6598e5a896b62e0cb999a3d23f8cb87fbd9eee44782aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1448c1c74f13ef8106f95eddb1f17db1b464998488fa1775245e60387efa29a8eec699268810435ab6ca7507a1f148ac33611d5c2020c6b463cc6b9697061b8433ed396da8d584d7ed6ed27cd743d9dea7887287ba5f156fad6dea0fc092e5ac1301;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed0c36ea91044798369378201aec3da0d00339a587682060aefa8675fd1b4bf0ec7564c4c202f9542cc3e4ad3ccc041a54b9c5eaa73f249c7cad77da9b79c8833e40d8d9528f1e83241555c61c9d527da8c096313af20ed21a93e749a19f581d4946;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24705769c451e5ffdb73a15f7fa4bbff19e296d63fe74f492be2cc6d3d358575ae9fe148c2d898223a3eb7fccef8b07c58a139d9053374a32014ec781968370b3f445f8a6249de6c5c4c56dfb8882e0211efc6e6519083fc45c66fc7125a84b82cfc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b238832254bba69892560a417c7caa094ab4a97229d628a71f6d08bc4e7fc6158321902449aeda01daf02f3e0aeeb4f72f17ac16fd8eec68fb57f7a293aa8e2cdb4052769fbf3d181e757b6a6248d5dc068345601a84ee2d06133ebbd85d5ff545e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe138381e6914e391bc2185b61c28c9669ddbf7e8cc3d3895e56a4c0703334fe9fff9eb0f85adb717aa9f48752ddad8cb11258649655929bd8611b4fbd94b05317e2497c9a378a91bc97cc93ec75ed07383f38829eb2ea93a042eac53b7d5ac17a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fd0ed97c57709db5ee06056df6667e2c3d35f4c636a2721185f4a7a6154e6811fbe2232bef99e1f38693b042b814055a12c6a4685e097c3c663fd785fcdb76ab3e602a337aff20a5c311f5757efa2569470005213250628b17b062e19c88aaf3a33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63a2eca4e0a8a489202fdcb141dae5e4580e78289e1ee15451534d0331ba07db9464b543b6b113942a89adc8519c51fa8c76a12e2d69ffe0cee42a535176c3c7ab90b43b99569994ed631428e65f3f330c87cf5bb9d13565ec7c5e7b7d0b10e4d1f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5ab65f1b45f8de3be801da7e66d76777151ae53817a006453949a98cba28177109b5b13b927c2685563014fc499e4ba42cc5bf0ba378a3b01f5f9781c35cf43055d292ca5d1545d1f830178fb84d6a7cacc19261caf336ceb12665fdc4a3a131d8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha842170293fc74aab21674d5bf9b38228db309caf277d177840f44fc1617c573c2a674ddae17d18dff6ca010c1ca7003c794349e306fba753255d964aa11302fe2f14555c6371c9d5e530474c025ca3d732cac90f78889ce61ac07026b82da28c6ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd68d08758ef69d275de176bb448618c77e3e6fb73009329db3aee78659052df58d072e22156972e1167e8dd7edfd7367c4d5393e595144b10bb0c179ec132b2c0ef349f13ee668737e793e1d3ee5f1752a32016ae03c3a8607493ddcea1d90a9b943;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h351d18e2814cf844f8915fc5793f0324a928ab509d2a5e53f060b5f662264a6cd05e1163fd18474b9511dd13635090af29e1a010fba722f43d5cae81a20ab9481a1dfff82abb10d0e9d5753cfc6cd741197b62449ab163e285cb78de8839c6c72cd2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h669ea9fe947909706250c268fffafb71fc7626a194e7990e82ce9cf10db494b5d1b08c9155adaee086782d3171d5b3c5c8a194944ed4925b7569e0ac6b1ac6526f4e6c9163abc4c5ea2f267f1586a3b62204b53b4333788b16a6430624516da94a7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b14f6d28d7f18b3211470736da04ee6e02091b7b92b883db13cdcde342f5cfd4cc1782309eb349bb6a9a8933a2b47fae2561439a1e53788f250c9f30cc74bcc2cf21a256ea1a23c4657b658f4eb887f90e57fb86f6882ca68325d1f707e783c0528;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfda5ae0f992c73050408dee6729554cd8972a4bd597ac013c8f00140ceb90531ec4de40ab3e527cf2a025b1a0d8fa8e40d3617268213d5246f8d8ce1e62d57a4131a39cb9daaa7fdcbd096bd04638aa00b4d973b7f1a228dba14e8d8ed76b6d307e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he25fb1ccad8b0bf666f84bc44459f044a65770425e840e9f7b1339870929884bb8ccfea27fb72310b2e0af47f44335f8c130f1eef0752f7f183814910815023a623c20fbe0aec89649c0c55fa32465cf70b0d7dbbe8a0f73aa42f5ff38c75a0146fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9915e343b92e7469212843b373bc4d9b7c209312bfaea946e858aa50417916b086ad7bdddb16dc30bf7c318633bd858c546b7f62cb1774e2e22e0352c2db98aa9300af1fd1095423e80da8e73ee10c38fb403f3bd0458c5e886681bdbad793243e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfff1c5cbb042ee77365d8c2c38746a6b7203e79c34f927d3159e3431e8f2096b774b019bdc76b007bf9d44eab2b35149ca0ea2e3e5e5e4b50d69dcd60d87241d9829bf4feb55efa1558dbe6436b932e056253ace372e4a6bed46bf89d40037bf24c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heef0c4e27796fb0eeb762825e4af712684fefd5b2abd6f8d157f651e83df00b5af7acc56d4f992d9ead3019709c20ab4d3c9cbc25d5edcca8aed26c54602b83c92a428e53d157726c253d6a23d1c5d4e799178ffae2485704e0c56bd350b65d5c112;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6ec6692c054ba56d77dbd6d56a744d569448b23c3ae50eaf05369e11b8ac2d21be74114bfcb887bbf69f3b688700927a71125b5d6209df32e6e1d7f4e7538bbc4109485ee8695984b8392a540a546f6830c3fc97038df113338d50c9cf07b4c84cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63653e9c51157ec67baf437794efb8e2a5ed2c46fca5b6075803dde7135ea4516594da887f5b735bdb87d2ee8f5d88c7abd7fa2c799853d4e8140c523a7b5a7ec04a87b6682ebcd9e609c45e8cd112e2d2a564e6a18fd65b3aa760b2ad32b540b364;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d4d405727d8b40cbf5421a34928815b0607b42f4708fea3167c47b745a3235668fa673eec7c038e066058ea9a99cb44f5dd09ea5352a7b2968f2ac72edb989f90c71366cc0d7b9d4b97fde10f43ce697a8e0db42c0f1bf10558d5c6b2fdc0414058;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fcf37028bf7d7bfeb0ed2cd0ba4e55d19c14320004ca66c06d68d6d5bf81352bb5bff97da1487dde4ecbb31f68cf9f18178b089b1f9fde07d1bf2659f8d3b72a5b86dc8345f67d1b874f44c4021a451621101cca57f6974d85cd651721cf08be774;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9bf2251af9e780e850e6120cf7eb1c3ae5af459b8a61e886c1fcc771354d5984b550ce4476c485a5e9e2ce5ee5428361c976b34032022a4094a292a696ed9c08b732d4848fb8d1958231c3b9486470b2ed1309225e94374bb25440d52e4ae3b4516;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7634c600fdd5b379d065a166b750f2d6a8504685471af2ee2a655450944dcf65df248967fdc3df995a15c182404fa99f0339ebb037671761609f275bba8c4ccc8db02f78e2db00a0731b32b4a35429a5508bf04da88e8eb9cbc36d2f56940204a923;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fbc93fc9d7430f2d5feb0ad2b84bc96bdaa8a9f6582a810cd45c6a8a94ebe5888fba0064096c3040614b4a0b76401ff2e2cdbbcf38f4546569985da891bf98af26d5e1ec1b81d629792f20bf463077d85580178c16bf9b0fbf2c087537cacb9c6a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3531ffe61aea72ae692c3c333b8c8d95eefe4bb17912c9ae9b919e1d6d53d18861e7a03fc4a1c9030a42849acb0a2f4f4719caf67a9238de8bb6c38544c471d26972422cb0218f39a47e0f104468d8e49d92ebf8c27730afb41e14460237b5e47b53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf820d121fd2eef5e089cc11ebd2f87b9d13fcef19ec1b6227ac2a33887555820a3039b4d6e56947f9f2df47073f661f113511f62d8426707a371b694c83d1553b78d9a53c83b2332a9c0295bc6077944df3c1fcd84cc306832b18784429fac07cdc5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h135f5aee38fa0bcd25d0f963eb9716b992ab55370637799e743edff567a2bd6f7209bed46a5a6bb358591596f38c8cd745f9c550d1e2b3b41831359abf5ecd8e0c4e91ce668e61532a2a1a9280c3bab2d507f3d75f07eaa80fae50f6a5fde1a62084;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97ee566277c20497d1bae6c85cc6a58f3a9c6847e85be7142b4230802ae1fbcb7111e63a2237fea48cef6f86228c9df61ef02be2cd1cbc4b4970369d604de434dacfc7ae1c02598c5ba8f3a1ebea973161008076eb6dd169ec73352f812e54644088;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1707fbc2177c7a49894d636880860149ef2f23e87a382d3c08e2825ebbfbdaadf2ce8fc88accdd18c7902bbe973605ac494d3ca8e64776429acf3aa4ca39a054784c63e11cbcd79cfe50d4bf9378500e49052c7c4c932677a0c8f89a10cf3cc73d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ca035648f16b0aa576debb6ea7cb5d05e750921434a043aaa9e29da310a14a755a9bc350b8e56a81b0b3f57a87c61ad78e697d0d3787a40e165203cdf408c9778acc6a39c546249cf7261ce79c9b974145b943d8bad02dc1c8cda6ea5906c4d4b1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bef7b764c6e92366f824a170226f6bfb530d1357fc2ce917e5c577a46eb25cf44cee0b47517f5420895bcbd626c62bdbb9b44a1522a59a9417d2703d93d58ab426492ff12e6328f5c6b6669db00ac34421f6c9550cfed7a6dfd0546a3c86bc064d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9551d272381f7ee23471cf5a7552d480e46e50e774a90580e63b5b84cbcde863791cad6a16a18932f9c1c699e66e9ba797db5030669917462b47320eba70eec30f12e4f63ae277dca715b0dc266ad8bf8ed0109ec4ba2b8bbf32953e7c81a6a24160;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cca196475cfdecad9a011fcf30bb83f90cc245907675c1e100fb1b779d6e32829bb0b5243524c25349128fb5087493e27efb2e8f2b35735f9eaf5f3a4d0013922af30225102b82353dd0614a26ba12c1b71ac7e92e22d06793915f0e6ce79a394e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h535f3e775c2c7fa55a384cdf6e3781db47a061a920bb2d492d97e138b0e2d5c8acd363d61c782510dd77db74c019ad83c04ff29143a141789966c8240fe1545d25b707e547e742081af6673753f1397989088119ba43f9e5b0394bbde8d6fa9d42f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7ab34054edc350e43f64bd4fa9b7d3c5eb1355684b81a6dee8c65d5b8b614eb7d56e5e8897f0c111291da60b6fdf451d3c4ab0bafad34502bbc681c333ebaa8bf922af68aa2da192a0b607d38e2a9f7f006c6aa25e49b8823f476d962a52d3997d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55a0f4021e0676ca0790b51a16da21019966e529b48492b1407afad533a763c3ca7c6c4c09a6a49400fb399487dc6cc64e65184cdd1129026886d6e62926a92eca8f30ce2a21718f1fb3bc27d2498a6f45a602a0f1cb5272d4ccf143b9ff2c0994c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3e554cf30115b66119eaea69b2d5892e0e4bfc7719119a4493902413e0a15068451cf83527457e2e95aa4d02bbc93302db178a6ead21c2994e2dfa1f3ced9682c8ec0dc07ccc502f532ae376ef1d5ce161429e8ec7ddc98b95c838402712416ebd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e6be1525111645674b1ed34e10bddf67346c0f8df662439872fa01d8adeed1c81129cbbdde47b48e5eec66ee6ddb136cec2e1735f5cfaeaec13db2e12f19977dd58be083625f8630ae764d76dd4c3deead99fc653c613a25b4b23febfc18b3246cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dca2273be9ea4db40cd88fa68ed295474fecbef18abf9e1fa6ac84440ed30bdeeb604ddac915e6bc9fc29bdaacef16f035d59ae2abbee4e05d766b772e48aa62964db2a29438e45968a853b1a3acf65307172d0f517746970024b52790ca88467be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf42c14f6bff8d8fab69775b60fcd427bc50913b93af49e914c96008365bc0771140f1fcb6e6ecd19151a160678f753977ab40b669448c7e9e5d1bbe3a0f91ed5953c60b02b723a2bbfd2a4a600c2f5968eabae30016542fcce15f4c4302254e34bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7935407f90c1525259617e0214074c4f3a0e0b37d7f011d825e9470772b80c74805cbd61ac3205ae09a11349225f5d5d6b3dc8d8e55a934b8e56a67b6ab8f92bac59ed498f280c818f3ca28e845cd64fedad59060d2799f6d682fa6d440953d0408;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5d3c9d36316afbba22fce05d5d4e7caeb43fef08bf4ce46556b6f5289097efec02b61c819e5a61269f3e8445e74f1412eebefcd8323f6d8b5192865f979a336cd8805c0d593bfcf3f5ea16ade78025ae64f33242ee778dc331b36576671fdbb38be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb32a1dc8eff3b69eaf1a010fc1062d4bf6a4b127ad6c053d4fab0901731cd42e1b8c1a6af3dbf1aa4ea64def6f718aebf0d847b71c3060f610ee6ad8d8e10c417b4f21d954b0942dcf57f506ac1a940876e986f801edd2190ea341dae5fc6f8baa2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7bb81eb9f858e3db1517c3db46063b43470609ad40c88e42f7b0a276f5b69590493bd9c66d22aa5d66530c669c0726531e5c71d58116745ddfdf1fb13084285bbfc91111cedde16b493553dd79588c140868bca0f8827d42901e69310a92653cea4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6be6f83fa54eaf2855c56334341ca232a93af9404eeea18cf3ddf702042e115008160bd3508a1b580c1b2bf5741076d3da3fd664107de899a5f27b0f3d40718e4efa4df86fb330f4bd4494d94df37342c17030b482d22f83528989a5856e975e1035;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha686e54d556ec94749fa3571efa097a61426883f2f9b0d97d2bb62529854f78e6bf225d3a34aa8b5a9d286586ef1259de839fefa265065e97a27f33b95468f6e3a34832aed36417d1bd4b3b87e5fc0e5f83209cd8c06cbb652b9b6a3cb7bc2e50429;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24d63bfd756ad7e88058e77757cd9237e6188d8809ee458766e8037a8ae8409c6343be0b0011bed00327b36e5289bdfd745140b93bd7ccac8333cf948f94e0e9d87049814604b4207645263efe335ba68aca81f5207e2a7f90fa170d5a850855e396;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha780a7ae5a893aaeaddb35d3c731d91ea540574ef06664851b3d60531dab59ff5a449a9319430d96465a1c1149770d66dc5d61f491469b4b910ee87bc71248285d57b95363fe273453753bc0482416096d7cd4db466070a0aae782980efa16ad9d05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde583f14b5f23e109917725280bde04b30c16a150f9999b0b9bab153d2861b0f88ad3be2a900940dc0398a899a27827885dd22a8fa0967ec1845b94d3bfb70e14a847ba1d7bd6148eecf74f6f2875c38175b34ad5fcf49e10b96d0103123938d91bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd09702ac4e2e713581d38e8816dcd95a7f6941102f1ce566c3b089c96db3dd3420e5c8f37584011333381d5d87c740fb03703ef915b62e59aff1ec8f3dc5d7cd04b14b833f08cc7a44034f66fe770ada5927aa0622a85c1a9ec32f663a96e28a2d17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29f4e1dd2e3c6735b290678a84dd7f8044a574243423d9b96ea2a591a0f63b93624bc252badf912cad7f7465c912707a4fdd4362563adf2c5ea3659cf252d50f8a9514eb491658629798df3d29e0cefd011d6bef8b5160f1483bdb60a89ee156ed96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74e06addc2e174241ed89386198c54314e3b4cab5558f780885593b64f2487ae8915d3f6490a852849239e70563173bce6b62fe1d9071626cc83d981b276ef5e9fb1550c69224ffb1bdef4025b13c79751e738b9ce3696c34774fc25a11b94028066;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed9c6502b1435b684d99c3863462e60ab798242401ce9aaa182805f72535c80a8de83e9b944f94d665981f58b4797828268f928a432135d922b1ea78b73f579ded5bab9be32cfbd4c83401aa731d4a12e2e9a745e97051a388e7fad54d002673ee8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e77cf6e577e98772f9ef27c3c18130fd697aab091f3555025b549657f00eacfd2af917789bd7097b3e11536987a148279a5c08314acf01e0724ff4981e69c62c54e172e331ae4e99f2a607b3e8527766b43875d5ebe482546754174d8d232bd4973;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cfbae53db3774167b9f13ec2da5e13c9029cee3dfdeb1535bcad3ded926d24261401f92f12d3ee3beb5bbb17ead0fb2aa8976bf75ca619ada38c8fbe824033f4e444f6d8d32fc7288a070593593e11fb32321ecadd0835cac5b94c5c5f4556f7926;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e176f9fa4a9baa0855475f7a068abe2e30f43dc98cdf5cb3677bd707fe546737946c0977ab44399c976b701c8aef9bb6ce3e42b41e391c9a040331a65378e970604466b7bef39ca476df0a0fd06a2bc5c8f8b52da9c0a938d11ad5e3f00e659f61d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24e38493eba6abfccfc5b958a66f7019adde5836ee3780099da8da976c968adefffdbd8e21a53803e1acc45be3e489daa555c5fd3009ea29718501af7821b22227a22be260609a67fc78e59228617be62000c0b7c92c3d2ba8c2042f573eb6447a77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74bea97ec1b58b8f81795713e9b6903977def15a80271d702388e1be902604df423cfc0b7932d23acec2ee8cebeec70268e95c624acb402be8abb88121a93bbe26dfbbd879bb9eb977f69123a41d14bb5881b6296cf0d775dd12908181acefbae809;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habd809dbcbf78eb831a0444703e49d8b758e958131cb0fee765ded46d16c630d9c282956f07f49d6a4a195aaf061be81d209541c8ef451e68bdcabea1393438e5937c926295cd797bd48a4a6a540cb78500b0172a3dd968ed7c82cc73afb80565e3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f950be1ce7115f75e32a9223ea4f0f779f26afb44671cc4b6eb836de2547698572f2deb13a098e5efee2acb64977194ccb2179af455fe9a953aa380aafcd400deb051ad5f96288cb4ab193d10d6634fc8b951c83720b84624bd9d349deb39656975;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ccc5e1d243eeccf035867d3f0ff8b38247350ad45b9f59aa8b66a3abaccf3de6169dc5ac82e2c15061c221e6314d9582872e054ca1d6e9f1084b978b93f57f2f20d2c2675a1beaf09651f8ee4b7da27b8602e930999ef3a7dbaf452efa3c1428a54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64f7c94f7ee8caedfd461d2eb02ed88817125ad26382c0db9ed7ac82576a3bbc50ff9a775611728c0131b2a43cb29311f501b03d994e33b318f2e43ce4b6946188ab2c1268957170fccd629717f9d921a4b2d02215010b68f7f84cebfb475d838810;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8448689dd44bac3f80e15c52c98b96d9f87a2a98d5ef4163083aa5e60214e33ee5550e613a8e7eee596cf2090691f1d17143ebee872c0ca21981004b8e3c26fb8a138d7e8ef38cf1d8222ab5b614d33052dd80c8f8e4ee8b9097cc95a516d1f8e29a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2a9e2ff2ba5bc8d27cc2d81fc59f283e5178b73c509e90b10e6402249f5e6439d3399c2aaa280f675ef5480f8f7848931e81fa662aa1d0c8ba718561fa7024c00349d53e83506c7bebdfea0d9e7817ffee1f8d6ee8b7d591da4b50e29dcd55be82b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf67225bcf1c13cf8ab7855e4f80c34cd33ee35574cca7a575891924b86283c7ef5383b7cb28f2fc84b945e554ce866d3b807c52162fa97c47df1631a889225992fce0fca4585920b27016b8a5bda20455ec1afef2af115c11ae23e11d562a8d05f89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h693a3d8fe9e480aebd09a53766ccff4da4e1bb0b757a4cdefa2e24727dac0f432e1c3a701cd2b01eada90a5a242939845e2f72521df2aec69bce8866a22d660fea874bba1f8421379514b502f38c02218b4e391231df5202273c7420a6cd6390abf6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h977ff4e05c51d19e00eb51eab30819fae20ceb3d9fb6ebc7b023156aa2391920d805fc3de1c7e59c804f089e90afe8049ce96f163d067ef0bd60a39742eee8f275f87798ccf4fb967075ad440e738a39a432476669ff077ed6728d560d46b2f793f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha01e5a0f69c302eb864fa09336c6c90691480919aafa0d7f0391466824600beddbb53128297eb9e796e264dcef79b790e68a2e7b852fe8e2d1f754fdbc19fc77d1b5406c6567c3946588363b822b973ca63a973147763ad8453a83b8904d10a22c9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h975b2f47de211fa1d036e1a9399dfeb219655ca169e336c8c566ae919bc2a6230bdb5e4050e6c1cec6c36f65ee6591fecc3e7a4e06748fc9460a8ba732794cff358d32a90d66bbe86d5eeb258fa5df057c8a866458d657bc1ea0304b24ad5a983fd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfcd46d05d25ed861174e664f952d8333271001659cd0715927feeb816849b03c06de544c13f419d7be2b80cf619c33801668a01441afaad9bf6f918d6c054a5b1e6cf78f89a70da6afe96c17fc7a4f444bf6a627576387bede9fc2f2b1c706c257b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h857671e44c6c81bd8399806b4453ffc25664278f70d7f5c51c650afa3debb0ab459d32bec3ede282b2134ae6187ff74295bfeae6c68524a9786d794a842281db71a8d4f3600c19d161efd553eb35dbb4dbcd0d762ef3c9c4f722afed065c11ae343c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe2dede46958286a219f72ad93030d546e34ad1352daf6a85aed412d558a07beafced96734b128d7a3dea547d396ee9b2a1e8f4f8448a2be2c42dd6159d30ac9b739a25673d7422f89153e66f2c2836aed2cb5e1128ca52ff3aa15c007c1fb7e5fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h215766330409ffa30293d1cd3fa2a58af2117a2cb9a7b500f3ecd1ba4f61eff68848a6528910c7e136d123ca90e0c1e3528af202d225c18fd1f4fce5fbb72483a6ece3d83c58df74231fed07847181af9cc91f3ea3ff75e7df9db11b06278a07e098;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e15a748d4cf96d98bb7deab56da88774bf719897ba290aa39cfbb0d92628bbc140efedf9186b43c8ab8174e5e4f593e39618aca4ea02478356c947fe7074f4c0b3ac1195b37616429a396e242aff5046694fb4b84db7e493853bac1da3e087d8e22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e8d00573ff608d85a20ec60f31ee68f507ca408669aaac580d35008207942b4d6230bf846a95d8eb7bd95190a85fefeadd6dd9b804bd8d480ac6ef1a974198e9ef0848276162c052f3fa016c020ed22be1373f8a228a8de7ebed85966c98bdf6dd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a86523cdeb66af3be6b2bc441a606e4256b5e0916e6f436831eb2d92b7d2a489922dca8ba6aea546ba6484b785b36f53089a48d32b127a2f4310b5fb5cba3774f3169e8264f20a339ec64e43d5a5891df61647ef5648ff2bceb211b6daeb721d252;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he688aef617764a8db9c73531f064fa7868d6cc692b9369f672bb093574a0f547087a068c9a0b6165fc4eb17b7324e9dff12dc05810b7e7e0d39773dd8d66fb066a3bdc61804eb47aedb787a4d8cc2bcd6b6609d566b0e3010bb14e72b3673a0b192b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb22819086b025fe8ce80e6e22ad6029ad42455f684c3eae056d835eec0f90d53363644c67f1c6f23555f07dbbd2ebba62f87da36ff6727349e551088e02f5ef441736ad153e41c9ecc37ce4fe9cc0b71b920dc0ba114d017bb089ec454a2eeba270;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ad34d7a88328bb65f51ef3204b411d6327f4cc9be818c1ef104b0335e64b124a343d2483c273eca726b9dba40210315882647f99d23d8958dc5da752845a2bcc068a01a7d578ebdc965f420f2cf208a51e07ba9a0d43396757347f288d9373476cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a49908c78e9faec7629ce7861e9c06e2552e490358b52c25c43d5ce65509c362cbed3a66522cc9501d797767d3fac5196848989d3879be52a93b73596c199ffdbf36004a76883a22b538950e27e6a578ab3226fa317cd5ab3f2d51a1f86abff5f1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heec2e3aab2fd6bc096718d0a41c5005fc44cbb1ca0056fb49f0eea666aae111f8efa69e33843280d2b3266694754d371bcb92f46aed86bb6f254de832e15a4ef23e909f6f60114e95677822200910305fbb9f73c175786a25b470936a205213f23a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93b13b0db75b96bc74741c48938aa1ae34029bad2a3d2527fd6a35eb977417b6d51542c8e2431acd54ba683ba341d34cb4f7b668c9bf2d7cae58e4d70e80b5f16548576eda67a8494addf693b87bc00576d82db92ee88457b058d9180ca67c035641;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc16c6f18321f6e13bdbf3109575142f22a30d2a35d9ccbc64f908fe501ff8dbb579311f408ecedaa996ace7226b502197434a4e70ebdd1d4e884c6566b842235869bcf2b87acbaacc6b3014f8d9064c47aa577543f563a6c24598a01bd583a814b19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce24239ec191728125c26afb8021fcffba7f290f1867a9c358ba13f72725290c486a722ad5c5ed1db4ba39275e6b5cd20eaa74ae1a34fde6515051f0c8b9bdb772277a71775c7ba10fef607d778853828fd79130b2617eacef1491fa486f3a37d8f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75de4a305d089b8f7a359b92240dbc27779a5ecfee65fa1bd9496756d2b6fab89e8668a3629fd79a89503ffc51444fa89622cbeb35b32d87e206083c5753f03e0c3ddf0fdf6d253eb6cd612503e0103a0f6ad0d7cbb29d1d8a3b07a83dd2325af41e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83fc8659a8dac520374346c0de03cb85d49d332befd60909bac24cb8377b01b518b314d1268fae5cb2783b30d7631b5357211feb0f1e41f4515fa9f3d65d6480bf27d7fbe02dc67999f9efed1deaf7e60a37489d0f57245d2198865a2f316ecfb58a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7cc8b8f516291d4ecf44b8aff5819e5d0b04e27444ed6fbe41aee9c3068657573af42ca12e90057c05c7d0ed50683405cf64f8b065022bfac442c60b812c08a7eee230b03dff612207b1ffed2a6144a9bb0bc9368240c393bf3de155546a7f4d985;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5f8f8559b384685116621881e7ffc282954752b56ecb895efa4d3f7dc9a4046044e382deb03f5ad7c9c29d09f13799c50b4a2dc578b45e4d4b4db6b523da153fd909ca8613266d7f98a9d2c291ae49592897baa62db220eb7132aa8a10721d0fe79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h286ae84ca3b73cc9a6bd7a0e20647928d00ed0159ae5d697a1eb9e891cd9109a75216c33b6031024164f025a1034e90263814b4555e5d5f97438e0ecb70a7fcf2a349545d79c70ac8a8f6443808c835a12354908732891a83fc6ae2610325c8ceaa6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5a4cdf88de17d56c2dae3b2d555b2fbcdc5548d52abcb0ec47036cfa20c70d355717b93657d1920a5e8ebbf17df7a2b88639d98287af999294c016018d20d7532848f985c36be1edbfde8577c07116f9189f9a3251dbc83a1da7958017b95963fa9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf6ad829c619c6f182f5520e2e41c9749e090d52d0f529473db21121daa8da94719d06a2fb616c3ec648d8072566084abd02cd36e2f6941f7ff558d473745b96273d22ce2a50be6db5e0561b2d09e5d81cfb7d58378e39a344de147e3481d882604;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3528a31e1fef8079dd40af1f6690416c94bd5b8d2e84c5a45b0dd7d6a3141a93b2ff8174c241ad974463d521434488091f149c96924c3e6e969ff50a7f50bf1be447c63ce04b932d7afe21be31630887d2851cca28359ddcbf1d459dc37b1a37a99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80809fce24d62856fa1df61dc2c36e2c9115fff7fe0e6b9e65d6ea3af2fce8cc9e0ba5a1c8dfc5eb26a6d27f8bf270f782531586b08ccb6d9f59188522a3d7d1f2cdcf0e7602ce800f685f0cd3218141da447ddc97753fa0a20811266d58010f9948;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h104100efada093316e04837b1c68fd15c56eaab3d931f3e6e6ef8b1fc286637f5eec06587fd602e584c01f87d403f4e538e47f4d51bbffd9e5fdadb12ebcd741e1b78e1aefcd5d412b98e719130455af42be562f04b66fc04bdd06efa8c5c37cf493;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h873fb63406d68459dfcaeae5e63e23e5b96b1a050381709aff5e9dc3f41d99f829f505771324db5b53b7a93b505e52b5b6323d27b249a30067368c806b862e0b7df1647d9179e41e2bd70d6cba499a6cd8cddffa9786dc5d1218f2ccc46184a9969b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a45ae18552754b9e8ee2b8332bed925565bd400bc5b52d1404c42845faad19290e46dd80631c51314cd49df9b551276507236724509fa29e189e0d510d581afbaa424cf42a492f9a35902431129f920dd1deaca3bbd42c0079229290e2656464bbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c717829771167d165c0b58b0265657d0b43edb245cbabc08e87f3a89c2d909991607dab0d1f4dd1a9551452c1a8bea57b8e92dc28a407989a122de8c95c4b35fbdf3b3a503c8dc18120e3992d84b41dd9034fbc80187e505bb5d0c3888c7ebcf659;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24fa25a84cca2ac37019ecb7490d510db4698b4b54a5f056f96e1c37c1a2034f8e63a584c02295251f77d05a4714fb8bf245380c667c067a9dd504bab809440755ba45dfc9fef426eb893a7ad30ed505d07dfebb61c7e8a906bc839f0174100f7749;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h873d337e6f4b9c74b58fb9ec545e55b5fbff477c22aa9d9d9df0fedf1253fcb98872c7f0962b8c098283f7a03a811ece570a301c1bf6d9f617a477772a826efcc19898d79c2d6f617a2ea69486ab8026503693ae7e92cc5e16ca7da4ffe20e5d0610;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha749ca29695effc90a97b7a3fea8f486ef3512691cd8c059f626cc85250b058c716f8b9b886787c478fffb2fca1fe6bfcf61cbcaed6ff2b65c296019ee81a823a72b40071e2389b47d79c66854c5935ddb2ff95bcd106e0ee586f339577471763efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8cf78b55ddd2b5c88eec511309d92be6ddf011213f53f4a719c9c336c4153ddaf8aab6a671f36ab302eae89aab89beb1c4cb749040782a18d03d5db89628ede53d8da90483c3edecac0ab67f290e0b24f7ee94a6fe92fda5f158925a7d9a94c105c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebe25f54f17fa588282036c4401fb11cbf3f9c64936918174a881ffc2d7bf04a1c2decf7281ea4be68024f1bf74c736a549a19c6320a90cbf6e3b27594a53decd66e879feedb570e27fd0e270232f5d3d0e5cc86c752c95886098881724d0fbe9baa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee8751354f5e1768aa7856f938d9206c5d43d6fa453343c22ab49a07199a9f02c9aa6cdce43dd4543319ab1bfc7b003401ba79a43a2e69d8fdce57a5d8439bb5a5d0d5f40569da1e63cc8cfc80d36fe7e3083a07f4a3a5eb424db6a7ecd1ee30c93b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2416c932cf01d490f74be58411ba1ccb1d4276b14ec7701f2459193dad152a7b44168f1111559c980bd92cb62e3cb91d41f32639f11dc95d830186d8b486e46d7f2849e305c2acb68cb1cbae6f577507efd526c55e42a87edf4f6aa66bb534b0ab7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab6138495b2404164b6fef12a352020161f28359f1d4cb8708090f703a385e45317c3f32ea23b87224bf25bfd5e1339020bfdc6f2a2fb3757f1ccf0b860c8919fed921cc1452f89d8c7bc2bb681275a30e5e8e1a5ee4128f275bd09a00498625a3d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb3ddfc706ef4cd3684429b83606ee3b99cfd43108ee0165d399b81a6aec37117e54dc33c960b5450603c9d599f17fbb7e4af9cd2b0376869f87005388b3f678e616976159fcec81daa1cce27cb4d576a46a8f825a3b615633b41a6e3ccc0e45782c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e5949cf5253f0d42049dfbff9eb422f820cac41ec768d1ce22f414af299807afae009db4e15030c67767521bba6b3d1e977e631091da9b7b9ff18fd05e7bb661936399511e41af1d29399f99e8280baec586a7d030375eb7f082b211424357b85c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha73a97b1c407b6a08630634a570cfe27915092f592922d68c6e25c0695523788dcc24e1f01e9b4b0291c97ef1127ee7d04b51181f2481e8313a96f53a8acfecfd7dab55771fdeb1b9739c146506f40fbc4efe3c47612be41643b368ff30886f6c147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11ed0000f9152bc0e47f4ed29c8ff2b3464d274e91f4754f686ed43582aae4c5c7753a7b5de679e2775a7055a0bc85db301fc0f1f9578086eea5f22292c76fda61030ac9c0c8909194fecf83247a388a925a5254ea65d229d445425e8a3e27dc53b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb35df8f61aaa3876ecf723ba267f9ce9388bf38ba234b8911b08865d4f87f7cef2f504c5dc982abd853cb1b737b264f19add4b6ce1cf5f5f0beb5a930f9d76d2b48c07b22b8f104a9a3df8e47cb57dbf20348d375214fc2ad78e7e6529c78e4daaa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32b65736b9f2f01653a58703208f3378852cfe6ef03c04617eb23a87089479ef7b234e228ea51bb5a19510b8782932387f5614afffbbfd9db5628663ca398646a337aaa1cfce10d872401a696801fcdc0caecf16d59b8512581d8e6a3c8dcc4c7fbe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1f1d56fe01676279b6acc52f57036529d20b60f350f59f865297b39f3a7e61b7d0d067742e3997b3f79701c68dbe0b10c7f75ce3a9bc49b5396a9d3e9b7162acf5347b5c0fe6d209e4b8c96503bc8a96f789b8eec4481907e23b231a48c22cb729c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9178885daf675879185406c5d15e145145b530284d7c7d235355553b98feb4aedb6e3eba3ef872a3fb674ebafc3df2366f2f963aac995d3379c814de2086595e5245cda6fcf5cd9441b8a1230651e078831f1dcba6d997d72d3903c44007afa458e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he22e0ea9b3ac51cb75dd3865ef492acae7a745706cfc228cae08d6f753b3e5aec201008474592460decd00c5de47f232db2401a437ede48ec4883c9c77bbcf96545bcdaeed8ebebb51b226977628bbd17ea1a1167577a969b17c638b0fe7041cffd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcef6d5e2c064a33e455e8005b3e204344d71c4b557f3ca6daa01049159884107fadba21472c7bf141b3d31fa3ff1ed4e2f10b571f848b2aa8660b4c97263be7fb94fe641108e0ee725914b076ae5000b87516b564f3c14d9167e29ed8a1372faa023;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f8aaffedc83cfd32964c4369c5e6c4f83f902c9fbd0603f2d658c8e47f5eaf93af777bd51e736a72452ac7bb3bc60150ead53f87967dc2b4df4d888033ddf9d769ebf473c4a326187009cf02ec853ea4ffa84d4ec87f0c351b8759a7b4e1eb324d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb71eb1a1c9e8e63cf84f1fc5836022c18754cd28dde97b69487041279d7000e17cbc36aed380a83e9a361318b8af401770862274da59ebede969109808cfbe9ee43c6b6bad9e18c602160fef62c074356c40aac08227dbc82cf31e97ad78bc0685d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he169447000d261ba5128c3967f1741c25e2734a102ed50f2036f5fcf1ec3501166a598d948fba5ae91bc79e402ca7b5deeedab889db9d0087151171e18b8e6ae6b5e8a54233647957f76dd7d9974570a42cac279a6c55c002dc982da9027f1908a84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e2d068b20507c1fcdf032915938fc8cce6c2eefa38ae0114819cbe94edd9a779fc3f347d3f0455f23dc3d7f8c1d284ba415e02d2aff2cd0b4aa029683b60729f7dc3859ad7fb34702314c81ddcc5ac3310bbd1cc37894e91b98e8bffdccd8a8cb9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3c38ab53dedadf3cd71529e8f928bd1028428a193f1db4aeaa6c425b5852a3ba824d5462730446fc1c2e06fd1d453630ef8e0670ffb0835f358a2f82939e472a3fca2dd85810e761051452c76efe406547365dcf2173e51d4eb6686e1d7eff0d454;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6351df2ce690566eb946903b83c8fb0a63d35c0012998d3d24908b07a76a54090117d943cfcf250b3dc5f0985eeaae1fd06bca06a6d208418c25b7916db23e67e0230256a71276cac519cca6b1d9c87345deffb87984f9f9ea5e6c89be9bba73a52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b4860df3273e9fb97f1c0f090b27873e22110279b4d5bc8604bd633f81125be6c7f7ca59539eead1f5089ab758a10b1e2cb92a0c5dfc7ebaab7bf9e897b9a6e949d1cc2794b59edecbfc8043a45e485c4186fc8813b1be9d7da8890d563b913433e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e2e1c28fc6fcb81f53a52c560ab065349170b082fdc1c649888933d6411a56393939bad414bdda9f4b5ec22ab85f9fef4904609133ee209f2d20a8dda48bf60a509a1d63bce97f01a272558343eaea6e292d79036f85f4d29f6b0cd80700d51fb8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea76e2e43d0fcc593cecacf918e900caab9e9de6f42507cbddf67dfb5d19cfe64d1930c10186dcbe3badb55c16d5e929b5cec22a69be4db29eda220ec01ee5395fbf5a27bc0da7d7aa2bd53d8070f896f78fd6298e66bd35fd9b033f25185ffb18d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9584acec8cff45417965ab41343380e00b64c015b5d61eaa1ffd6d902de134becceb2ceec8b1a864be878ef2ecc42e88ae898767c088a3fa9020a1e93e736d53bd7ee5372201500cf0329e26ce492362b0a6b84c9958d69293ca0a444a68f61912ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69d3c66f8df0e4d9582c5d748ffffb1bb1ccc9cfbcc4cca28aa992c376a6516b369cfdc0ac74587b15bc374956092fd74026cb312bb603fcf1946d13c6b156f074b8728ba8c55783c46d6f9d660e022a8a36a67a82f35d8834273ff8e4b1257cd527;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11a3bd3acebc63d400797e277088187ba9e4f511470389a847d18f8b053aaf965a2ed9b7ded943600bc4de62c0cfaeaa613e41538243f2a5f058d721f89ba0afc89f87844d27d688893c0e8665f5f76cb3519c86c0582a5c9bda24c16028e45f1bec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83c46dd1237b4f7406d78780e8deae2357a064ba5879118f4d1ee89903fa72af9cdc7664ec9e8a1b235e47844f4e21c0580e66ada22abf03fe4578b0f22991317888416ca6cf82245e7119f9f2f88232281a52cb23a013f8c429d22bcd9e349c2a6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde8cd4a4f8eb620d86fa59a0aab4eee25f978bba5602a8a84f4ec740550814226db7cc7a86813c24fd7ca5aa99a7f8fb6c87b596173399ffa6ad6573a254dd89f002ec736933310a551bf2c72c5cd7d28e4ef3cefd7b0c914afa0d2dd0333efbc31d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h782476f9f43798e5d9e4455cfece0a72d33bb590cd2cc8cb0c3b8a4efbda9688837b3c5d901de3538fc8478acf3d96e0a48719ef390858eb67249375d7d99956d550a354b779437cb844548fdfd49d980d7c6009a8047234ea9313d5ac615ed795f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8148dd32209d88169ced7502627fc7a09e87c09a070ac221480cedbe63cb78f7aede6d522bfb859ebc8336a6d6e381e74180ecee2fc81fd2485ce21b42c73152eee2d4f7cbe2aceeb7aa8052a13d5fa7a38443e9bf422925ab2c40c907d414e304a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5629314170bdb14d4e93e5af1deea26906620d530ab36a3cdc4fe760db0b4e3f48f932934c34012ab271b507e1e4cfb4ca3d1e5f9a8feec58e798002cc718763b5d8f47ec502d678a77c1195237d7addf8dc7d738d8b010ecaf5b014a635374951ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he88702fec99a033f04630e1692b5a14a68eb49d906cab4ec643128d3c1a13f327ff7ac051caf1118d7de4e7386e6097d4a8f9c1f8214758abbbe32bce89f40145cd9bed5d638ec2e1a3c8f3775133822b6fa554c061c1298fcc36393d8fda16ca612;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd80a27991a582fc24ade2af1ca148557273c6f08472debcc8f68b344983c30baf1f291ae9c547d64d58626d363d9350980dc4044adb1e0b5b41f2f539ba90aa9715fc3e81da496e0a9d1f1068a5aa93ed4e11ff8cd74d5b277a0aab5f87e68e34a25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d06fc53cebacb3622864c15135a18156ddc575dbc10f50320c8c4a61616cbeccad9a9c22126981396f926f41ad7726d3f128a334b8a81c0686846cdf57e9d7e000cc451e0eabdd7ef8fd61dd0a48f69cabaada8702c26af96f6d32662a1b528f474;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h269a42707a98b0b8f20f3d482d84e85b1ea376a7324b66ebab7968989520917a62d81069af4a73f4a46ec78f05a799757b958f3b2cee206faaad1735ef992d86b128ebb725ebb65ac1eda82182fc69be5c3b73752f8ee164e9e7d10f8ed8d06713fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae7c2bcb02ecbadf190f5f89852a9abb230089ed1a29712bf209dbd648c9c83a332e765b7b560460709b02e37b1bf9c935ad2e6953c12de278d56f91ff4e150939546486010563a4f1a0526910beab8e0b6fc142bac8f879694a4e0c296a9271e3ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39324bf8971b76c850feffcd22e51ecabc23d3669e2f1e332fe1797caf1337ef9202e824884899192e535f47a592591e08455d430d4507d1ee30a296184802a6595ac1b6a7a39069e63cd196994867ab7fed3597e735cda4ac81b961b2220e430386;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f4d1279b72b0de6f609cfc1312dc8dc88415014b4fe03826b0c50e6f5a83155b47f7eff8ca9b50c8945eb7055890222376731e0a16e134238595e4e33fc2905df9f4724da93aede28f522bc9b37b09b8caf68c69e571ec46dec8a70a6cf1089a0dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heba3b3cd80ed2ecdbc769fafb13fde79587fc8280acf0adddc61bd5424ce2ae0e17529d9282316c9c3f409e032036ae32912e8e72c5d1cef16bd306050f1eaa149e0730a327b41ca07793c823fe615a0d8d2fb9ef1dcd366fc198d0cd1f3b37d01a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b63d6efbc4100e123254962baedac9e46188986fd85cac63c35d434f38fefdada705eedc7d45b93ddd04e87b79ba9b0d40f6c07fe72fe61afcb005bb0b9a92e355bb904a616d4cd0569a3802dd27b17d40795ecc1613d9a841136a7fbbb6b2ff79a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38d9c07a01493a5752fe9deb416ade4a4607f9d76bc82f30cf98c0230fc1642327bb8605dba83718ee82ba7c265732931ce7f0259f1287e2e31f3bdc9a8ef5c2a9ac38e3e771715ce7c5eb07094f504cdcbb73db925a04ce6c5c1b3c50094d72acca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7221a4ea8abd54b76578579cbb9dc827a08ea88a20fe7c19bda812aff064eee1db89d9f01f52241b11cbdca9e4aa25da51ad4604d206adfa83586ec17950936d1af19eff5091f0ac759204c0a752117ee1a1cebc33e7ef7ea6d77523374c18428715;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e28a92b5ac7377c988ccb8163fb253a18c424043d9596dee7e195c0dee71969788e9b22c3df8090b4053de4f5b615056a6433ea3b8f910dfff3316db6144cce015469edb2293aa7cd90d20913bd351c12492871e3884021732c82e1df7fe9b6ce4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6f036d3c7250651ea11890a6977de07d427d7dcb37a3c890d1b1880940974aa812c81979654484a65aae006452351054c79701bdb2c7e1a2686691721da361907a4136d8ad20322ce0c709d878682693b79819d361fdaa9b907ecc2c1536830478a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae06260e02b58db0ab4e8b49d80775cb82a1a5c9429820167f6c25edac86416d4f2edbcfdd6dcaedbc7f10f52995506d9d851b7558eb231425265955920059eadc13bcf2377347edec8c7bdee887d01857f72e3c6f9ee64419adce9be0289e1d53a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7257a97f3800d1304c1c77536f86c28109b2f3301fdedb0c985826609915874a22287b59ac1fd3e855b1242280770cbbbf66039bb58fd3bd8f56411da28373138f6f92239788ad21c91be01be8100bcd2580a438667ae738383423c7052945130b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdba9aecc162746018fc0c5162259b1f53dc39c033cc6ae801f9d95dad546eb8e48e215300a6b1c105b25d7ad0ff6757a37ab3a500c3d1fccb298e27557bbf3da6f1667c04c22df6da05b737494215e93d9fbcdd32ac72a8da36464296264a54b207;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50f054a01b7525482616e4be7159a9f65fe2d5216c6a1449809c926c2f1885c0fbbe9206854ca774e259b9a6556ab381b4aa5144c62fa4c3f9da96c4d6bb4b5e8fb8b57fb7c8135bba45e108c114e87b88692fbace5bfbb324e0b96e1cc10fddd6f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24996fb20a6fd36f1218b7713454ac837ee3810f6c0015c8f036445bd354c396026474a80fbd1810becc1f9899ac283bf449b08d90874c23d7589eb52cad11a84b0d270cc49f1f94db6b80085cf604e8752bc83c684fe4d9d15eb5e3e7a87b0c0378;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h388817d3cb4d6fb9506a42be45e705693983ed400871e4ffaeaca476daa3b7969834369b58a246f304ee500c5a2ec1aa76ce5adab92657626496cbe34faa3c9b0d8fc9f477d3c970c60fa2477912563976e00bb3da0907f7e256ec071bbcc79910e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57100e7dcbb223c758ccf6decb38908c09cd1760540e36ad20b144b4fcb24400c9411ebd11cca8df3c627f74a33c3cb1d7c83fbb46bf140910d2c2eed10421bfd359253349a6b71d9fa7c22f5c0f97170339f02361c67955d66b0856af2f54533170;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14017da0915b6c777975c3f66075d185dbecb063ee01873885b18d1b3d466a86c06808b75304ea73917096bad873f31dbe422180a00f3a87c06edb0470ac8eba0e3f024c60c29967807d2e2067f8f415a27d73c6d55e3f1d7ab4eb8c240779447344;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb029170c5deaedf58408824dceea30b461526eaa2a473739e1d7944446defc667efa020aece3dfde1d9d420f84dfa1e406be5585b3f4f7d6f24f14002add5192cf720cbdcabe6067ebde82a6091b52af5ad1c752499418952f415b0f5d49a7b6930b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4b292a1bdfe87b7527f7bfe205c9e7e985390f6400961044071caea0a8efecb509095c4b0fd71b6e7f729b61ab698a8d2086d078678a00baf3a80c9492194808b3429e1919dbfb3d202208b32d0b004c4843b28813adda325fe5deac52589c7b9f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5db7a1a591a5e92a08197f3aa3a5dd91b0165e8a2b6863cdebe400a2a5201caa1d021177eaac486f2e93f0f2b29a4dcb63f70bba3fc04563b791d446a6c1b6e574ae6c8b33ea76097e362701f1260f6aabc0867817385b8789923d76189588936f6c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ada2ac05b94517e6cdfe7780920d1b6fe659d99a1b09c3ef681f68727b0f165da0820bdd4f2a9a443285d1f106f0f048ff87fa3cb5920099f4c136a7425261645e40bff1b664d35a96e078297147002097a3b15edeeef0be14423b22252b3df52fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ba119a169a52a6ef688c41081009ac29bdc2b3c0af04814dab39e914d540a70fce19927781497eddc5db1544f9943ad60c12b27e779e831af244196e0e707efd4883cc0ae1b27c2aae3b34d746adf24329527f908fcde580023616abdca7c17f0fe;
        #1
        $finish();
    end
endmodule
